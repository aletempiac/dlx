
module DLX_IR_SIZE32_PC_SIZE32_DW01_inc_1 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106;

  XNOR2_X2 U2 ( .A(A[4]), .B(n54), .ZN(SUM[4]) );
  INV_X1 U3 ( .A(n32), .ZN(n54) );
  NOR2_X1 U4 ( .A1(n72), .A2(n24), .ZN(n1) );
  NAND2_X1 U5 ( .A1(n1), .A2(n2), .ZN(n66) );
  AND2_X1 U6 ( .A1(n3), .A2(A[26]), .ZN(n2) );
  INV_X1 U7 ( .A(n25), .ZN(n3) );
  OR2_X1 U8 ( .A1(n24), .A2(n72), .ZN(n4) );
  OR2_X1 U9 ( .A1(n20), .A2(n21), .ZN(n5) );
  OR2_X2 U10 ( .A1(n5), .A2(n6), .ZN(n85) );
  OR2_X1 U11 ( .A1(n7), .A2(n39), .ZN(n6) );
  INV_X1 U12 ( .A(A[18]), .ZN(n7) );
  INV_X1 U13 ( .A(A[25]), .ZN(n24) );
  NOR2_X1 U14 ( .A1(n24), .A2(n72), .ZN(n23) );
  NOR2_X1 U15 ( .A1(n59), .A2(n60), .ZN(n57) );
  XNOR2_X1 U16 ( .A(n57), .B(n58), .ZN(SUM[31]) );
  OR2_X2 U17 ( .A1(n20), .A2(n21), .ZN(n89) );
  NOR2_X2 U18 ( .A1(n43), .A2(n101), .ZN(n42) );
  OR2_X2 U19 ( .A1(n8), .A2(n9), .ZN(n101) );
  NOR2_X2 U20 ( .A1(n41), .A2(n85), .ZN(n40) );
  NAND2_X1 U21 ( .A1(n30), .A2(A[8]), .ZN(n8) );
  OR2_X1 U22 ( .A1(n10), .A2(n36), .ZN(n9) );
  INV_X1 U23 ( .A(A[10]), .ZN(n10) );
  NAND2_X1 U24 ( .A1(n40), .A2(A[20]), .ZN(n11) );
  OR2_X1 U25 ( .A1(n11), .A2(n12), .ZN(n76) );
  OR2_X1 U26 ( .A1(n13), .A2(n34), .ZN(n12) );
  INV_X1 U27 ( .A(A[22]), .ZN(n13) );
  OR2_X1 U28 ( .A1(n11), .A2(n12), .ZN(n14) );
  OR2_X2 U29 ( .A1(n14), .A2(n15), .ZN(n72) );
  OR2_X1 U30 ( .A1(n16), .A2(n29), .ZN(n15) );
  INV_X1 U31 ( .A(A[24]), .ZN(n16) );
  NAND2_X1 U32 ( .A1(n42), .A2(A[12]), .ZN(n17) );
  OR2_X1 U33 ( .A1(n17), .A2(n18), .ZN(n93) );
  OR2_X1 U34 ( .A1(n19), .A2(n27), .ZN(n18) );
  INV_X1 U35 ( .A(A[14]), .ZN(n19) );
  OR2_X1 U36 ( .A1(n17), .A2(n18), .ZN(n20) );
  OR2_X1 U37 ( .A1(n22), .A2(n45), .ZN(n21) );
  INV_X1 U38 ( .A(A[16]), .ZN(n22) );
  NOR2_X1 U39 ( .A1(n103), .A2(n36), .ZN(n35) );
  INV_X32 U40 ( .A(A[27]), .ZN(n25) );
  INV_X1 U41 ( .A(n26), .ZN(n94) );
  NOR2_X1 U42 ( .A1(n27), .A2(n97), .ZN(n26) );
  INV_X32 U43 ( .A(A[13]), .ZN(n27) );
  INV_X1 U44 ( .A(n28), .ZN(n73) );
  NOR2_X1 U45 ( .A1(n29), .A2(n76), .ZN(n28) );
  INV_X1 U46 ( .A(n35), .ZN(n102) );
  INV_X1 U47 ( .A(A[11]), .ZN(n43) );
  INV_X32 U48 ( .A(A[23]), .ZN(n29) );
  AND2_X1 U49 ( .A1(A[1]), .A2(A[0]), .ZN(n37) );
  INV_X1 U50 ( .A(n37), .ZN(n62) );
  INV_X2 U51 ( .A(n30), .ZN(n48) );
  INV_X2 U52 ( .A(n31), .ZN(n51) );
  NAND2_X1 U53 ( .A1(A[6]), .A2(n31), .ZN(n104) );
  NAND2_X1 U54 ( .A1(A[4]), .A2(n32), .ZN(n105) );
  AND2_X2 U55 ( .A1(A[7]), .A2(n49), .ZN(n30) );
  AND2_X2 U56 ( .A1(A[5]), .A2(n52), .ZN(n31) );
  NOR2_X1 U57 ( .A1(n34), .A2(n80), .ZN(n33) );
  INV_X1 U58 ( .A(A[9]), .ZN(n36) );
  INV_X1 U59 ( .A(n33), .ZN(n77) );
  AND2_X2 U60 ( .A1(A[3]), .A2(n55), .ZN(n32) );
  INV_X32 U61 ( .A(A[21]), .ZN(n34) );
  NOR2_X1 U62 ( .A1(n39), .A2(n89), .ZN(n38) );
  INV_X1 U63 ( .A(n38), .ZN(n86) );
  INV_X32 U64 ( .A(A[17]), .ZN(n39) );
  INV_X1 U65 ( .A(n42), .ZN(n98) );
  INV_X1 U66 ( .A(n40), .ZN(n81) );
  INV_X32 U67 ( .A(A[19]), .ZN(n41) );
  NOR2_X1 U68 ( .A1(n45), .A2(n93), .ZN(n44) );
  INV_X1 U69 ( .A(n44), .ZN(n90) );
  INV_X32 U70 ( .A(A[15]), .ZN(n45) );
  NAND2_X1 U71 ( .A1(A[8]), .A2(n30), .ZN(n103) );
  NAND2_X1 U72 ( .A1(A[28]), .A2(n65), .ZN(n64) );
  XNOR2_X1 U73 ( .A(A[6]), .B(n51), .ZN(SUM[6]) );
  XNOR2_X1 U74 ( .A(A[2]), .B(n62), .ZN(SUM[2]) );
  XNOR2_X1 U75 ( .A(A[26]), .B(n4), .ZN(SUM[26]) );
  XNOR2_X1 U76 ( .A(A[16]), .B(n90), .ZN(SUM[16]) );
  XNOR2_X1 U77 ( .A(A[22]), .B(n77), .ZN(SUM[22]) );
  XNOR2_X1 U78 ( .A(A[12]), .B(n98), .ZN(SUM[12]) );
  INV_X1 U79 ( .A(A[0]), .ZN(SUM[0]) );
  XNOR2_X1 U80 ( .A(A[10]), .B(n102), .ZN(SUM[10]) );
  XNOR2_X1 U81 ( .A(A[8]), .B(n48), .ZN(SUM[8]) );
  XNOR2_X1 U82 ( .A(A[20]), .B(n81), .ZN(SUM[20]) );
  XNOR2_X1 U83 ( .A(A[18]), .B(n86), .ZN(SUM[18]) );
  XNOR2_X1 U84 ( .A(A[28]), .B(n66), .ZN(SUM[28]) );
  XNOR2_X1 U85 ( .A(A[0]), .B(n83), .ZN(SUM[1]) );
  XNOR2_X1 U86 ( .A(A[24]), .B(n73), .ZN(SUM[24]) );
  XNOR2_X1 U87 ( .A(A[14]), .B(n94), .ZN(SUM[14]) );
  NAND2_X1 U88 ( .A1(A[29]), .A2(n61), .ZN(n59) );
  NAND2_X1 U89 ( .A1(A[26]), .A2(n23), .ZN(n69) );
  NAND2_X1 U90 ( .A1(A[20]), .A2(n40), .ZN(n80) );
  NAND2_X1 U91 ( .A1(A[12]), .A2(n42), .ZN(n97) );
  NAND2_X1 U92 ( .A1(A[2]), .A2(n37), .ZN(n106) );
  XNOR2_X1 U93 ( .A(n46), .B(n47), .ZN(SUM[9]) );
  INV_X2 U94 ( .A(A[9]), .ZN(n47) );
  XNOR2_X1 U95 ( .A(n49), .B(n50), .ZN(SUM[7]) );
  INV_X2 U96 ( .A(A[7]), .ZN(n50) );
  XNOR2_X1 U97 ( .A(n52), .B(n53), .ZN(SUM[5]) );
  INV_X2 U98 ( .A(A[5]), .ZN(n53) );
  XNOR2_X1 U99 ( .A(n55), .B(n56), .ZN(SUM[3]) );
  INV_X2 U100 ( .A(A[3]), .ZN(n56) );
  INV_X2 U101 ( .A(A[31]), .ZN(n58) );
  INV_X2 U102 ( .A(A[30]), .ZN(n60) );
  XNOR2_X2 U103 ( .A(A[30]), .B(n59), .ZN(SUM[30]) );
  XNOR2_X1 U104 ( .A(n61), .B(n63), .ZN(SUM[29]) );
  INV_X2 U105 ( .A(A[29]), .ZN(n63) );
  INV_X1 U106 ( .A(n64), .ZN(n61) );
  INV_X1 U107 ( .A(n66), .ZN(n65) );
  XNOR2_X1 U108 ( .A(n67), .B(n68), .ZN(SUM[27]) );
  INV_X2 U109 ( .A(A[27]), .ZN(n68) );
  INV_X1 U110 ( .A(n69), .ZN(n67) );
  XNOR2_X1 U111 ( .A(n70), .B(n71), .ZN(SUM[25]) );
  INV_X2 U112 ( .A(A[25]), .ZN(n71) );
  INV_X1 U113 ( .A(n72), .ZN(n70) );
  XNOR2_X1 U114 ( .A(n74), .B(n75), .ZN(SUM[23]) );
  INV_X2 U115 ( .A(A[23]), .ZN(n75) );
  INV_X1 U116 ( .A(n76), .ZN(n74) );
  XNOR2_X1 U117 ( .A(n78), .B(n79), .ZN(SUM[21]) );
  INV_X2 U118 ( .A(A[21]), .ZN(n79) );
  INV_X1 U119 ( .A(n80), .ZN(n78) );
  INV_X2 U120 ( .A(A[1]), .ZN(n83) );
  XNOR2_X1 U121 ( .A(n82), .B(n84), .ZN(SUM[19]) );
  INV_X2 U122 ( .A(A[19]), .ZN(n84) );
  INV_X1 U123 ( .A(n85), .ZN(n82) );
  XNOR2_X1 U124 ( .A(n87), .B(n88), .ZN(SUM[17]) );
  INV_X2 U125 ( .A(A[17]), .ZN(n88) );
  INV_X1 U126 ( .A(n89), .ZN(n87) );
  XNOR2_X1 U127 ( .A(n91), .B(n92), .ZN(SUM[15]) );
  INV_X2 U128 ( .A(A[15]), .ZN(n92) );
  INV_X1 U129 ( .A(n93), .ZN(n91) );
  XNOR2_X1 U130 ( .A(n95), .B(n96), .ZN(SUM[13]) );
  INV_X2 U131 ( .A(A[13]), .ZN(n96) );
  INV_X1 U132 ( .A(n97), .ZN(n95) );
  XNOR2_X1 U133 ( .A(n99), .B(n100), .ZN(SUM[11]) );
  INV_X2 U134 ( .A(A[11]), .ZN(n100) );
  INV_X1 U135 ( .A(n101), .ZN(n99) );
  INV_X1 U136 ( .A(n103), .ZN(n46) );
  INV_X1 U137 ( .A(n104), .ZN(n49) );
  INV_X1 U138 ( .A(n105), .ZN(n52) );
  INV_X1 U139 ( .A(n106), .ZN(n55) );
endmodule


module FA_1 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U1 ( .A(Ci), .B(n10), .Z(S) );
  INV_X1 U2 ( .A(n11), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n10), .B2(Ci), .ZN(n11) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n10) );
endmodule


module FA_2 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U1 ( .A(Ci), .B(n11), .Z(S) );
  INV_X1 U2 ( .A(n12), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
endmodule


module FA_3 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8;

  XOR2_X1 U1 ( .A(Ci), .B(n7), .Z(S) );
  INV_X1 U2 ( .A(n8), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n7) );
endmodule


module FA_4 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10;

  XOR2_X1 U1 ( .A(n8), .B(Ci), .Z(S) );
  INV_X1 U2 ( .A(n9), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(n10), .B1(n8), .B2(Ci), .ZN(n9) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n8) );
  CLKBUF_X1 U5 ( .A(A), .Z(n10) );
endmodule


module FA_5 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8;

  XOR2_X1 U1 ( .A(Ci), .B(n7), .Z(S) );
  INV_X1 U2 ( .A(n8), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n7) );
endmodule


module FA_6 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U1 ( .A(Ci), .B(n11), .Z(S) );
  INV_X1 U2 ( .A(n12), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
endmodule


module FA_7 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8;

  XOR2_X1 U1 ( .A(Ci), .B(n7), .Z(S) );
  INV_X1 U2 ( .A(n8), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n7) );
endmodule


module FA_8 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U1 ( .A(n8), .B(Ci), .Z(S) );
  INV_X1 U2 ( .A(n9), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n8) );
endmodule


module FA_9 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U1 ( .A(Ci), .B(n12), .Z(S) );
  INV_X1 U2 ( .A(n13), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n12), .B2(Ci), .ZN(n13) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n12) );
endmodule


module FA_10 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U1 ( .A(Ci), .B(n12), .Z(S) );
  INV_X1 U2 ( .A(n13), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n12), .B2(Ci), .ZN(n13) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n12) );
endmodule


module FA_11 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8;

  XOR2_X1 U1 ( .A(Ci), .B(n7), .Z(S) );
  INV_X1 U2 ( .A(n8), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n7) );
endmodule


module FA_12 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11;

  XOR2_X1 U1 ( .A(Ci), .B(n10), .Z(S) );
  INV_X1 U2 ( .A(n11), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n10), .B2(Ci), .ZN(n11) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n10) );
endmodule


module FA_13 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U1 ( .A(Ci), .B(n12), .Z(S) );
  INV_X1 U2 ( .A(n13), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n12), .B2(Ci), .ZN(n13) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n12) );
endmodule


module FA_14 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U1 ( .A(Ci), .B(n12), .Z(S) );
  INV_X1 U2 ( .A(n13), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n12), .B2(Ci), .ZN(n13) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n12) );
endmodule


module FA_15 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8;

  XOR2_X1 U1 ( .A(Ci), .B(n7), .Z(S) );
  INV_X1 U2 ( .A(n8), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n7) );
endmodule


module FA_16 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10;

  XOR2_X1 U1 ( .A(Ci), .B(n9), .Z(S) );
  INV_X1 U2 ( .A(n10), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n10) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
endmodule


module FA_17 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U1 ( .A(Ci), .B(n12), .Z(S) );
  INV_X1 U2 ( .A(n13), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n12), .B2(Ci), .ZN(n13) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n12) );
endmodule


module FA_18 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8;

  XOR2_X1 U1 ( .A(Ci), .B(n7), .Z(S) );
  INV_X1 U2 ( .A(n8), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n7) );
endmodule


module FA_19 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8;

  XOR2_X1 U1 ( .A(Ci), .B(n7), .Z(S) );
  INV_X1 U2 ( .A(n8), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n7) );
endmodule


module FA_20 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10;

  XOR2_X1 U1 ( .A(Ci), .B(n9), .Z(S) );
  INV_X1 U2 ( .A(n10), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n10) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
endmodule


module FA_21 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U1 ( .A(Ci), .B(n12), .Z(S) );
  INV_X1 U2 ( .A(n13), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n12), .B2(Ci), .ZN(n13) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n12) );
endmodule


module FA_22 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8;

  XOR2_X1 U1 ( .A(Ci), .B(n7), .Z(S) );
  INV_X1 U2 ( .A(n8), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n7) );
endmodule


module FA_23 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8;

  XOR2_X1 U1 ( .A(Ci), .B(n7), .Z(S) );
  INV_X1 U2 ( .A(n8), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n7) );
endmodule


module FA_24 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10;

  XOR2_X1 U1 ( .A(Ci), .B(n9), .Z(S) );
  INV_X1 U2 ( .A(n10), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n10) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
endmodule


module FA_25 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U1 ( .A(Ci), .B(n12), .Z(S) );
  INV_X1 U2 ( .A(n13), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n12), .B2(Ci), .ZN(n13) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n12) );
endmodule


module FA_26 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8;

  XOR2_X1 U1 ( .A(Ci), .B(n7), .Z(S) );
  INV_X1 U2 ( .A(n8), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n7) );
endmodule


module FA_27 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8;

  XOR2_X1 U1 ( .A(Ci), .B(n7), .Z(S) );
  INV_X1 U2 ( .A(n8), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n7) );
endmodule


module FA_28 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  XOR2_X1 U1 ( .A(Ci), .B(n11), .Z(S) );
  INV_X1 U2 ( .A(n10), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n10) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  CLKBUF_X1 U5 ( .A(n9), .Z(n11) );
endmodule


module FA_29 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U1 ( .A(Ci), .B(n8), .Z(S) );
  INV_X1 U2 ( .A(n9), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n8) );
endmodule


module FA_30 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8;

  XOR2_X1 U1 ( .A(Ci), .B(n7), .Z(S) );
  INV_X1 U2 ( .A(n8), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n7) );
endmodule


module FA_31 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8;

  XOR2_X1 U1 ( .A(Ci), .B(n7), .Z(S) );
  INV_X1 U2 ( .A(n8), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n7) );
endmodule


module FA_32 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10;

  XOR2_X1 U1 ( .A(Ci), .B(n10), .Z(S) );
  INV_X1 U2 ( .A(n9), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n8) );
  CLKBUF_X1 U5 ( .A(n8), .Z(n10) );
endmodule


module FA_33 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U1 ( .A(Ci), .B(n8), .Z(S) );
  INV_X1 U2 ( .A(n9), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n8) );
endmodule


module FA_34 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8;

  XOR2_X1 U1 ( .A(Ci), .B(n7), .Z(S) );
  INV_X1 U2 ( .A(n8), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n7) );
endmodule


module FA_35 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8;

  XOR2_X1 U1 ( .A(Ci), .B(n7), .Z(S) );
  INV_X1 U2 ( .A(n8), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n7) );
endmodule


module FA_36 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  XOR2_X1 U1 ( .A(Ci), .B(n11), .Z(S) );
  INV_X1 U2 ( .A(n10), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n10) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  CLKBUF_X1 U5 ( .A(n9), .Z(n11) );
endmodule


module FA_37 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U1 ( .A(Ci), .B(n8), .Z(S) );
  INV_X1 U2 ( .A(n9), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n8) );
endmodule


module FA_38 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8;

  XOR2_X1 U1 ( .A(Ci), .B(n7), .Z(S) );
  INV_X1 U2 ( .A(n8), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n7) );
endmodule


module FA_39 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8;

  XOR2_X1 U1 ( .A(Ci), .B(n7), .Z(S) );
  INV_X1 U2 ( .A(n8), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n7) );
endmodule


module FA_40 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10;

  XOR2_X1 U1 ( .A(Ci), .B(n10), .Z(S) );
  INV_X1 U2 ( .A(n9), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n8) );
  CLKBUF_X1 U5 ( .A(n8), .Z(n10) );
endmodule


module FA_41 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U1 ( .A(Ci), .B(n8), .Z(S) );
  INV_X1 U2 ( .A(n9), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n8) );
endmodule


module FA_42 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8;

  XOR2_X1 U1 ( .A(Ci), .B(n7), .Z(S) );
  INV_X1 U2 ( .A(n8), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n7) );
endmodule


module FA_43 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9, n10;

  XOR2_X1 U1 ( .A(Ci), .B(n7), .Z(S) );
  INV_X1 U2 ( .A(n8), .ZN(Co) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n7) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n7), .A2(Ci), .ZN(n10) );
  AND2_X1 U6 ( .A1(n9), .A2(n10), .ZN(n8) );
endmodule


module FA_44 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U1 ( .A(n8), .B(Ci), .Z(S) );
  INV_X1 U2 ( .A(n9), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n8) );
endmodule


module FA_45 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U1 ( .A(Ci), .B(n8), .Z(S) );
  INV_X1 U2 ( .A(n9), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n8) );
endmodule


module FA_46 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8;

  XOR2_X1 U1 ( .A(Ci), .B(n7), .Z(S) );
  INV_X1 U2 ( .A(n8), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n7) );
endmodule


module FA_47 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8;

  XOR2_X1 U1 ( .A(Ci), .B(n7), .Z(S) );
  INV_X1 U2 ( .A(n8), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n7) );
endmodule


module FA_48 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8;

  XOR2_X1 U1 ( .A(Ci), .B(n7), .Z(S) );
  INV_X1 U2 ( .A(n8), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n7) );
endmodule


module FA_49 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U1 ( .A(Ci), .B(n8), .Z(S) );
  INV_X1 U2 ( .A(n9), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n8) );
endmodule


module FA_50 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8;

  XOR2_X1 U1 ( .A(Ci), .B(n7), .Z(S) );
  INV_X1 U2 ( .A(n8), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n7) );
endmodule


module FA_51 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8;

  XOR2_X1 U1 ( .A(Ci), .B(n7), .Z(S) );
  INV_X1 U2 ( .A(n8), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n7) );
endmodule


module FA_52 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U1 ( .A(Ci), .B(n8), .Z(S) );
  INV_X1 U2 ( .A(n9), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n8) );
endmodule


module FA_53 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U1 ( .A(Ci), .B(n8), .Z(S) );
  INV_X1 U2 ( .A(n9), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n8) );
endmodule


module FA_54 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8;

  XOR2_X1 U1 ( .A(Ci), .B(n7), .Z(S) );
  INV_X1 U2 ( .A(n8), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n7) );
endmodule


module FA_55 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8;

  XOR2_X1 U1 ( .A(Ci), .B(n7), .Z(S) );
  INV_X1 U2 ( .A(n8), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n7) );
endmodule


module FA_56 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U1 ( .A(Ci), .B(n8), .Z(S) );
  INV_X1 U2 ( .A(n9), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n8) );
endmodule


module FA_57 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9;

  XOR2_X1 U1 ( .A(Ci), .B(n8), .Z(S) );
  INV_X1 U2 ( .A(n9), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n8), .B2(Ci), .ZN(n9) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n8) );
endmodule


module FA_58 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n10, n11, n12;

  XOR2_X1 U1 ( .A(n10), .B(n8), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n8) );
  NAND2_X1 U2 ( .A1(n11), .A2(n12), .ZN(Co) );
  CLKBUF_X1 U3 ( .A(Ci), .Z(n10) );
  NAND2_X1 U5 ( .A1(B), .A2(A), .ZN(n11) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n8), .ZN(n12) );
endmodule


module FA_59 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8;

  XOR2_X1 U1 ( .A(Ci), .B(n7), .Z(S) );
  INV_X1 U2 ( .A(n8), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(Ci), .B2(n7), .ZN(n8) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n7) );
endmodule


module FA_60 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n12, n13;

  XOR2_X1 U1 ( .A(n12), .B(Ci), .Z(S) );
  INV_X1 U2 ( .A(n13), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n12), .B2(Ci), .ZN(n13) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n12) );
endmodule


module FA_61 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10;

  XOR2_X1 U1 ( .A(Ci), .B(n9), .Z(S) );
  INV_X1 U2 ( .A(n10), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n10) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
endmodule


module FA_62 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8;

  XOR2_X1 U1 ( .A(Ci), .B(n7), .Z(S) );
  INV_X1 U2 ( .A(n8), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n7), .B2(Ci), .ZN(n8) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n7) );
endmodule


module FA_63 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  XOR2_X1 U1 ( .A(n9), .B(n7), .Z(S) );
  INV_X1 U2 ( .A(n8), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(Ci), .B2(n7), .ZN(n8) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n7) );
  CLKBUF_X1 U5 ( .A(Ci), .Z(n9) );
endmodule


module FA_0 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n12, n13, n14, n15;

  XOR2_X1 U1 ( .A(n10), .B(Ci), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n10) );
  OAI22_X1 U2 ( .A1(n12), .A2(n13), .B1(n14), .B2(n15), .ZN(Co) );
  INV_X1 U3 ( .A(B), .ZN(n12) );
  INV_X1 U5 ( .A(A), .ZN(n13) );
  INV_X1 U6 ( .A(n10), .ZN(n14) );
  INV_X1 U7 ( .A(Ci), .ZN(n15) );
endmodule


module RCA_N4_1 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:1] CTMP;

  FA_4 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_3 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_2 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_2 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:1] CTMP;

  FA_8 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_7 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_6 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_5 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_3 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:1] CTMP;

  FA_12 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_11 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_10 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_9 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_4 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:1] CTMP;

  FA_16 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_15 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_14 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_13 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_5 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:1] CTMP;

  FA_20 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_19 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_18 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_17 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_6 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:1] CTMP;

  FA_24 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_23 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_22 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_21 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_7 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:1] CTMP;

  FA_28 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_27 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_26 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_25 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_8 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:1] CTMP;

  FA_32 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_31 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_30 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_29 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_9 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:1] CTMP;

  FA_36 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_35 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_34 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_33 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_10 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:1] CTMP;

  FA_40 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_39 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_38 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_37 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_11 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:1] CTMP;

  FA_44 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_43 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_42 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_41 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_12 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:1] CTMP;

  FA_48 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_47 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_46 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_45 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_13 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:1] CTMP;

  FA_52 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_51 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_50 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_49 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_14 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:1] CTMP;

  FA_56 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_55 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_54 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_53 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_15 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:1] CTMP;

  FA_60 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_59 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_58 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_57 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_0 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:1] CTMP;

  FA_0 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_63 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_62 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_61 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module CSB_1 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_N4_2 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_N4_1 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX2_X2 U3 ( .A(sum0[3]), .B(sum1[3]), .S(Ci), .Z(S[3]) );
  MUX2_X1 U4 ( .A(sum0[2]), .B(sum1[2]), .S(Ci), .Z(S[2]) );
  MUX2_X2 U5 ( .A(sum0[0]), .B(sum1[0]), .S(Ci), .Z(S[0]) );
  MUX2_X2 U6 ( .A(sum0[1]), .B(sum1[1]), .S(Ci), .Z(S[1]) );
endmodule


module CSB_2 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  MUX2_X1 U4 ( .A(sum0[2]), .B(sum1[2]), .S(Ci), .Z(S[2]) );
  MUX2_X1 U5 ( .A(sum0[1]), .B(sum1[1]), .S(Ci), .Z(S[1]) );
  RCA_N4_4 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_N4_3 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX2_X1 U3 ( .A(sum0[0]), .B(sum1[0]), .S(Ci), .Z(S[0]) );
  MUX2_X1 U6 ( .A(sum0[3]), .B(sum1[3]), .S(Ci), .Z(S[3]) );
endmodule


module CSB_3 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  MUX2_X1 U3 ( .A(sum0[3]), .B(sum1[3]), .S(Ci), .Z(S[3]) );
  MUX2_X1 U4 ( .A(sum0[2]), .B(sum1[2]), .S(Ci), .Z(S[2]) );
  RCA_N4_6 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_N4_5 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX2_X1 U5 ( .A(sum0[0]), .B(sum1[0]), .S(Ci), .Z(S[0]) );
  MUX2_X1 U6 ( .A(sum0[1]), .B(sum1[1]), .S(Ci), .Z(S[1]) );
endmodule


module CSB_4 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_N4_8 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_N4_7 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX2_X1 U5 ( .A(sum0[1]), .B(sum1[1]), .S(Ci), .Z(S[1]) );
  MUX2_X1 U4 ( .A(sum0[2]), .B(sum1[2]), .S(Ci), .Z(S[2]) );
  MUX2_X1 U3 ( .A(sum0[3]), .B(sum1[3]), .S(Ci), .Z(S[3]) );
  MUX2_X1 U6 ( .A(sum0[0]), .B(sum1[0]), .S(Ci), .Z(S[0]) );
endmodule


module CSB_5 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  MUX2_X1 U3 ( .A(sum0[3]), .B(sum1[3]), .S(Ci), .Z(S[3]) );
  MUX2_X1 U4 ( .A(sum0[2]), .B(sum1[2]), .S(Ci), .Z(S[2]) );
  MUX2_X1 U5 ( .A(sum0[1]), .B(sum1[1]), .S(Ci), .Z(S[1]) );
  RCA_N4_10 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_N4_9 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX2_X1 U6 ( .A(sum0[0]), .B(sum1[0]), .S(Ci), .Z(S[0]) );
endmodule


module CSB_6 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  MUX2_X1 U3 ( .A(sum0[3]), .B(sum1[3]), .S(Ci), .Z(S[3]) );
  MUX2_X1 U4 ( .A(sum0[2]), .B(sum1[2]), .S(Ci), .Z(S[2]) );
  MUX2_X1 U5 ( .A(sum0[1]), .B(sum1[1]), .S(Ci), .Z(S[1]) );
  MUX2_X1 U6 ( .A(sum0[0]), .B(sum1[0]), .S(Ci), .Z(S[0]) );
  RCA_N4_12 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_N4_11 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
endmodule


module CSB_7 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  MUX2_X1 U4 ( .A(sum0[2]), .B(sum1[2]), .S(Ci), .Z(S[2]) );
  MUX2_X1 U5 ( .A(sum0[1]), .B(sum1[1]), .S(Ci), .Z(S[1]) );
  MUX2_X1 U6 ( .A(sum0[0]), .B(sum1[0]), .S(Ci), .Z(S[0]) );
  RCA_N4_14 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_N4_13 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX2_X2 U3 ( .A(sum0[3]), .B(sum1[3]), .S(Ci), .Z(S[3]) );
endmodule


module CSB_0 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  MUX2_X1 U4 ( .A(sum0[2]), .B(sum1[2]), .S(Ci), .Z(S[2]) );
  MUX2_X1 U5 ( .A(sum0[1]), .B(sum1[1]), .S(Ci), .Z(S[1]) );
  MUX2_X1 U6 ( .A(sum0[0]), .B(sum1[0]), .S(Ci), .Z(S[0]) );
  RCA_N4_0 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_N4_15 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX2_X2 U3 ( .A(sum0[3]), .B(sum1[3]), .S(Ci), .Z(S[3]) );
endmodule


module G_1 ( pi, gi, gj, gout );
  input pi, gi, gj;
  output gout;
  wire   n5, n6, n7;

  OAI21_X2 U1 ( .B1(n5), .B2(n6), .A(n7), .ZN(gout) );
  INV_X1 U2 ( .A(gj), .ZN(n5) );
  INV_X1 U3 ( .A(pi), .ZN(n6) );
  INV_X1 U4 ( .A(gi), .ZN(n7) );
endmodule


module G_2 ( pi, gi, gj, gout );
  input pi, gi, gj;
  output gout;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(gout) );
  AOI21_X1 U2 ( .B1(gj), .B2(pi), .A(gi), .ZN(n4) );
endmodule


module G_3 ( pi, gi, gj, gout );
  input pi, gi, gj;
  output gout;
  wire   n6;

  INV_X1 U1 ( .A(n6), .ZN(gout) );
  AOI21_X1 U2 ( .B1(gj), .B2(pi), .A(gi), .ZN(n6) );
endmodule


module G_4 ( pi, gi, gj, gout );
  input pi, gi, gj;
  output gout;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(gout) );
  AOI21_X1 U2 ( .B1(pi), .B2(gj), .A(gi), .ZN(n4) );
endmodule


module PG_1 ( pi, gi, pj, gj, pout, gout );
  input pi, gi, pj, gj;
  output pout, gout;
  wire   n4;

  AND2_X1 U1 ( .A1(pj), .A2(pi), .ZN(pout) );
  INV_X1 U2 ( .A(n4), .ZN(gout) );
  AOI21_X1 U3 ( .B1(gj), .B2(pi), .A(gi), .ZN(n4) );
endmodule


module PG_2 ( pi, gi, pj, gj, pout, gout );
  input pi, gi, pj, gj;
  output pout, gout;
  wire   n4;

  AND2_X1 U1 ( .A1(pj), .A2(pi), .ZN(pout) );
  INV_X1 U2 ( .A(n4), .ZN(gout) );
  AOI21_X1 U3 ( .B1(gj), .B2(pi), .A(gi), .ZN(n4) );
endmodule


module G_5 ( pi, gi, gj, gout );
  input pi, gi, gj;
  output gout;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(gout) );
  AOI21_X1 U2 ( .B1(pi), .B2(gj), .A(gi), .ZN(n4) );
endmodule


module G_6 ( pi, gi, gj, gout );
  input pi, gi, gj;
  output gout;
  wire   n6;

  INV_X1 U1 ( .A(n6), .ZN(gout) );
  AOI21_X1 U2 ( .B1(gj), .B2(pi), .A(gi), .ZN(n6) );
endmodule


module PG_3 ( pi, gi, pj, gj, pout, gout );
  input pi, gi, pj, gj;
  output pout, gout;
  wire   n4;

  AND2_X1 U1 ( .A1(pj), .A2(pi), .ZN(pout) );
  INV_X1 U2 ( .A(n4), .ZN(gout) );
  AOI21_X1 U3 ( .B1(gj), .B2(pi), .A(gi), .ZN(n4) );
endmodule


module PG_4 ( pi, gi, pj, gj, pout, gout );
  input pi, gi, pj, gj;
  output pout, gout;
  wire   n7;

  AND2_X1 U1 ( .A1(pj), .A2(pi), .ZN(pout) );
  INV_X1 U2 ( .A(n7), .ZN(gout) );
  AOI21_X1 U3 ( .B1(gj), .B2(pi), .A(gi), .ZN(n7) );
endmodule


module PG_5 ( pi, gi, pj, gj, pout, gout );
  input pi, gi, pj, gj;
  output pout, gout;
  wire   n6;

  AND2_X1 U1 ( .A1(pj), .A2(pi), .ZN(pout) );
  INV_X1 U2 ( .A(n6), .ZN(gout) );
  AOI21_X1 U3 ( .B1(gj), .B2(pi), .A(gi), .ZN(n6) );
endmodule


module G_7 ( pi, gi, gj, gout );
  input pi, gi, gj;
  output gout;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(gout) );
  AOI21_X1 U2 ( .B1(gj), .B2(pi), .A(gi), .ZN(n4) );
endmodule


module PG_6 ( pi, gi, pj, gj, pout, gout );
  input pi, gi, pj, gj;
  output pout, gout;
  wire   n4;

  AND2_X1 U1 ( .A1(pj), .A2(pi), .ZN(pout) );
  INV_X1 U2 ( .A(n4), .ZN(gout) );
  AOI21_X1 U3 ( .B1(gj), .B2(pi), .A(gi), .ZN(n4) );
endmodule


module PG_7 ( pi, gi, pj, gj, pout, gout );
  input pi, gi, pj, gj;
  output pout, gout;
  wire   n4;

  AND2_X1 U1 ( .A1(pj), .A2(pi), .ZN(pout) );
  INV_X1 U2 ( .A(n4), .ZN(gout) );
  AOI21_X1 U3 ( .B1(gj), .B2(pi), .A(gi), .ZN(n4) );
endmodule


module PG_8 ( pi, gi, pj, gj, pout, gout );
  input pi, gi, pj, gj;
  output pout, gout;
  wire   n4;

  AND2_X1 U1 ( .A1(pj), .A2(pi), .ZN(pout) );
  INV_X1 U2 ( .A(n4), .ZN(gout) );
  AOI21_X1 U3 ( .B1(gj), .B2(pi), .A(gi), .ZN(n4) );
endmodule


module PG_9 ( pi, gi, pj, gj, pout, gout );
  input pi, gi, pj, gj;
  output pout, gout;
  wire   n4;

  AND2_X1 U1 ( .A1(pj), .A2(pi), .ZN(pout) );
  INV_X1 U2 ( .A(n4), .ZN(gout) );
  AOI21_X1 U3 ( .B1(gj), .B2(pi), .A(gi), .ZN(n4) );
endmodule


module PG_10 ( pi, gi, pj, gj, pout, gout );
  input pi, gi, pj, gj;
  output pout, gout;
  wire   n4;

  AND2_X1 U1 ( .A1(pj), .A2(pi), .ZN(pout) );
  INV_X1 U2 ( .A(n4), .ZN(gout) );
  AOI21_X1 U3 ( .B1(gj), .B2(pi), .A(gi), .ZN(n4) );
endmodule


module PG_11 ( pi, gi, pj, gj, pout, gout );
  input pi, gi, pj, gj;
  output pout, gout;
  wire   n4;

  AND2_X1 U1 ( .A1(pj), .A2(pi), .ZN(pout) );
  INV_X1 U2 ( .A(n4), .ZN(gout) );
  AOI21_X1 U3 ( .B1(gj), .B2(pi), .A(gi), .ZN(n4) );
endmodule


module PG_12 ( pi, gi, pj, gj, pout, gout );
  input pi, gi, pj, gj;
  output pout, gout;
  wire   n4;

  AND2_X1 U1 ( .A1(pj), .A2(pi), .ZN(pout) );
  INV_X1 U2 ( .A(n4), .ZN(gout) );
  AOI21_X1 U3 ( .B1(gj), .B2(pi), .A(gi), .ZN(n4) );
endmodule


module G_8 ( pi, gi, gj, gout );
  input pi, gi, gj;
  output gout;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(gout) );
  AOI21_X1 U2 ( .B1(gj), .B2(pi), .A(gi), .ZN(n4) );
endmodule


module PG_13 ( pi, gi, pj, gj, pout, gout );
  input pi, gi, pj, gj;
  output pout, gout;
  wire   n4;

  AND2_X1 U1 ( .A1(pj), .A2(pi), .ZN(pout) );
  INV_X1 U2 ( .A(n4), .ZN(gout) );
  AOI21_X1 U3 ( .B1(gj), .B2(pi), .A(gi), .ZN(n4) );
endmodule


module PG_14 ( pi, gi, pj, gj, pout, gout );
  input pi, gi, pj, gj;
  output pout, gout;
  wire   n4;

  AND2_X1 U1 ( .A1(pj), .A2(pi), .ZN(pout) );
  INV_X1 U2 ( .A(n4), .ZN(gout) );
  AOI21_X1 U3 ( .B1(gj), .B2(pi), .A(gi), .ZN(n4) );
endmodule


module PG_15 ( pi, gi, pj, gj, pout, gout );
  input pi, gi, pj, gj;
  output pout, gout;
  wire   n4;

  AND2_X1 U1 ( .A1(pj), .A2(pi), .ZN(pout) );
  INV_X1 U2 ( .A(n4), .ZN(gout) );
  AOI21_X1 U3 ( .B1(gj), .B2(pi), .A(gi), .ZN(n4) );
endmodule


module PG_16 ( pi, gi, pj, gj, pout, gout );
  input pi, gi, pj, gj;
  output pout, gout;
  wire   n4;

  AND2_X1 U1 ( .A1(pj), .A2(pi), .ZN(pout) );
  INV_X1 U2 ( .A(n4), .ZN(gout) );
  AOI21_X1 U3 ( .B1(gj), .B2(pi), .A(gi), .ZN(n4) );
endmodule


module PG_17 ( pi, gi, pj, gj, pout, gout );
  input pi, gi, pj, gj;
  output pout, gout;
  wire   n4;

  AND2_X1 U1 ( .A1(pi), .A2(pj), .ZN(pout) );
  INV_X1 U2 ( .A(n4), .ZN(gout) );
  AOI21_X1 U3 ( .B1(pi), .B2(gj), .A(gi), .ZN(n4) );
endmodule


module PG_18 ( pi, gi, pj, gj, pout, gout );
  input pi, gi, pj, gj;
  output pout, gout;
  wire   n4;

  AND2_X1 U1 ( .A1(pj), .A2(pi), .ZN(pout) );
  INV_X1 U2 ( .A(n4), .ZN(gout) );
  AOI21_X1 U3 ( .B1(gj), .B2(pi), .A(gi), .ZN(n4) );
endmodule


module PG_19 ( pi, gi, pj, gj, pout, gout );
  input pi, gi, pj, gj;
  output pout, gout;
  wire   n4;

  AND2_X1 U1 ( .A1(pj), .A2(pi), .ZN(pout) );
  INV_X1 U2 ( .A(n4), .ZN(gout) );
  AOI21_X1 U3 ( .B1(pi), .B2(gj), .A(gi), .ZN(n4) );
endmodule


module PG_20 ( pi, gi, pj, gj, pout, gout );
  input pi, gi, pj, gj;
  output pout, gout;
  wire   n4;

  AND2_X1 U1 ( .A1(pj), .A2(pi), .ZN(pout) );
  INV_X1 U2 ( .A(n4), .ZN(gout) );
  AOI21_X1 U3 ( .B1(gj), .B2(pi), .A(gi), .ZN(n4) );
endmodule


module PG_21 ( pi, gi, pj, gj, pout, gout );
  input pi, gi, pj, gj;
  output pout, gout;
  wire   n6, n7, n8;

  OAI21_X1 U1 ( .B1(n6), .B2(n7), .A(n8), .ZN(gout) );
  INV_X1 U2 ( .A(pi), .ZN(n6) );
  INV_X1 U3 ( .A(gj), .ZN(n7) );
  INV_X1 U4 ( .A(gi), .ZN(n8) );
  AND2_X1 U5 ( .A1(pi), .A2(pj), .ZN(pout) );
endmodule


module PG_22 ( pi, gi, pj, gj, pout, gout );
  input pi, gi, pj, gj;
  output pout, gout;
  wire   n5;

  AND2_X1 U1 ( .A1(pi), .A2(pj), .ZN(pout) );
  INV_X1 U2 ( .A(n5), .ZN(gout) );
  AOI21_X1 U3 ( .B1(pi), .B2(gj), .A(gi), .ZN(n5) );
endmodule


module PG_23 ( pi, gi, pj, gj, pout, gout );
  input pi, gi, pj, gj;
  output pout, gout;
  wire   n5;

  AND2_X1 U1 ( .A1(pi), .A2(pj), .ZN(pout) );
  INV_X1 U2 ( .A(n5), .ZN(gout) );
  AOI21_X1 U3 ( .B1(pi), .B2(gj), .A(gi), .ZN(n5) );
endmodule


module PG_24 ( pi, gi, pj, gj, pout, gout );
  input pi, gi, pj, gj;
  output pout, gout;
  wire   n5;

  AND2_X1 U1 ( .A1(pj), .A2(pi), .ZN(pout) );
  INV_X1 U2 ( .A(n5), .ZN(gout) );
  AOI21_X1 U3 ( .B1(gj), .B2(pi), .A(gi), .ZN(n5) );
endmodule


module PG_25 ( pi, gi, pj, gj, pout, gout );
  input pi, gi, pj, gj;
  output pout, gout;
  wire   n7;

  AND2_X1 U1 ( .A1(pi), .A2(pj), .ZN(pout) );
  INV_X1 U2 ( .A(n7), .ZN(gout) );
  AOI21_X1 U3 ( .B1(pi), .B2(gj), .A(gi), .ZN(n7) );
endmodule


module PG_26 ( pi, gi, pj, gj, pout, gout );
  input pi, gi, pj, gj;
  output pout, gout;
  wire   n7;

  AND2_X1 U1 ( .A1(pi), .A2(pj), .ZN(pout) );
  INV_X1 U2 ( .A(n7), .ZN(gout) );
  AOI21_X1 U3 ( .B1(gj), .B2(pi), .A(gi), .ZN(n7) );
endmodule


module PG_0 ( pi, gi, pj, gj, pout, gout );
  input pi, gi, pj, gj;
  output pout, gout;
  wire   n7;

  AND2_X1 U1 ( .A1(pi), .A2(pj), .ZN(pout) );
  INV_X1 U2 ( .A(n7), .ZN(gout) );
  AOI21_X1 U3 ( .B1(pi), .B2(gj), .A(gi), .ZN(n7) );
endmodule


module G_0 ( pi, gi, gj, gout );
  input pi, gi, gj;
  output gout;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(gout) );
  AOI21_X1 U2 ( .B1(gj), .B2(pi), .A(gi), .ZN(n4) );
endmodule


module prop_gen_1 ( a, b, prop, gen );
  input a, b;
  output prop, gen;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(prop) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(gen) );
endmodule


module prop_gen_2 ( a, b, prop, gen );
  input a, b;
  output prop, gen;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(prop) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(gen) );
endmodule


module prop_gen_3 ( a, b, prop, gen );
  input a, b;
  output prop, gen;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(prop) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(gen) );
endmodule


module prop_gen_4 ( a, b, prop, gen );
  input a, b;
  output prop, gen;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(prop) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(gen) );
endmodule


module prop_gen_5 ( a, b, prop, gen );
  input a, b;
  output prop, gen;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(prop) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(gen) );
endmodule


module prop_gen_6 ( a, b, prop, gen );
  input a, b;
  output prop, gen;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(prop) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(gen) );
endmodule


module prop_gen_7 ( a, b, prop, gen );
  input a, b;
  output prop, gen;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(prop) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(gen) );
endmodule


module prop_gen_8 ( a, b, prop, gen );
  input a, b;
  output prop, gen;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(prop) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(gen) );
endmodule


module prop_gen_9 ( a, b, prop, gen );
  input a, b;
  output prop, gen;


  XOR2_X1 U1 ( .A(a), .B(b), .Z(prop) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(gen) );
endmodule


module prop_gen_10 ( a, b, prop, gen );
  input a, b;
  output prop, gen;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(prop) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(gen) );
endmodule


module prop_gen_11 ( a, b, prop, gen );
  input a, b;
  output prop, gen;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(prop) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(gen) );
endmodule


module prop_gen_12 ( a, b, prop, gen );
  input a, b;
  output prop, gen;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(prop) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(gen) );
endmodule


module prop_gen_13 ( a, b, prop, gen );
  input a, b;
  output prop, gen;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(prop) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(gen) );
endmodule


module prop_gen_14 ( a, b, prop, gen );
  input a, b;
  output prop, gen;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(prop) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(gen) );
endmodule


module prop_gen_15 ( a, b, prop, gen );
  input a, b;
  output prop, gen;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(prop) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(gen) );
endmodule


module prop_gen_16 ( a, b, prop, gen );
  input a, b;
  output prop, gen;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(prop) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(gen) );
endmodule


module prop_gen_17 ( a, b, prop, gen );
  input a, b;
  output prop, gen;


  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(gen) );
  XOR2_X1 U1 ( .A(a), .B(b), .Z(prop) );
endmodule


module prop_gen_18 ( a, b, prop, gen );
  input a, b;
  output prop, gen;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(prop) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(gen) );
endmodule


module prop_gen_19 ( a, b, prop, gen );
  input a, b;
  output prop, gen;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(prop) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(gen) );
endmodule


module prop_gen_20 ( a, b, prop, gen );
  input a, b;
  output prop, gen;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(prop) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(gen) );
endmodule


module prop_gen_21 ( a, b, prop, gen );
  input a, b;
  output prop, gen;


  XOR2_X1 U1 ( .A(a), .B(b), .Z(prop) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(gen) );
endmodule


module prop_gen_22 ( a, b, prop, gen );
  input a, b;
  output prop, gen;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(prop) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(gen) );
endmodule


module prop_gen_23 ( a, b, prop, gen );
  input a, b;
  output prop, gen;
  wire   n1;

  XOR2_X1 U1 ( .A(b), .B(a), .Z(prop) );
  AND2_X1 U2 ( .A1(b), .A2(n1), .ZN(gen) );
  CLKBUF_X1 U3 ( .A(a), .Z(n1) );
endmodule


module prop_gen_24 ( a, b, prop, gen );
  input a, b;
  output prop, gen;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(prop) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(gen) );
endmodule


module prop_gen_25 ( a, b, prop, gen );
  input a, b;
  output prop, gen;


  XOR2_X1 U1 ( .A(a), .B(b), .Z(prop) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(gen) );
endmodule


module prop_gen_26 ( a, b, prop, gen );
  input a, b;
  output prop, gen;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(prop) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(gen) );
endmodule


module prop_gen_27 ( a, b, prop, gen );
  input a, b;
  output prop, gen;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(prop) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(gen) );
endmodule


module prop_gen_28 ( a, b, prop, gen );
  input a, b;
  output prop, gen;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(prop) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(gen) );
endmodule


module prop_gen_29 ( a, b, prop, gen );
  input a, b;
  output prop, gen;
  wire   n1;

  AND2_X1 U2 ( .A1(b), .A2(n1), .ZN(gen) );
  XOR2_X1 U1 ( .A(b), .B(a), .Z(prop) );
  CLKBUF_X1 U3 ( .A(a), .Z(n1) );
endmodule


module prop_gen_30 ( a, b, prop, gen );
  input a, b;
  output prop, gen;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(prop) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(gen) );
endmodule


module prop_gen_0 ( a, b, prop, gen );
  input a, b;
  output prop, gen;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(prop) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(gen) );
endmodule


module prop_gen_Cin ( a, b, cin, prop, gen );
  input a, b, cin;
  output prop, gen;
  wire   n20, n21, n22;

  XOR2_X1 U1 ( .A(b), .B(n22), .Z(prop) );
  OAI21_X1 U5 ( .B1(a), .B2(b), .A(cin), .ZN(n20) );
  NAND2_X1 U2 ( .A1(n20), .A2(n21), .ZN(gen) );
  NAND2_X1 U3 ( .A1(a), .A2(b), .ZN(n21) );
  CLKBUF_X1 U4 ( .A(a), .Z(n22) );
endmodule


module shifter ( R, Offset, .Conf({\Conf[1] , \Conf[0] }), Shift_OUT );
  input [31:0] R;
  input [4:0] Offset;
  output [31:0] Shift_OUT;
  input \Conf[1] , \Conf[0] ;
  wire   \finegrainsel[0] , n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497;
  assign \finegrainsel[0]  = Offset[0];

  AOI221_X1 U2 ( .B1(n324), .B2(R[21]), .C1(n325), .C2(R[5]), .A(n479), .ZN(
        n281) );
  AOI221_X1 U3 ( .B1(n324), .B2(R[25]), .C1(n325), .C2(R[9]), .A(n326), .ZN(
        n256) );
  AOI222_X1 U4 ( .A1(n423), .A2(R[31]), .B1(R[7]), .B2(n298), .C1(R[15]), .C2(
        n299), .ZN(n430) );
  NOR3_X2 U5 ( .A1(n470), .A2(Offset[3]), .A3(n372), .ZN(n324) );
  NOR2_X2 U6 ( .A1(n486), .A2(n487), .ZN(n257) );
  NOR2_X2 U7 ( .A1(n483), .A2(n486), .ZN(n259) );
  NOR3_X2 U8 ( .A1(Offset[3]), .A2(Offset[4]), .A3(n470), .ZN(n325) );
  NOR3_X2 U9 ( .A1(n371), .A2(Offset[3]), .A3(n372), .ZN(n338) );
  NOR3_X4 U10 ( .A1(n470), .A2(Offset[4]), .A3(n370), .ZN(n423) );
  NOR2_X2 U11 ( .A1(n484), .A2(n487), .ZN(n270) );
  NOR3_X4 U12 ( .A1(n371), .A2(Offset[4]), .A3(n370), .ZN(n298) );
  NOR2_X4 U13 ( .A1(n483), .A2(n484), .ZN(n268) );
  NOR3_X4 U14 ( .A1(Offset[3]), .A2(Offset[4]), .A3(n371), .ZN(n299) );
  MUX2_X1 U15 ( .A(n247), .B(n248), .S(\finegrainsel[0] ), .Z(Shift_OUT[9]) );
  MUX2_X1 U16 ( .A(n249), .B(n247), .S(\finegrainsel[0] ), .Z(Shift_OUT[8]) );
  INV_X1 U17 ( .A(n250), .ZN(n247) );
  OAI221_X1 U18 ( .B1(n251), .B2(n252), .C1(n253), .C2(n254), .A(n255), .ZN(
        n250) );
  AOI22_X1 U19 ( .A1(n256), .A2(n257), .B1(n258), .B2(n259), .ZN(n255) );
  MUX2_X1 U20 ( .A(n260), .B(n249), .S(\finegrainsel[0] ), .Z(Shift_OUT[7]) );
  INV_X1 U21 ( .A(n261), .ZN(n249) );
  OAI221_X1 U22 ( .B1(n262), .B2(n263), .C1(n264), .C2(n265), .A(n266), .ZN(
        n261) );
  AOI22_X1 U23 ( .A1(n267), .A2(n268), .B1(n269), .B2(n270), .ZN(n266) );
  MUX2_X1 U24 ( .A(n271), .B(n260), .S(\finegrainsel[0] ), .Z(Shift_OUT[6]) );
  INV_X1 U25 ( .A(n272), .ZN(n260) );
  OAI221_X1 U26 ( .B1(n251), .B2(n254), .C1(n262), .C2(n273), .A(n274), .ZN(
        n272) );
  AOI22_X1 U27 ( .A1(n256), .A2(n259), .B1(n258), .B2(n270), .ZN(n274) );
  INV_X1 U28 ( .A(n275), .ZN(n273) );
  MUX2_X1 U29 ( .A(n276), .B(n271), .S(\finegrainsel[0] ), .Z(Shift_OUT[5]) );
  INV_X1 U30 ( .A(n277), .ZN(n271) );
  OAI221_X1 U31 ( .B1(n265), .B2(n263), .C1(n264), .C2(n253), .A(n278), .ZN(
        n277) );
  AOI22_X1 U32 ( .A1(n269), .A2(n268), .B1(n279), .B2(n257), .ZN(n278) );
  MUX2_X1 U33 ( .A(n280), .B(n276), .S(\finegrainsel[0] ), .Z(Shift_OUT[4]) );
  AOI221_X1 U34 ( .B1(n259), .B2(n275), .C1(n257), .C2(n281), .A(n282), .ZN(
        n276) );
  INV_X1 U35 ( .A(n283), .ZN(n282) );
  AOI22_X1 U36 ( .A1(n256), .A2(n270), .B1(n258), .B2(n268), .ZN(n283) );
  MUX2_X1 U37 ( .A(n284), .B(n280), .S(\finegrainsel[0] ), .Z(Shift_OUT[3]) );
  INV_X1 U38 ( .A(n285), .ZN(n280) );
  OAI221_X1 U39 ( .B1(n253), .B2(n263), .C1(n264), .C2(n251), .A(n286), .ZN(
        n285) );
  AOI22_X1 U40 ( .A1(n287), .A2(n257), .B1(n279), .B2(n259), .ZN(n286) );
  INV_X1 U41 ( .A(n288), .ZN(n279) );
  INV_X1 U42 ( .A(n289), .ZN(n263) );
  MUX2_X1 U43 ( .A(n290), .B(n291), .S(\finegrainsel[0] ), .Z(Shift_OUT[31])
         );
  OAI221_X1 U44 ( .B1(n292), .B2(n251), .C1(n293), .C2(n253), .A(n294), .ZN(
        n291) );
  AOI22_X1 U45 ( .A1(n259), .A2(n295), .B1(n257), .B2(n296), .ZN(n294) );
  INV_X1 U46 ( .A(n297), .ZN(n295) );
  AOI221_X1 U47 ( .B1(R[22]), .B2(n298), .C1(R[30]), .C2(n299), .A(n300), .ZN(
        n292) );
  OAI221_X1 U48 ( .B1(n301), .B2(n302), .C1(n303), .C2(n304), .A(n305), .ZN(
        n300) );
  MUX2_X1 U49 ( .A(n306), .B(n290), .S(\finegrainsel[0] ), .Z(Shift_OUT[30])
         );
  INV_X1 U50 ( .A(n307), .ZN(n290) );
  OAI221_X1 U51 ( .B1(n308), .B2(n309), .C1(n253), .C2(n310), .A(n311), .ZN(
        n307) );
  AOI22_X1 U52 ( .A1(n312), .A2(n259), .B1(n313), .B2(n257), .ZN(n311) );
  OAI221_X1 U53 ( .B1(n314), .B2(n315), .C1(n316), .C2(n317), .A(n268), .ZN(
        n309) );
  OAI221_X1 U54 ( .B1(n318), .B2(n302), .C1(n319), .C2(n304), .A(n305), .ZN(
        n308) );
  MUX2_X1 U55 ( .A(n320), .B(n284), .S(\finegrainsel[0] ), .Z(Shift_OUT[2]) );
  AOI221_X1 U56 ( .B1(n257), .B2(n321), .C1(n270), .C2(n275), .A(n322), .ZN(
        n284) );
  INV_X1 U57 ( .A(n323), .ZN(n322) );
  AOI22_X1 U58 ( .A1(n256), .A2(n268), .B1(n281), .B2(n259), .ZN(n323) );
  OAI221_X1 U59 ( .B1(n327), .B2(n328), .C1(n329), .C2(n316), .A(n330), .ZN(
        n326) );
  MUX2_X1 U60 ( .A(n331), .B(n306), .S(\finegrainsel[0] ), .Z(Shift_OUT[29])
         );
  AOI221_X1 U61 ( .B1(n268), .B2(n293), .C1(n270), .C2(n297), .A(n332), .ZN(
        n306) );
  OAI22_X1 U62 ( .A1(n296), .A2(n265), .B1(n333), .B2(n262), .ZN(n332) );
  INV_X1 U63 ( .A(n334), .ZN(n293) );
  OAI221_X1 U64 ( .B1(n316), .B2(n335), .C1(n314), .C2(n336), .A(n337), .ZN(
        n334) );
  MUX2_X1 U66 ( .A(n341), .B(n331), .S(\finegrainsel[0] ), .Z(Shift_OUT[28])
         );
  INV_X1 U67 ( .A(n342), .ZN(n331) );
  OAI221_X1 U68 ( .B1(n251), .B2(n310), .C1(n253), .C2(n343), .A(n344), .ZN(
        n342) );
  AOI22_X1 U69 ( .A1(n313), .A2(n259), .B1(n345), .B2(n257), .ZN(n344) );
  OAI221_X1 U70 ( .B1(n316), .B2(n346), .C1(n314), .C2(n347), .A(n348), .ZN(
        n310) );
  MUX2_X1 U72 ( .A(n349), .B(n341), .S(\finegrainsel[0] ), .Z(Shift_OUT[27])
         );
  AOI221_X1 U73 ( .B1(n268), .B2(n297), .C1(n270), .C2(n350), .A(n351), .ZN(
        n341) );
  OAI22_X1 U74 ( .A1(n333), .A2(n265), .B1(n352), .B2(n262), .ZN(n351) );
  AOI221_X1 U75 ( .B1(R[18]), .B2(n298), .C1(n299), .C2(R[26]), .A(n353), .ZN(
        n297) );
  OAI221_X1 U76 ( .B1(n304), .B2(n354), .C1(n302), .C2(n355), .A(n305), .ZN(
        n353) );
  INV_X1 U77 ( .A(n339), .ZN(n302) );
  INV_X1 U78 ( .A(n338), .ZN(n304) );
  MUX2_X1 U79 ( .A(n356), .B(n349), .S(\finegrainsel[0] ), .Z(Shift_OUT[26])
         );
  AOI221_X1 U80 ( .B1(n268), .B2(n312), .C1(n270), .C2(n313), .A(n357), .ZN(
        n349) );
  OAI22_X1 U81 ( .A1(n358), .A2(n265), .B1(n359), .B2(n262), .ZN(n357) );
  INV_X1 U82 ( .A(n360), .ZN(n313) );
  INV_X1 U83 ( .A(n343), .ZN(n312) );
  OAI221_X1 U84 ( .B1(n314), .B2(n327), .C1(n316), .C2(n361), .A(n362), .ZN(
        n343) );
  MUX2_X1 U86 ( .A(n363), .B(n356), .S(\finegrainsel[0] ), .Z(Shift_OUT[25])
         );
  AOI221_X1 U87 ( .B1(n268), .B2(n350), .C1(n270), .C2(n364), .A(n365), .ZN(
        n356) );
  OAI22_X1 U88 ( .A1(n352), .A2(n265), .B1(n366), .B2(n262), .ZN(n365) );
  INV_X1 U89 ( .A(n296), .ZN(n350) );
  OAI221_X1 U90 ( .B1(n314), .B2(n367), .C1(n316), .C2(n368), .A(n369), .ZN(
        n296) );
  NOR3_X1 U92 ( .A1(n370), .A2(n371), .A3(n372), .ZN(n339) );
  MUX2_X1 U93 ( .A(n373), .B(n363), .S(\finegrainsel[0] ), .Z(Shift_OUT[24])
         );
  AOI221_X1 U94 ( .B1(n259), .B2(n374), .C1(n257), .C2(n375), .A(n376), .ZN(
        n363) );
  OAI22_X1 U95 ( .A1(n360), .A2(n251), .B1(n358), .B2(n253), .ZN(n376) );
  OAI211_X1 U96 ( .C1(n377), .C2(n378), .A(n379), .B(n380), .ZN(n360) );
  AOI222_X1 U97 ( .A1(R[23]), .A2(n299), .B1(n338), .B2(R[7]), .C1(R[15]), 
        .C2(n298), .ZN(n380) );
  MUX2_X1 U98 ( .A(n381), .B(n373), .S(\finegrainsel[0] ), .Z(Shift_OUT[23])
         );
  AOI221_X1 U99 ( .B1(n268), .B2(n364), .C1(n270), .C2(n382), .A(n383), .ZN(
        n373) );
  OAI22_X1 U100 ( .A1(n366), .A2(n265), .B1(n384), .B2(n262), .ZN(n383) );
  INV_X1 U101 ( .A(n333), .ZN(n364) );
  OAI211_X1 U102 ( .C1(n378), .C2(n385), .A(n379), .B(n386), .ZN(n333) );
  AOI222_X1 U103 ( .A1(R[22]), .A2(n299), .B1(n338), .B2(R[6]), .C1(R[14]), 
        .C2(n298), .ZN(n386) );
  MUX2_X1 U104 ( .A(n387), .B(n381), .S(\finegrainsel[0] ), .Z(Shift_OUT[22])
         );
  AOI221_X1 U105 ( .B1(n268), .B2(n345), .C1(n270), .C2(n374), .A(n388), .ZN(
        n381) );
  OAI22_X1 U106 ( .A1(n389), .A2(n265), .B1(n390), .B2(n262), .ZN(n388) );
  INV_X1 U107 ( .A(n358), .ZN(n345) );
  OAI211_X1 U108 ( .C1(n378), .C2(n317), .A(n379), .B(n391), .ZN(n358) );
  AOI222_X1 U109 ( .A1(R[21]), .A2(n299), .B1(n338), .B2(R[5]), .C1(R[13]), 
        .C2(n298), .ZN(n391) );
  MUX2_X1 U110 ( .A(n392), .B(n387), .S(\finegrainsel[0] ), .Z(Shift_OUT[21])
         );
  AOI221_X1 U111 ( .B1(n268), .B2(n382), .C1(n270), .C2(n393), .A(n394), .ZN(
        n387) );
  OAI22_X1 U112 ( .A1(n384), .A2(n265), .B1(n395), .B2(n262), .ZN(n394) );
  INV_X1 U113 ( .A(n352), .ZN(n382) );
  OAI211_X1 U114 ( .C1(n378), .C2(n335), .A(n379), .B(n396), .ZN(n352) );
  AOI222_X1 U115 ( .A1(R[20]), .A2(n299), .B1(n338), .B2(R[4]), .C1(R[12]), 
        .C2(n298), .ZN(n396) );
  MUX2_X1 U116 ( .A(n397), .B(n392), .S(\finegrainsel[0] ), .Z(Shift_OUT[20])
         );
  AOI221_X1 U117 ( .B1(n268), .B2(n374), .C1(n270), .C2(n375), .A(n398), .ZN(
        n392) );
  OAI22_X1 U118 ( .A1(n390), .A2(n265), .B1(n399), .B2(n262), .ZN(n398) );
  INV_X1 U119 ( .A(n389), .ZN(n375) );
  INV_X1 U120 ( .A(n359), .ZN(n374) );
  OAI211_X1 U121 ( .C1(n378), .C2(n346), .A(n379), .B(n400), .ZN(n359) );
  AOI222_X1 U122 ( .A1(R[19]), .A2(n299), .B1(n338), .B2(R[3]), .C1(R[11]), 
        .C2(n298), .ZN(n400) );
  MUX2_X1 U123 ( .A(n401), .B(n320), .S(\finegrainsel[0] ), .Z(Shift_OUT[1])
         );
  INV_X1 U124 ( .A(n402), .ZN(n320) );
  OAI221_X1 U125 ( .B1(n262), .B2(n403), .C1(n253), .C2(n288), .A(n404), .ZN(
        n402) );
  AOI22_X1 U126 ( .A1(n289), .A2(n268), .B1(n287), .B2(n259), .ZN(n404) );
  AOI221_X1 U127 ( .B1(n324), .B2(R[24]), .C1(n325), .C2(R[8]), .A(n405), .ZN(
        n289) );
  OAI221_X1 U128 ( .B1(n367), .B2(n328), .C1(n406), .C2(n316), .A(n330), .ZN(
        n405) );
  MUX2_X1 U129 ( .A(n407), .B(n397), .S(\finegrainsel[0] ), .Z(Shift_OUT[19])
         );
  AOI221_X1 U130 ( .B1(n268), .B2(n393), .C1(n270), .C2(n408), .A(n409), .ZN(
        n397) );
  OAI22_X1 U131 ( .A1(n395), .A2(n265), .B1(n410), .B2(n262), .ZN(n409) );
  INV_X1 U132 ( .A(n366), .ZN(n393) );
  OAI211_X1 U133 ( .C1(n411), .C2(n378), .A(n379), .B(n412), .ZN(n366) );
  AOI222_X1 U134 ( .A1(R[18]), .A2(n299), .B1(n338), .B2(R[2]), .C1(n298), 
        .C2(R[10]), .ZN(n412) );
  MUX2_X1 U135 ( .A(n413), .B(n407), .S(\finegrainsel[0] ), .Z(Shift_OUT[18])
         );
  AOI221_X1 U136 ( .B1(n259), .B2(n414), .C1(n257), .C2(n415), .A(n416), .ZN(
        n407) );
  OAI22_X1 U137 ( .A1(n389), .A2(n251), .B1(n390), .B2(n253), .ZN(n416) );
  OAI211_X1 U138 ( .C1(n378), .C2(n361), .A(n379), .B(n417), .ZN(n389) );
  AOI222_X1 U139 ( .A1(R[17]), .A2(n299), .B1(n338), .B2(R[1]), .C1(R[9]), 
        .C2(n298), .ZN(n417) );
  MUX2_X1 U140 ( .A(n418), .B(n413), .S(\finegrainsel[0] ), .Z(Shift_OUT[17])
         );
  AOI221_X1 U141 ( .B1(n268), .B2(n408), .C1(n270), .C2(n419), .A(n420), .ZN(
        n413) );
  OAI22_X1 U142 ( .A1(n410), .A2(n265), .B1(n421), .B2(n262), .ZN(n420) );
  INV_X1 U143 ( .A(n384), .ZN(n408) );
  OAI211_X1 U144 ( .C1(n378), .C2(n368), .A(n379), .B(n422), .ZN(n384) );
  AOI222_X1 U145 ( .A1(R[16]), .A2(n299), .B1(n338), .B2(R[0]), .C1(R[8]), 
        .C2(n298), .ZN(n422) );
  MUX2_X1 U147 ( .A(n425), .B(n418), .S(\finegrainsel[0] ), .Z(Shift_OUT[16])
         );
  AOI221_X1 U148 ( .B1(n259), .B2(n415), .C1(n257), .C2(n426), .A(n427), .ZN(
        n418) );
  OAI22_X1 U149 ( .A1(n390), .A2(n251), .B1(n399), .B2(n253), .ZN(n427) );
  INV_X1 U150 ( .A(n414), .ZN(n399) );
  OAI211_X1 U151 ( .C1(n378), .C2(n428), .A(n497), .B(n430), .ZN(n390) );
  MUX2_X1 U152 ( .A(n431), .B(n425), .S(\finegrainsel[0] ), .Z(Shift_OUT[15])
         );
  AOI221_X1 U153 ( .B1(n268), .B2(n419), .C1(n270), .C2(n432), .A(n433), .ZN(
        n425) );
  OAI22_X1 U154 ( .A1(n421), .A2(n265), .B1(n434), .B2(n262), .ZN(n433) );
  INV_X1 U155 ( .A(n395), .ZN(n419) );
  OAI211_X1 U156 ( .C1(n328), .C2(n385), .A(n497), .B(n435), .ZN(n395) );
  AOI222_X1 U157 ( .A1(R[14]), .A2(n299), .B1(R[6]), .B2(n298), .C1(R[22]), 
        .C2(n325), .ZN(n435) );
  MUX2_X1 U158 ( .A(n436), .B(n431), .S(\finegrainsel[0] ), .Z(Shift_OUT[14])
         );
  INV_X1 U159 ( .A(n437), .ZN(n431) );
  OAI221_X1 U160 ( .B1(n265), .B2(n438), .C1(n262), .C2(n252), .A(n439), .ZN(
        n437) );
  AOI22_X1 U161 ( .A1(n414), .A2(n268), .B1(n415), .B2(n270), .ZN(n439) );
  AOI211_X1 U162 ( .C1(n325), .C2(R[21]), .A(n424), .B(n440), .ZN(n414) );
  OAI222_X1 U163 ( .A1(n317), .A2(n328), .B1(n318), .B2(n314), .C1(n319), .C2(
        n316), .ZN(n440) );
  INV_X1 U164 ( .A(R[5]), .ZN(n318) );
  MUX2_X1 U165 ( .A(n441), .B(n436), .S(\finegrainsel[0] ), .Z(Shift_OUT[13])
         );
  AOI221_X1 U166 ( .B1(n257), .B2(n267), .C1(n268), .C2(n432), .A(n442), .ZN(
        n436) );
  OAI22_X1 U167 ( .A1(n421), .A2(n253), .B1(n265), .B2(n434), .ZN(n442) );
  INV_X1 U168 ( .A(n410), .ZN(n432) );
  OAI211_X1 U169 ( .C1(n378), .C2(n336), .A(n497), .B(n443), .ZN(n410) );
  AOI222_X1 U170 ( .A1(R[28]), .A2(n423), .B1(R[4]), .B2(n298), .C1(R[12]), 
        .C2(n299), .ZN(n443) );
  MUX2_X1 U171 ( .A(n444), .B(n441), .S(\finegrainsel[0] ), .Z(Shift_OUT[12])
         );
  INV_X1 U172 ( .A(n445), .ZN(n441) );
  OAI221_X1 U173 ( .B1(n265), .B2(n252), .C1(n262), .C2(n254), .A(n446), .ZN(
        n445) );
  AOI22_X1 U174 ( .A1(n415), .A2(n268), .B1(n426), .B2(n270), .ZN(n446) );
  INV_X1 U175 ( .A(n447), .ZN(n415) );
  OAI211_X1 U176 ( .C1(n328), .C2(n346), .A(n497), .B(n448), .ZN(n447) );
  AOI222_X1 U177 ( .A1(R[11]), .A2(n299), .B1(R[3]), .B2(n298), .C1(R[19]), 
        .C2(n325), .ZN(n448) );
  MUX2_X1 U178 ( .A(n449), .B(n444), .S(\finegrainsel[0] ), .Z(Shift_OUT[11])
         );
  AOI221_X1 U179 ( .B1(n267), .B2(n259), .C1(n257), .C2(n269), .A(n450), .ZN(
        n444) );
  OAI22_X1 U180 ( .A1(n421), .A2(n251), .B1(n253), .B2(n434), .ZN(n450) );
  INV_X1 U181 ( .A(n451), .ZN(n421) );
  AOI211_X1 U182 ( .C1(R[18]), .C2(n325), .A(n424), .B(n452), .ZN(n451) );
  OAI222_X1 U183 ( .A1(n411), .A2(n328), .B1(n314), .B2(n355), .C1(n354), .C2(
        n316), .ZN(n452) );
  INV_X1 U184 ( .A(n298), .ZN(n314) );
  INV_X1 U185 ( .A(n496), .ZN(n424) );
  MUX2_X1 U186 ( .A(n248), .B(n449), .S(\finegrainsel[0] ), .Z(Shift_OUT[10])
         );
  INV_X1 U187 ( .A(n453), .ZN(n449) );
  OAI221_X1 U188 ( .B1(n253), .B2(n252), .C1(n265), .C2(n254), .A(n454), .ZN(
        n453) );
  AOI22_X1 U189 ( .A1(n258), .A2(n257), .B1(n426), .B2(n268), .ZN(n454) );
  INV_X1 U190 ( .A(n438), .ZN(n426) );
  OAI211_X1 U191 ( .C1(n378), .C2(n327), .A(n497), .B(n455), .ZN(n438) );
  AOI222_X1 U192 ( .A1(R[25]), .A2(n423), .B1(R[1]), .B2(n298), .C1(R[9]), 
        .C2(n299), .ZN(n455) );
  AOI221_X1 U193 ( .B1(n423), .B2(R[19]), .C1(n325), .C2(R[11]), .A(n456), 
        .ZN(n258) );
  OAI221_X1 U194 ( .B1(n346), .B2(n457), .C1(n458), .C2(n316), .A(n330), .ZN(
        n456) );
  INV_X1 U195 ( .A(R[3]), .ZN(n458) );
  OAI221_X1 U196 ( .B1(n328), .B2(n315), .C1(n378), .C2(n319), .A(n459), .ZN(
        n254) );
  AOI221_X1 U197 ( .B1(R[29]), .B2(n324), .C1(R[5]), .C2(n299), .A(n494), .ZN(
        n459) );
  INV_X1 U198 ( .A(R[21]), .ZN(n315) );
  INV_X1 U199 ( .A(n259), .ZN(n265) );
  OAI221_X1 U200 ( .B1(n377), .B2(n457), .C1(n378), .C2(n461), .A(n462), .ZN(
        n252) );
  INV_X1 U202 ( .A(R[15]), .ZN(n461) );
  AOI221_X1 U203 ( .B1(n270), .B2(n267), .C1(n259), .C2(n269), .A(n463), .ZN(
        n248) );
  OAI22_X1 U204 ( .A1(n262), .A2(n264), .B1(n251), .B2(n434), .ZN(n463) );
  OAI211_X1 U205 ( .C1(n378), .C2(n367), .A(n497), .B(n464), .ZN(n434) );
  AOI222_X1 U206 ( .A1(R[24]), .A2(n423), .B1(R[0]), .B2(n298), .C1(R[8]), 
        .C2(n299), .ZN(n464) );
  INV_X1 U208 ( .A(R[16]), .ZN(n367) );
  INV_X1 U209 ( .A(n268), .ZN(n251) );
  OAI221_X1 U210 ( .B1(n457), .B2(n411), .C1(n378), .C2(n354), .A(n465), .ZN(
        n264) );
  AOI221_X1 U211 ( .B1(R[18]), .B2(n423), .C1(R[2]), .C2(n299), .A(n494), .ZN(
        n465) );
  INV_X1 U213 ( .A(R[26]), .ZN(n411) );
  AOI221_X1 U214 ( .B1(n423), .B2(R[20]), .C1(n325), .C2(R[12]), .A(n466), 
        .ZN(n269) );
  OAI221_X1 U215 ( .B1(n335), .B2(n457), .C1(n467), .C2(n316), .A(n330), .ZN(
        n466) );
  INV_X1 U216 ( .A(R[4]), .ZN(n467) );
  AOI221_X1 U217 ( .B1(n423), .B2(R[22]), .C1(n325), .C2(R[14]), .A(n468), 
        .ZN(n267) );
  OAI221_X1 U218 ( .B1(n385), .B2(n457), .C1(n301), .C2(n316), .A(n330), .ZN(
        n468) );
  INV_X1 U220 ( .A(n305), .ZN(n340) );
  NAND2_X1 U221 ( .A1(R[31]), .A2(Conf[1]), .ZN(n305) );
  INV_X1 U222 ( .A(n299), .ZN(n316) );
  INV_X1 U223 ( .A(n470), .ZN(n371) );
  INV_X1 U224 ( .A(R[30]), .ZN(n385) );
  MUX2_X1 U225 ( .A(n471), .B(n401), .S(\finegrainsel[0] ), .Z(Shift_OUT[0])
         );
  AOI221_X1 U226 ( .B1(n270), .B2(n281), .C1(n268), .C2(n275), .A(n472), .ZN(
        n401) );
  INV_X1 U227 ( .A(n473), .ZN(n472) );
  AOI21_X1 U228 ( .B1(n321), .B2(n259), .A(n474), .ZN(n473) );
  AOI211_X1 U229 ( .C1(R[9]), .C2(n423), .A(n475), .B(n262), .ZN(n474) );
  OAI222_X1 U230 ( .A1(n378), .A2(n329), .B1(n457), .B2(n327), .C1(n476), .C2(
        n361), .ZN(n475) );
  INV_X1 U231 ( .A(R[25]), .ZN(n361) );
  INV_X1 U232 ( .A(R[17]), .ZN(n327) );
  INV_X1 U233 ( .A(R[1]), .ZN(n329) );
  AOI221_X1 U234 ( .B1(n325), .B2(R[3]), .C1(n423), .C2(R[11]), .A(n477), .ZN(
        n321) );
  OAI22_X1 U235 ( .A1(n347), .A2(n457), .B1(n346), .B2(n476), .ZN(n477) );
  INV_X1 U236 ( .A(R[27]), .ZN(n346) );
  INV_X1 U237 ( .A(R[19]), .ZN(n347) );
  AOI221_X1 U238 ( .B1(n325), .B2(R[7]), .C1(n423), .C2(R[15]), .A(n478), .ZN(
        n275) );
  OAI22_X1 U239 ( .A1(n428), .A2(n457), .B1(n476), .B2(n377), .ZN(n478) );
  INV_X1 U240 ( .A(R[31]), .ZN(n377) );
  INV_X1 U241 ( .A(R[23]), .ZN(n428) );
  OAI22_X1 U242 ( .A1(n319), .A2(n328), .B1(n317), .B2(n476), .ZN(n479) );
  INV_X1 U243 ( .A(R[29]), .ZN(n317) );
  INV_X1 U244 ( .A(R[13]), .ZN(n319) );
  OAI221_X1 U245 ( .B1(n480), .B2(n262), .C1(n287), .C2(n253), .A(n481), .ZN(
        n471) );
  AOI22_X1 U246 ( .A1(n259), .A2(n403), .B1(n268), .B2(n288), .ZN(n481) );
  OAI221_X1 U247 ( .B1(n328), .B2(n303), .C1(n378), .C2(n301), .A(n482), .ZN(
        n288) );
  AOI22_X1 U248 ( .A1(R[22]), .A2(n324), .B1(R[30]), .B2(n469), .ZN(n482) );
  INV_X1 U249 ( .A(R[6]), .ZN(n301) );
  INV_X1 U250 ( .A(R[14]), .ZN(n303) );
  OAI221_X1 U251 ( .B1(n355), .B2(n378), .C1(n328), .C2(n354), .A(n485), .ZN(
        n403) );
  AOI22_X1 U252 ( .A1(n324), .A2(R[18]), .B1(R[26]), .B2(n469), .ZN(n485) );
  INV_X1 U253 ( .A(R[10]), .ZN(n354) );
  INV_X1 U254 ( .A(n423), .ZN(n328) );
  INV_X1 U255 ( .A(R[2]), .ZN(n355) );
  INV_X1 U256 ( .A(n270), .ZN(n253) );
  INV_X1 U257 ( .A(n486), .ZN(n484) );
  AOI221_X1 U258 ( .B1(n325), .B2(R[4]), .C1(n423), .C2(R[12]), .A(n488), .ZN(
        n287) );
  OAI22_X1 U259 ( .A1(n336), .A2(n457), .B1(n335), .B2(n476), .ZN(n488) );
  INV_X1 U260 ( .A(R[28]), .ZN(n335) );
  INV_X1 U261 ( .A(n324), .ZN(n457) );
  INV_X1 U262 ( .A(R[20]), .ZN(n336) );
  INV_X1 U263 ( .A(n257), .ZN(n262) );
  INV_X1 U264 ( .A(n483), .ZN(n487) );
  NAND2_X1 U265 ( .A1(n489), .A2(n490), .ZN(n483) );
  MUX2_X1 U266 ( .A(n470), .B(n491), .S(Offset[1]), .Z(n489) );
  NAND2_X1 U267 ( .A1(\finegrainsel[0] ), .A2(n470), .ZN(n491) );
  XNOR2_X1 U268 ( .A(n492), .B(Offset[2]), .ZN(n486) );
  NAND2_X1 U269 ( .A1(n470), .A2(n490), .ZN(n492) );
  OR2_X1 U270 ( .A1(\finegrainsel[0] ), .A2(Offset[1]), .ZN(n490) );
  AOI221_X1 U271 ( .B1(R[8]), .B2(n423), .C1(R[16]), .C2(n324), .A(n493), .ZN(
        n480) );
  OAI22_X1 U272 ( .A1(n476), .A2(n368), .B1(n378), .B2(n406), .ZN(n493) );
  INV_X1 U273 ( .A(R[0]), .ZN(n406) );
  INV_X1 U274 ( .A(n325), .ZN(n378) );
  INV_X1 U275 ( .A(R[24]), .ZN(n368) );
  INV_X1 U276 ( .A(n469), .ZN(n476) );
  NOR3_X1 U277 ( .A1(n370), .A2(n470), .A3(n372), .ZN(n469) );
  INV_X1 U278 ( .A(Offset[4]), .ZN(n372) );
  INV_X1 U279 ( .A(Offset[3]), .ZN(n370) );
  NOR2_X1 U280 ( .A1(Conf[1]), .A2(Conf[0]), .ZN(n470) );
  OAI221_X1 U65 ( .B1(Offset[4]), .B2(Offset[3]), .C1(Conf[1]), .C2(Conf[0]), 
        .A(n340), .ZN(n379) );
  AND2_X2 U71 ( .A1(n469), .A2(n340), .ZN(n494) );
  INV_X4 U85 ( .A(n494), .ZN(n330) );
  AOI221_X4 U91 ( .B1(n338), .B2(R[9]), .C1(n339), .C2(R[1]), .A(n340), .ZN(
        n362) );
  AOI21_X1 U146 ( .B1(n340), .B2(n324), .A(n494), .ZN(n429) );
  INV_X1 U201 ( .A(n429), .ZN(n495) );
  INV_X1 U207 ( .A(n495), .ZN(n496) );
  INV_X1 U212 ( .A(n495), .ZN(n497) );
  AOI221_X4 U219 ( .B1(n338), .B2(R[12]), .C1(n339), .C2(R[4]), .A(n340), .ZN(
        n337) );
  AOI221_X4 U281 ( .B1(n338), .B2(R[11]), .C1(n339), .C2(R[3]), .A(n340), .ZN(
        n348) );
  AOI221_X4 U282 ( .B1(n338), .B2(R[8]), .C1(n339), .C2(R[0]), .A(n340), .ZN(
        n369) );
  AOI221_X4 U283 ( .B1(R[23]), .B2(n423), .C1(R[7]), .C2(n299), .A(n494), .ZN(
        n462) );
endmodule


module ComparatorUnit ( A_MSB, B_MSB, SUBIN, COUT, SIGN_UNSIGN, .OP({\OP[2] , 
        \OP[1] , \OP[0] }), CU_OUT );
  input [31:0] SUBIN;
  output [31:0] CU_OUT;
  input A_MSB, B_MSB, COUT, SIGN_UNSIGN, \OP[2] , \OP[1] , \OP[0] ;
  wire   net123593, n39, n50, n41, n40, net124999, net124998, net124924,
         net124922, net125054, net125029, net125028, net125025, net125024,
         net125023, net125022, net125021, net124992, net124989, net124976,
         net124927, n34, n32, n30, net125020, net124983, net124980, net124995,
         net125095, net125050, net124982, net124967, net124965, net124964,
         net124963, net124925, net123651, net123650, net123620, net123618, n36,
         n31, net125090, net125007, net125006, net125005, net125004, net125002,
         net124994, net124993, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81;
  assign CU_OUT[31] = 1'b0;
  assign CU_OUT[30] = 1'b0;
  assign CU_OUT[29] = 1'b0;
  assign CU_OUT[28] = 1'b0;
  assign CU_OUT[27] = 1'b0;
  assign CU_OUT[26] = 1'b0;
  assign CU_OUT[25] = 1'b0;
  assign CU_OUT[24] = 1'b0;
  assign CU_OUT[23] = 1'b0;
  assign CU_OUT[22] = 1'b0;
  assign CU_OUT[21] = 1'b0;
  assign CU_OUT[20] = 1'b0;
  assign CU_OUT[19] = 1'b0;
  assign CU_OUT[18] = 1'b0;
  assign CU_OUT[17] = 1'b0;
  assign CU_OUT[16] = 1'b0;
  assign CU_OUT[15] = 1'b0;
  assign CU_OUT[14] = 1'b0;
  assign CU_OUT[13] = 1'b0;
  assign CU_OUT[12] = 1'b0;
  assign CU_OUT[11] = 1'b0;
  assign CU_OUT[10] = 1'b0;
  assign CU_OUT[9] = 1'b0;
  assign CU_OUT[8] = 1'b0;
  assign CU_OUT[7] = 1'b0;
  assign CU_OUT[6] = 1'b0;
  assign CU_OUT[5] = 1'b0;
  assign CU_OUT[4] = 1'b0;
  assign CU_OUT[3] = 1'b0;
  assign CU_OUT[2] = 1'b0;
  assign CU_OUT[1] = 1'b0;

  INV_X1 U67 ( .A(A_MSB), .ZN(n40) );
  XOR2_X1 U76 ( .A(B_MSB), .B(A_MSB), .Z(n50) );
  AND2_X1 U75 ( .A1(SIGN_UNSIGN), .A2(n50), .ZN(n41) );
  INV_X2 syn379 ( .A(n40), .ZN(net124999) );
  NAND3_X1 syn369 ( .A1(n80), .A2(net125028), .A3(net124989), .ZN(n81) );
  NOR2_X2 syn362 ( .A1(net125022), .A2(net125023), .ZN(n79) );
  OAI21_X1 U63 ( .B1(net123593), .B2(n39), .A(n34), .ZN(n30) );
  NAND2_X2 syn489 ( .A1(OP[0]), .A2(net125029), .ZN(net124922) );
  NAND3_X1 syn361 ( .A1(net125024), .A2(net125025), .A3(n71), .ZN(net125023)
         );
  INV_X1 U64 ( .A(OP[1]), .ZN(n34) );
  INV_X2 syn92 ( .A(OP[0]), .ZN(net124925) );
  AOI22_X1 U58 ( .A1(n30), .A2(OP[2]), .B1(n31), .B2(n32), .ZN(CU_OUT[0]) );
  NAND3_X1 syn309 ( .A1(net125004), .A2(net125005), .A3(net125007), .ZN(
        net125006) );
  NOR2_X2 syn294 ( .A1(n41), .A2(SUBIN[1]), .ZN(n60) );
  INV_X2 syn411 ( .A(SUBIN[15]), .ZN(n62) );
  NOR2_X2 syn312 ( .A1(SUBIN[0]), .A2(SUBIN[10]), .ZN(n63) );
  NOR2_X2 syn316 ( .A1(SUBIN[4]), .A2(SUBIN[9]), .ZN(n64) );
  NAND3_X1 syn319 ( .A1(n63), .A2(n66), .A3(n64), .ZN(n65) );
  NOR2_X2 syn320 ( .A1(SUBIN[8]), .A2(SUBIN[5]), .ZN(n67) );
  NOR2_X2 syn324 ( .A1(SUBIN[6]), .A2(SUBIN[2]), .ZN(n68) );
  NAND3_X1 syn327 ( .A1(n67), .A2(n70), .A3(n68), .ZN(n69) );
  NAND2_X1 U59 ( .A1(net124983), .A2(net124964), .ZN(n74) );
  OR2_X1 U60 ( .A1(SUBIN[25]), .A2(SUBIN[26]), .ZN(net124983) );
  CLKBUF_X1 U61 ( .A(n72), .Z(n53) );
  AND4_X1 U62 ( .A1(n58), .A2(n59), .A3(net125090), .A4(net124993), .ZN(n54)
         );
  NAND2_X1 U65 ( .A1(net125021), .A2(n53), .ZN(net125022) );
  OAI21_X1 U66 ( .B1(net125029), .B2(n34), .A(OP[0]), .ZN(net124976) );
  AND4_X1 U68 ( .A1(net124989), .A2(n72), .A3(n55), .A4(n56), .ZN(net125020)
         );
  INV_X1 U69 ( .A(SUBIN[25]), .ZN(n55) );
  INV_X1 U70 ( .A(SUBIN[26]), .ZN(n56) );
  OAI211_X1 U71 ( .C1(net125095), .C2(net123650), .A(n73), .B(n74), .ZN(
        net124965) );
  NOR2_X1 U72 ( .A1(net124963), .A2(net124967), .ZN(net123593) );
  NOR2_X1 U73 ( .A1(n81), .A2(net124992), .ZN(n78) );
  OAI211_X1 U74 ( .C1(n54), .C2(net123650), .A(n57), .B(net123620), .ZN(n31)
         );
  INV_X1 U77 ( .A(net124965), .ZN(n57) );
  NAND4_X1 U78 ( .A1(n58), .A2(n59), .A3(net124994), .A4(net124993), .ZN(
        net124963) );
  INV_X1 U79 ( .A(net124995), .ZN(n58) );
  INV_X1 U80 ( .A(OP[0]), .ZN(n59) );
  NOR2_X1 U81 ( .A1(net125002), .A2(net125006), .ZN(net124994) );
  NOR2_X1 U82 ( .A1(n65), .A2(n69), .ZN(net124993) );
  NAND2_X1 U83 ( .A1(net125090), .A2(net124993), .ZN(net124992) );
  INV_X1 U84 ( .A(SUBIN[7]), .ZN(n70) );
  INV_X1 U85 ( .A(SUBIN[11]), .ZN(n66) );
  NAND3_X1 U86 ( .A1(n60), .A2(n62), .A3(n61), .ZN(net125002) );
  NOR2_X1 U87 ( .A1(net125002), .A2(net125006), .ZN(net125090) );
  NOR2_X1 U88 ( .A1(SUBIN[14]), .A2(SUBIN[13]), .ZN(n61) );
  INV_X1 U89 ( .A(SUBIN[12]), .ZN(net125007) );
  NOR2_X1 U90 ( .A1(SUBIN[17]), .A2(SUBIN[16]), .ZN(net125005) );
  NOR2_X1 U91 ( .A1(SUBIN[18]), .A2(SUBIN[19]), .ZN(net125004) );
  MUX2_X2 U92 ( .A(net124998), .B(net124999), .S(n41), .Z(net124924) );
  NAND2_X1 U93 ( .A1(n36), .A2(OP[1]), .ZN(net123620) );
  AND2_X1 U94 ( .A1(net125050), .A2(n75), .ZN(n73) );
  NAND2_X1 U95 ( .A1(net124964), .A2(SUBIN[27]), .ZN(n75) );
  INV_X1 U96 ( .A(net123650), .ZN(net124964) );
  OR2_X1 U97 ( .A1(n72), .A2(net123650), .ZN(net125050) );
  INV_X1 U98 ( .A(SUBIN[24]), .ZN(n72) );
  NAND2_X1 U99 ( .A1(net124924), .A2(net124925), .ZN(n36) );
  NAND2_X1 U100 ( .A1(n36), .A2(net124922), .ZN(n39) );
  INV_X1 U101 ( .A(OP[1]), .ZN(net123618) );
  OR2_X1 U102 ( .A1(OP[2]), .A2(net123651), .ZN(net123650) );
  INV_X1 U103 ( .A(net123618), .ZN(net123651) );
  AND3_X1 U104 ( .A1(net124980), .A2(net124982), .A3(n71), .ZN(net125095) );
  NAND2_X1 U105 ( .A1(net125020), .A2(net125095), .ZN(net124967) );
  INV_X1 U106 ( .A(SUBIN[23]), .ZN(n71) );
  NOR2_X1 U107 ( .A1(SUBIN[29]), .A2(SUBIN[28]), .ZN(net124982) );
  NAND2_X1 U108 ( .A1(n76), .A2(n77), .ZN(net124995) );
  INV_X1 U109 ( .A(net124995), .ZN(net125028) );
  NOR2_X1 U110 ( .A1(SUBIN[22]), .A2(SUBIN[21]), .ZN(n77) );
  NOR2_X2 U111 ( .A1(SUBIN[20]), .A2(SUBIN[3]), .ZN(n76) );
  NOR2_X1 U112 ( .A1(SUBIN[30]), .A2(SUBIN[31]), .ZN(net124980) );
  INV_X1 U113 ( .A(SUBIN[27]), .ZN(net124989) );
  INV_X1 U114 ( .A(net124927), .ZN(n32) );
  AOI21_X1 U115 ( .B1(n78), .B2(n79), .A(net124976), .ZN(net124927) );
  INV_X1 U116 ( .A(net124924), .ZN(net125029) );
  INV_X1 U117 ( .A(SUBIN[30]), .ZN(net125025) );
  INV_X1 U118 ( .A(SUBIN[31]), .ZN(net125024) );
  NOR2_X1 U119 ( .A1(net125054), .A2(SUBIN[25]), .ZN(net125021) );
  CLKBUF_X1 U120 ( .A(SUBIN[26]), .Z(net125054) );
  NOR2_X1 U121 ( .A1(SUBIN[29]), .A2(SUBIN[28]), .ZN(n80) );
  INV_X1 U122 ( .A(COUT), .ZN(net124998) );
endmodule


module logicunit ( A, B, SEL, LU_OUT );
  input [31:0] A;
  input [31:0] B;
  input [2:0] SEL;
  output [31:0] LU_OUT;
  wire   n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128;

  MUX2_X1 U1 ( .A(n65), .B(n66), .S(B[9]), .Z(LU_OUT[9]) );
  MUX2_X1 U2 ( .A(SEL[0]), .B(SEL[2]), .S(A[9]), .Z(n66) );
  AND2_X1 U3 ( .A1(A[9]), .A2(SEL[1]), .ZN(n65) );
  MUX2_X1 U4 ( .A(n67), .B(n68), .S(B[8]), .Z(LU_OUT[8]) );
  MUX2_X1 U5 ( .A(SEL[0]), .B(SEL[2]), .S(A[8]), .Z(n68) );
  AND2_X1 U6 ( .A1(SEL[1]), .A2(A[8]), .ZN(n67) );
  MUX2_X1 U7 ( .A(n69), .B(n70), .S(B[7]), .Z(LU_OUT[7]) );
  MUX2_X1 U8 ( .A(SEL[0]), .B(SEL[2]), .S(A[7]), .Z(n70) );
  AND2_X1 U9 ( .A1(SEL[1]), .A2(A[7]), .ZN(n69) );
  MUX2_X1 U10 ( .A(n71), .B(n72), .S(B[6]), .Z(LU_OUT[6]) );
  MUX2_X1 U11 ( .A(SEL[0]), .B(SEL[2]), .S(A[6]), .Z(n72) );
  AND2_X1 U12 ( .A1(SEL[1]), .A2(A[6]), .ZN(n71) );
  MUX2_X1 U13 ( .A(n73), .B(n74), .S(B[5]), .Z(LU_OUT[5]) );
  MUX2_X1 U14 ( .A(SEL[0]), .B(SEL[2]), .S(A[5]), .Z(n74) );
  AND2_X1 U15 ( .A1(SEL[1]), .A2(A[5]), .ZN(n73) );
  MUX2_X1 U16 ( .A(n75), .B(n76), .S(B[4]), .Z(LU_OUT[4]) );
  MUX2_X1 U17 ( .A(SEL[0]), .B(SEL[2]), .S(A[4]), .Z(n76) );
  AND2_X1 U18 ( .A1(SEL[1]), .A2(A[4]), .ZN(n75) );
  MUX2_X1 U19 ( .A(n77), .B(n78), .S(B[3]), .Z(LU_OUT[3]) );
  MUX2_X1 U20 ( .A(SEL[0]), .B(SEL[2]), .S(A[3]), .Z(n78) );
  AND2_X1 U21 ( .A1(SEL[1]), .A2(A[3]), .ZN(n77) );
  MUX2_X1 U22 ( .A(n79), .B(n80), .S(B[31]), .Z(LU_OUT[31]) );
  MUX2_X1 U23 ( .A(SEL[0]), .B(SEL[2]), .S(A[31]), .Z(n80) );
  AND2_X1 U24 ( .A1(SEL[1]), .A2(A[31]), .ZN(n79) );
  MUX2_X1 U25 ( .A(n81), .B(n82), .S(B[30]), .Z(LU_OUT[30]) );
  MUX2_X1 U26 ( .A(SEL[0]), .B(SEL[2]), .S(A[30]), .Z(n82) );
  AND2_X1 U27 ( .A1(SEL[1]), .A2(A[30]), .ZN(n81) );
  MUX2_X1 U28 ( .A(n83), .B(n84), .S(B[2]), .Z(LU_OUT[2]) );
  MUX2_X1 U29 ( .A(SEL[0]), .B(SEL[2]), .S(A[2]), .Z(n84) );
  AND2_X1 U30 ( .A1(SEL[1]), .A2(A[2]), .ZN(n83) );
  MUX2_X1 U31 ( .A(n85), .B(n86), .S(B[29]), .Z(LU_OUT[29]) );
  MUX2_X1 U32 ( .A(SEL[0]), .B(SEL[2]), .S(A[29]), .Z(n86) );
  AND2_X1 U33 ( .A1(SEL[1]), .A2(A[29]), .ZN(n85) );
  MUX2_X1 U34 ( .A(n87), .B(n88), .S(B[28]), .Z(LU_OUT[28]) );
  MUX2_X1 U35 ( .A(SEL[0]), .B(SEL[2]), .S(A[28]), .Z(n88) );
  AND2_X1 U36 ( .A1(SEL[1]), .A2(A[28]), .ZN(n87) );
  MUX2_X1 U37 ( .A(n89), .B(n90), .S(B[27]), .Z(LU_OUT[27]) );
  MUX2_X1 U38 ( .A(SEL[0]), .B(SEL[2]), .S(A[27]), .Z(n90) );
  AND2_X1 U39 ( .A1(SEL[1]), .A2(A[27]), .ZN(n89) );
  MUX2_X1 U40 ( .A(n91), .B(n92), .S(B[26]), .Z(LU_OUT[26]) );
  MUX2_X1 U41 ( .A(SEL[0]), .B(SEL[2]), .S(A[26]), .Z(n92) );
  AND2_X1 U42 ( .A1(SEL[1]), .A2(A[26]), .ZN(n91) );
  MUX2_X1 U43 ( .A(n93), .B(n94), .S(B[25]), .Z(LU_OUT[25]) );
  MUX2_X1 U44 ( .A(SEL[0]), .B(SEL[2]), .S(A[25]), .Z(n94) );
  AND2_X1 U45 ( .A1(SEL[1]), .A2(A[25]), .ZN(n93) );
  MUX2_X1 U46 ( .A(n95), .B(n96), .S(B[24]), .Z(LU_OUT[24]) );
  MUX2_X1 U47 ( .A(SEL[0]), .B(SEL[2]), .S(A[24]), .Z(n96) );
  AND2_X1 U48 ( .A1(SEL[1]), .A2(A[24]), .ZN(n95) );
  MUX2_X1 U49 ( .A(n97), .B(n98), .S(B[23]), .Z(LU_OUT[23]) );
  MUX2_X1 U50 ( .A(SEL[0]), .B(SEL[2]), .S(A[23]), .Z(n98) );
  AND2_X1 U51 ( .A1(SEL[1]), .A2(A[23]), .ZN(n97) );
  MUX2_X1 U52 ( .A(n99), .B(n100), .S(B[22]), .Z(LU_OUT[22]) );
  MUX2_X1 U53 ( .A(SEL[0]), .B(SEL[2]), .S(A[22]), .Z(n100) );
  AND2_X1 U54 ( .A1(SEL[1]), .A2(A[22]), .ZN(n99) );
  MUX2_X1 U55 ( .A(n101), .B(n102), .S(B[21]), .Z(LU_OUT[21]) );
  MUX2_X1 U56 ( .A(SEL[0]), .B(SEL[2]), .S(A[21]), .Z(n102) );
  AND2_X1 U57 ( .A1(SEL[1]), .A2(A[21]), .ZN(n101) );
  MUX2_X1 U58 ( .A(n103), .B(n104), .S(B[20]), .Z(LU_OUT[20]) );
  MUX2_X1 U59 ( .A(SEL[0]), .B(SEL[2]), .S(A[20]), .Z(n104) );
  AND2_X1 U60 ( .A1(SEL[1]), .A2(A[20]), .ZN(n103) );
  MUX2_X1 U61 ( .A(n105), .B(n106), .S(B[1]), .Z(LU_OUT[1]) );
  MUX2_X1 U62 ( .A(SEL[0]), .B(SEL[2]), .S(A[1]), .Z(n106) );
  AND2_X1 U63 ( .A1(SEL[1]), .A2(A[1]), .ZN(n105) );
  MUX2_X1 U64 ( .A(n107), .B(n108), .S(B[19]), .Z(LU_OUT[19]) );
  MUX2_X1 U65 ( .A(SEL[0]), .B(SEL[2]), .S(A[19]), .Z(n108) );
  AND2_X1 U66 ( .A1(SEL[1]), .A2(A[19]), .ZN(n107) );
  MUX2_X1 U67 ( .A(n109), .B(n110), .S(B[18]), .Z(LU_OUT[18]) );
  MUX2_X1 U68 ( .A(SEL[0]), .B(SEL[2]), .S(A[18]), .Z(n110) );
  AND2_X1 U69 ( .A1(SEL[1]), .A2(A[18]), .ZN(n109) );
  MUX2_X1 U70 ( .A(n111), .B(n112), .S(B[17]), .Z(LU_OUT[17]) );
  MUX2_X1 U71 ( .A(SEL[0]), .B(SEL[2]), .S(A[17]), .Z(n112) );
  AND2_X1 U72 ( .A1(SEL[1]), .A2(A[17]), .ZN(n111) );
  MUX2_X1 U73 ( .A(n113), .B(n114), .S(B[16]), .Z(LU_OUT[16]) );
  MUX2_X1 U74 ( .A(SEL[0]), .B(SEL[2]), .S(A[16]), .Z(n114) );
  AND2_X1 U75 ( .A1(SEL[1]), .A2(A[16]), .ZN(n113) );
  MUX2_X1 U76 ( .A(n115), .B(n116), .S(B[15]), .Z(LU_OUT[15]) );
  MUX2_X1 U77 ( .A(SEL[0]), .B(SEL[2]), .S(A[15]), .Z(n116) );
  AND2_X1 U78 ( .A1(SEL[1]), .A2(A[15]), .ZN(n115) );
  MUX2_X1 U79 ( .A(n117), .B(n118), .S(B[14]), .Z(LU_OUT[14]) );
  MUX2_X1 U80 ( .A(SEL[0]), .B(SEL[2]), .S(A[14]), .Z(n118) );
  AND2_X1 U81 ( .A1(SEL[1]), .A2(A[14]), .ZN(n117) );
  MUX2_X1 U82 ( .A(n119), .B(n120), .S(B[13]), .Z(LU_OUT[13]) );
  MUX2_X1 U83 ( .A(SEL[0]), .B(SEL[2]), .S(A[13]), .Z(n120) );
  AND2_X1 U84 ( .A1(SEL[1]), .A2(A[13]), .ZN(n119) );
  MUX2_X1 U85 ( .A(n121), .B(n122), .S(B[12]), .Z(LU_OUT[12]) );
  MUX2_X1 U86 ( .A(SEL[0]), .B(SEL[2]), .S(A[12]), .Z(n122) );
  AND2_X1 U87 ( .A1(SEL[1]), .A2(A[12]), .ZN(n121) );
  MUX2_X1 U88 ( .A(n123), .B(n124), .S(B[11]), .Z(LU_OUT[11]) );
  MUX2_X1 U89 ( .A(SEL[0]), .B(SEL[2]), .S(A[11]), .Z(n124) );
  AND2_X1 U90 ( .A1(SEL[1]), .A2(A[11]), .ZN(n123) );
  MUX2_X1 U91 ( .A(n125), .B(n126), .S(B[10]), .Z(LU_OUT[10]) );
  MUX2_X1 U92 ( .A(SEL[0]), .B(SEL[2]), .S(A[10]), .Z(n126) );
  AND2_X1 U93 ( .A1(SEL[1]), .A2(A[10]), .ZN(n125) );
  MUX2_X1 U94 ( .A(n127), .B(n128), .S(B[0]), .Z(LU_OUT[0]) );
  MUX2_X1 U95 ( .A(SEL[0]), .B(SEL[2]), .S(A[0]), .Z(n128) );
  AND2_X1 U96 ( .A1(SEL[1]), .A2(A[0]), .ZN(n127) );
endmodule


module sumgen_N_blocks8 ( A, B, Ci, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] Ci;
  output [31:0] S;


  CSB_0 CSBI_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(S[3:0]) );
  CSB_7 CSBI_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(S[7:4]) );
  CSB_6 CSBI_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), .S(S[11:8]) );
  CSB_5 CSBI_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), .S(S[15:12]) );
  CSB_4 CSBI_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), .S(S[19:16]) );
  CSB_3 CSBI_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), .S(S[23:20]) );
  CSB_2 CSBI_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), .S(S[27:24]) );
  CSB_1 CSBI_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), .S(S[31:28]) );
endmodule


module STCG_N32_L5 ( A, B, cin, cout );
  input [31:0] A;
  input [31:0] B;
  output [7:0] cout;
  input cin;
  wire   \gen[0][31] , \gen[0][30] , \gen[0][29] , \gen[0][28] , \gen[0][27] ,
         \gen[0][26] , \gen[0][25] , \gen[0][24] , \gen[0][23] , \gen[0][22] ,
         \gen[0][21] , \gen[0][20] , \gen[0][19] , \gen[0][18] , \gen[0][17] ,
         \gen[0][16] , \gen[0][15] , \gen[0][14] , \gen[0][13] , \gen[0][12] ,
         \gen[0][11] , \gen[0][10] , \gen[0][9] , \gen[0][8] , \gen[0][7] ,
         \gen[0][6] , \gen[0][5] , \gen[0][4] , \gen[0][3] , \gen[0][2] ,
         \gen[0][1] , \gen[0][0] , \gen[1][31] , \gen[1][29] , \gen[1][27] ,
         \gen[1][25] , \gen[1][23] , \gen[1][21] , \gen[1][19] , \gen[1][17] ,
         \gen[1][15] , \gen[1][13] , \gen[1][11] , \gen[1][9] , \gen[1][7] ,
         \gen[1][5] , \gen[1][3] , \gen[1][1] , \gen[2][31] , \gen[2][23] ,
         \gen[2][15] , \gen[2][7] , \gen[3][31] , \gen[3][15] , \gen[4][31] ,
         \gen[4][27] , \prop[0][31] , \prop[0][30] , \prop[0][29] ,
         \prop[0][28] , \prop[0][27] , \prop[0][26] , \prop[0][25] ,
         \prop[0][24] , \prop[0][23] , \prop[0][22] , \prop[0][21] ,
         \prop[0][20] , \prop[0][19] , \prop[0][18] , \prop[0][17] ,
         \prop[0][16] , \prop[0][15] , \prop[0][14] , \prop[0][13] ,
         \prop[0][12] , \prop[0][11] , \prop[0][10] , \prop[0][9] ,
         \prop[0][8] , \prop[0][7] , \prop[0][6] , \prop[0][5] , \prop[0][4] ,
         \prop[0][3] , \prop[0][2] , \prop[0][1] , \prop[1][31] ,
         \prop[1][29] , \prop[1][27] , \prop[1][25] , \prop[1][23] ,
         \prop[1][21] , \prop[1][19] , \prop[1][17] , \prop[1][15] ,
         \prop[1][13] , \prop[1][11] , \prop[1][9] , \prop[1][7] ,
         \prop[1][5] , \prop[1][3] , \prop[2][31] , \prop[2][27] ,
         \prop[2][23] , \prop[2][19] , \prop[2][15] , \prop[2][11] ,
         \prop[2][7] , \prop[3][31] , \prop[3][23] , \prop[3][15] ,
         \prop[4][31] , \prop[4][27] , n1, n22, n23, n24, n37, n26, n36, n29,
         n30, n32, n33;

  prop_gen_Cin prop_gen_Cin0 ( .a(A[0]), .b(B[0]), .cin(cin), .gen(\gen[0][0] ) );
  prop_gen_0 prop_gen_i_1 ( .a(A[1]), .b(B[1]), .prop(\prop[0][1] ), .gen(
        \gen[0][1] ) );
  prop_gen_30 prop_gen_i_2 ( .a(A[2]), .b(B[2]), .prop(\prop[0][2] ), .gen(
        \gen[0][2] ) );
  prop_gen_29 prop_gen_i_3 ( .a(A[3]), .b(B[3]), .prop(\prop[0][3] ), .gen(
        \gen[0][3] ) );
  prop_gen_28 prop_gen_i_4 ( .a(A[4]), .b(B[4]), .prop(\prop[0][4] ), .gen(
        \gen[0][4] ) );
  prop_gen_27 prop_gen_i_5 ( .a(A[5]), .b(B[5]), .prop(\prop[0][5] ), .gen(
        \gen[0][5] ) );
  prop_gen_26 prop_gen_i_6 ( .a(A[6]), .b(B[6]), .prop(\prop[0][6] ), .gen(
        \gen[0][6] ) );
  prop_gen_25 prop_gen_i_7 ( .a(A[7]), .b(B[7]), .prop(\prop[0][7] ), .gen(
        \gen[0][7] ) );
  prop_gen_24 prop_gen_i_8 ( .a(A[8]), .b(B[8]), .prop(\prop[0][8] ), .gen(
        \gen[0][8] ) );
  prop_gen_23 prop_gen_i_9 ( .a(A[9]), .b(B[9]), .prop(\prop[0][9] ), .gen(
        \gen[0][9] ) );
  prop_gen_22 prop_gen_i_10 ( .a(A[10]), .b(B[10]), .prop(\prop[0][10] ), 
        .gen(\gen[0][10] ) );
  prop_gen_21 prop_gen_i_11 ( .a(A[11]), .b(B[11]), .prop(\prop[0][11] ), 
        .gen(\gen[0][11] ) );
  prop_gen_20 prop_gen_i_12 ( .a(A[12]), .b(B[12]), .prop(\prop[0][12] ), 
        .gen(\gen[0][12] ) );
  prop_gen_19 prop_gen_i_13 ( .a(A[13]), .b(B[13]), .prop(\prop[0][13] ), 
        .gen(\gen[0][13] ) );
  prop_gen_18 prop_gen_i_14 ( .a(A[14]), .b(B[14]), .prop(\prop[0][14] ), 
        .gen(\gen[0][14] ) );
  prop_gen_17 prop_gen_i_15 ( .a(A[15]), .b(B[15]), .prop(\prop[0][15] ), 
        .gen(\gen[0][15] ) );
  prop_gen_16 prop_gen_i_16 ( .a(A[16]), .b(B[16]), .prop(\prop[0][16] ), 
        .gen(\gen[0][16] ) );
  prop_gen_15 prop_gen_i_17 ( .a(A[17]), .b(B[17]), .prop(\prop[0][17] ), 
        .gen(\gen[0][17] ) );
  prop_gen_14 prop_gen_i_18 ( .a(A[18]), .b(B[18]), .prop(\prop[0][18] ), 
        .gen(\gen[0][18] ) );
  prop_gen_13 prop_gen_i_19 ( .a(A[19]), .b(B[19]), .prop(\prop[0][19] ), 
        .gen(\gen[0][19] ) );
  prop_gen_12 prop_gen_i_20 ( .a(A[20]), .b(B[20]), .prop(\prop[0][20] ), 
        .gen(\gen[0][20] ) );
  prop_gen_11 prop_gen_i_21 ( .a(A[21]), .b(B[21]), .prop(\prop[0][21] ), 
        .gen(\gen[0][21] ) );
  prop_gen_10 prop_gen_i_22 ( .a(A[22]), .b(B[22]), .prop(\prop[0][22] ), 
        .gen(\gen[0][22] ) );
  prop_gen_9 prop_gen_i_23 ( .a(A[23]), .b(B[23]), .prop(\prop[0][23] ), .gen(
        \gen[0][23] ) );
  prop_gen_8 prop_gen_i_24 ( .a(A[24]), .b(B[24]), .prop(\prop[0][24] ), .gen(
        \gen[0][24] ) );
  prop_gen_7 prop_gen_i_25 ( .a(A[25]), .b(B[25]), .prop(\prop[0][25] ), .gen(
        \gen[0][25] ) );
  prop_gen_6 prop_gen_i_26 ( .a(A[26]), .b(B[26]), .prop(\prop[0][26] ), .gen(
        \gen[0][26] ) );
  prop_gen_5 prop_gen_i_27 ( .a(A[27]), .b(B[27]), .prop(\prop[0][27] ), .gen(
        \gen[0][27] ) );
  prop_gen_4 prop_gen_i_28 ( .a(A[28]), .b(B[28]), .prop(\prop[0][28] ), .gen(
        \gen[0][28] ) );
  prop_gen_3 prop_gen_i_29 ( .a(A[29]), .b(B[29]), .prop(\prop[0][29] ), .gen(
        \gen[0][29] ) );
  prop_gen_2 prop_gen_i_30 ( .a(A[30]), .b(B[30]), .prop(\prop[0][30] ), .gen(
        \gen[0][30] ) );
  prop_gen_1 prop_gen_i_31 ( .a(A[31]), .b(B[31]), .prop(\prop[0][31] ), .gen(
        \gen[0][31] ) );
  G_0 G_1_1_1 ( .pi(\prop[0][1] ), .gi(\gen[0][1] ), .gj(\gen[0][0] ), .gout(
        \gen[1][1] ) );
  PG_0 PG_0_i_1_3 ( .pi(\prop[0][3] ), .gi(\gen[0][3] ), .pj(\prop[0][2] ), 
        .gj(\gen[0][2] ), .pout(\prop[1][3] ), .gout(\gen[1][3] ) );
  PG_26 PG_0_i_1_5 ( .pi(\prop[0][5] ), .gi(\gen[0][5] ), .pj(\prop[0][4] ), 
        .gj(\gen[0][4] ), .pout(\prop[1][5] ), .gout(\gen[1][5] ) );
  PG_25 PG_0_i_1_7 ( .pi(\prop[0][7] ), .gi(\gen[0][7] ), .pj(\prop[0][6] ), 
        .gj(\gen[0][6] ), .pout(\prop[1][7] ), .gout(\gen[1][7] ) );
  PG_24 PG_0_i_1_9 ( .pi(\prop[0][9] ), .gi(\gen[0][9] ), .pj(\prop[0][8] ), 
        .gj(\gen[0][8] ), .pout(\prop[1][9] ), .gout(\gen[1][9] ) );
  PG_23 PG_0_i_1_11 ( .pi(\prop[0][11] ), .gi(\gen[0][11] ), .pj(\prop[0][10] ), .gj(\gen[0][10] ), .pout(\prop[1][11] ), .gout(\gen[1][11] ) );
  PG_22 PG_0_i_1_13 ( .pi(\prop[0][13] ), .gi(\gen[0][13] ), .pj(\prop[0][12] ), .gj(\gen[0][12] ), .pout(\prop[1][13] ), .gout(\gen[1][13] ) );
  PG_21 PG_0_i_1_15 ( .pi(\prop[0][15] ), .gi(\gen[0][15] ), .pj(\prop[0][14] ), .gj(\gen[0][14] ), .pout(\prop[1][15] ), .gout(\gen[1][15] ) );
  PG_20 PG_0_i_1_17 ( .pi(\prop[0][17] ), .gi(\gen[0][17] ), .pj(\prop[0][16] ), .gj(\gen[0][16] ), .pout(\prop[1][17] ), .gout(\gen[1][17] ) );
  PG_19 PG_0_i_1_19 ( .pi(\prop[0][19] ), .gi(\gen[0][19] ), .pj(\prop[0][18] ), .gj(\gen[0][18] ), .pout(\prop[1][19] ), .gout(\gen[1][19] ) );
  PG_18 PG_0_i_1_21 ( .pi(\prop[0][21] ), .gi(\gen[0][21] ), .pj(\prop[0][20] ), .gj(\gen[0][20] ), .pout(\prop[1][21] ), .gout(\gen[1][21] ) );
  PG_17 PG_0_i_1_23 ( .pi(\prop[0][23] ), .gi(\gen[0][23] ), .pj(\prop[0][22] ), .gj(\gen[0][22] ), .pout(\prop[1][23] ), .gout(\gen[1][23] ) );
  PG_16 PG_0_i_1_25 ( .pi(\prop[0][25] ), .gi(\gen[0][25] ), .pj(\prop[0][24] ), .gj(\gen[0][24] ), .pout(\prop[1][25] ), .gout(\gen[1][25] ) );
  PG_15 PG_0_i_1_27 ( .pi(\prop[0][27] ), .gi(\gen[0][27] ), .pj(\prop[0][26] ), .gj(\gen[0][26] ), .pout(\prop[1][27] ), .gout(\gen[1][27] ) );
  PG_14 PG_0_i_1_29 ( .pi(\prop[0][29] ), .gi(\gen[0][29] ), .pj(\prop[0][28] ), .gj(\gen[0][28] ), .pout(\prop[1][29] ), .gout(\gen[1][29] ) );
  PG_13 PG_0_i_1_31 ( .pi(\prop[0][31] ), .gi(\gen[0][31] ), .pj(\prop[0][30] ), .gj(\gen[0][30] ), .pout(\prop[1][31] ), .gout(\gen[1][31] ) );
  G_8 G_23_2_3 ( .pi(\prop[1][3] ), .gi(\gen[1][3] ), .gj(\gen[1][1] ), .gout(
        n37) );
  PG_12 PG_0_i_2_7 ( .pi(\prop[1][7] ), .gi(\gen[1][7] ), .pj(\prop[1][5] ), 
        .gj(\gen[1][5] ), .pout(\prop[2][7] ), .gout(\gen[2][7] ) );
  PG_11 PG_0_i_2_11 ( .pi(\prop[1][11] ), .gi(\gen[1][11] ), .pj(\prop[1][9] ), 
        .gj(\gen[1][9] ), .pout(\prop[2][11] ), .gout(n24) );
  PG_10 PG_0_i_2_15 ( .pi(\prop[1][15] ), .gi(\gen[1][15] ), .pj(\prop[1][13] ), .gj(\gen[1][13] ), .pout(\prop[2][15] ), .gout(\gen[2][15] ) );
  PG_9 PG_0_i_2_19 ( .pi(\prop[1][19] ), .gi(\gen[1][19] ), .pj(\prop[1][17] ), 
        .gj(\gen[1][17] ), .pout(\prop[2][19] ), .gout(n22) );
  PG_8 PG_0_i_2_23 ( .pi(\prop[1][23] ), .gi(\gen[1][23] ), .pj(\prop[1][21] ), 
        .gj(\gen[1][21] ), .pout(\prop[2][23] ), .gout(\gen[2][23] ) );
  PG_7 PG_0_i_2_27 ( .pi(\prop[1][27] ), .gi(\gen[1][27] ), .pj(\prop[1][25] ), 
        .gj(\gen[1][25] ), .pout(\prop[2][27] ), .gout(n1) );
  PG_6 PG_0_i_2_31 ( .pi(\prop[1][31] ), .gi(\gen[1][31] ), .pj(\prop[1][29] ), 
        .gj(\gen[1][29] ), .pout(\prop[2][31] ), .gout(\gen[2][31] ) );
  G_7 G_23_3_7 ( .pi(\prop[2][7] ), .gi(\gen[2][7] ), .gj(n37), .gout(n26) );
  PG_5 PG_0_i_3_15 ( .pi(\prop[2][15] ), .gi(\gen[2][15] ), .pj(\prop[2][11] ), 
        .gj(n24), .pout(\prop[3][15] ), .gout(\gen[3][15] ) );
  PG_4 PG_0_i_3_23 ( .pi(\prop[2][23] ), .gi(\gen[2][23] ), .pj(\prop[2][19] ), 
        .gj(n22), .pout(\prop[3][23] ), .gout(n23) );
  PG_3 PG_0_i_3_31 ( .pi(\prop[2][31] ), .gi(\gen[2][31] ), .pj(\prop[2][27] ), 
        .gj(n1), .pout(\prop[3][31] ), .gout(\gen[3][31] ) );
  G_6 G_jk_4_15_1_0 ( .pi(\prop[3][15] ), .gi(\gen[3][15] ), .gj(n26), .gout(
        n36) );
  G_5 G_jk1_4_15_1_0 ( .pi(\prop[2][11] ), .gi(n30), .gj(n33), .gout(cout[2])
         );
  PG_2 PG_jk_4_31_1_0 ( .pi(\prop[3][31] ), .gi(\gen[3][31] ), .pj(
        \prop[3][23] ), .gj(n29), .pout(\prop[4][31] ), .gout(\gen[4][31] ) );
  PG_1 PG_jk1_4_31_1_0 ( .pi(\prop[2][27] ), .gi(n1), .pj(\prop[3][23] ), .gj(
        n23), .pout(\prop[4][27] ), .gout(\gen[4][27] ) );
  G_4 G_jk_5_31_2_0 ( .pi(\prop[4][31] ), .gi(\gen[4][31] ), .gj(n32), .gout(
        cout[7]) );
  G_3 G_jk_5_31_2_1 ( .pi(\prop[4][27] ), .gi(\gen[4][27] ), .gj(n36), .gout(
        cout[6]) );
  G_2 G_jk_5_31_1_0 ( .pi(\prop[3][23] ), .gi(n29), .gj(n36), .gout(cout[5])
         );
  G_1 G_jk1_5_31_1_0 ( .pi(\prop[2][19] ), .gi(n22), .gj(n36), .gout(cout[4])
         );
  CLKBUF_X1 U1 ( .A(n23), .Z(n29) );
  BUF_X2 U2 ( .A(n36), .Z(cout[3]) );
  CLKBUF_X1 U3 ( .A(n24), .Z(n30) );
  BUF_X1 U4 ( .A(n33), .Z(cout[1]) );
  CLKBUF_X1 U5 ( .A(n26), .Z(n33) );
  CLKBUF_X1 U6 ( .A(cout[3]), .Z(n32) );
  CLKBUF_X1 U7 ( .A(n37), .Z(cout[0]) );
endmodule


module BTB_PC_SIZE32_BTBSIZE5_DW01_cmp6_0 ( A, B, TC, LT, GT, EQ, LE, GE, NE
 );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47;

  NOR4_X1 U1 ( .A1(n1), .A2(n2), .A3(n3), .A4(n4), .ZN(EQ) );
  NAND4_X1 U2 ( .A1(n5), .A2(n6), .A3(n7), .A4(n8), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B[3]), .B(A[3]), .ZN(n8) );
  XNOR2_X1 U4 ( .A(B[4]), .B(A[4]), .ZN(n7) );
  XNOR2_X1 U5 ( .A(B[5]), .B(A[5]), .ZN(n6) );
  XNOR2_X1 U6 ( .A(B[6]), .B(A[6]), .ZN(n5) );
  NAND4_X1 U7 ( .A1(n9), .A2(n10), .A3(n11), .A4(n12), .ZN(n3) );
  OAI22_X1 U8 ( .A1(n13), .A2(n14), .B1(B[1]), .B2(n13), .ZN(n12) );
  INV_X1 U9 ( .A(A[1]), .ZN(n14) );
  AND2_X1 U10 ( .A1(B[0]), .A2(n15), .ZN(n13) );
  OAI22_X1 U11 ( .A1(A[1]), .A2(n16), .B1(n16), .B2(n17), .ZN(n11) );
  INV_X1 U12 ( .A(B[1]), .ZN(n17) );
  NOR2_X1 U13 ( .A1(n15), .A2(B[0]), .ZN(n16) );
  INV_X1 U14 ( .A(A[0]), .ZN(n15) );
  XNOR2_X1 U15 ( .A(B[31]), .B(A[31]), .ZN(n10) );
  XNOR2_X1 U16 ( .A(B[2]), .B(A[2]), .ZN(n9) );
  NAND2_X1 U17 ( .A1(n18), .A2(n19), .ZN(n2) );
  NOR4_X1 U18 ( .A1(n20), .A2(n21), .A3(n22), .A4(n23), .ZN(n19) );
  XOR2_X1 U19 ( .A(B[10]), .B(A[10]), .Z(n23) );
  XOR2_X1 U20 ( .A(B[9]), .B(A[9]), .Z(n22) );
  XOR2_X1 U21 ( .A(B[8]), .B(A[8]), .Z(n21) );
  XOR2_X1 U22 ( .A(B[7]), .B(A[7]), .Z(n20) );
  NOR4_X1 U23 ( .A1(n24), .A2(n25), .A3(n26), .A4(n27), .ZN(n18) );
  XOR2_X1 U24 ( .A(B[14]), .B(A[14]), .Z(n27) );
  XOR2_X1 U25 ( .A(B[13]), .B(A[13]), .Z(n26) );
  XOR2_X1 U26 ( .A(B[12]), .B(A[12]), .Z(n25) );
  XOR2_X1 U27 ( .A(B[11]), .B(A[11]), .Z(n24) );
  NAND4_X1 U28 ( .A1(n28), .A2(n29), .A3(n30), .A4(n31), .ZN(n1) );
  NOR4_X1 U29 ( .A1(n32), .A2(n33), .A3(n34), .A4(n35), .ZN(n31) );
  XOR2_X1 U30 ( .A(B[18]), .B(A[18]), .Z(n35) );
  XOR2_X1 U31 ( .A(B[17]), .B(A[17]), .Z(n34) );
  XOR2_X1 U32 ( .A(B[16]), .B(A[16]), .Z(n33) );
  XOR2_X1 U33 ( .A(B[15]), .B(A[15]), .Z(n32) );
  NOR4_X1 U34 ( .A1(n36), .A2(n37), .A3(n38), .A4(n39), .ZN(n30) );
  XOR2_X1 U35 ( .A(B[22]), .B(A[22]), .Z(n39) );
  XOR2_X1 U36 ( .A(B[21]), .B(A[21]), .Z(n38) );
  XOR2_X1 U37 ( .A(B[20]), .B(A[20]), .Z(n37) );
  XOR2_X1 U38 ( .A(B[19]), .B(A[19]), .Z(n36) );
  NOR4_X1 U39 ( .A1(n40), .A2(n41), .A3(n42), .A4(n43), .ZN(n29) );
  XOR2_X1 U40 ( .A(B[26]), .B(A[26]), .Z(n43) );
  XOR2_X1 U41 ( .A(B[25]), .B(A[25]), .Z(n42) );
  XOR2_X1 U42 ( .A(B[24]), .B(A[24]), .Z(n41) );
  XOR2_X1 U43 ( .A(B[23]), .B(A[23]), .Z(n40) );
  NOR4_X1 U44 ( .A1(n44), .A2(n45), .A3(n46), .A4(n47), .ZN(n28) );
  XOR2_X1 U45 ( .A(B[30]), .B(A[30]), .Z(n47) );
  XOR2_X1 U46 ( .A(B[29]), .B(A[29]), .Z(n46) );
  XOR2_X1 U47 ( .A(B[28]), .B(A[28]), .Z(n45) );
  XOR2_X1 U48 ( .A(B[27]), .B(A[27]), .Z(n44) );
endmodule


module ForwardingUnit_NUMBIT32_ADDRESS_WIDTH_RF5 ( CLK, RST, RS1, RS2, RD_XM, 
        RD_MW, REGWRITE_XM, REGWRITE_MW, ForwardA, forwardB, ForwardC, 
        ForwardD );
  input [4:0] RS1;
  input [4:0] RS2;
  input [4:0] RD_XM;
  input [4:0] RD_MW;
  output [1:0] ForwardA;
  output [1:0] forwardB;
  output [1:0] ForwardD;
  input CLK, RST, REGWRITE_XM, REGWRITE_MW;
  output ForwardC;
  wire   N13, N14, N15, N16, N17, N18, N19, N20, n19, n20, n21, n61, n62, n63,
         n64, n65, net78471, net78472, net78473, net78475, net78476, net78477,
         net78478, net78479, net78481, net78482, net78630, net78629, net78628,
         net78621, net78620, net78618, net78611, net78608, net78606, net78605,
         net78601, net78593, net78592, net78566, net78565, net78564, net78563,
         net78562, net78559, net78558, net95388, net95387, net95500, net95502,
         net95508, net95512, net95523, net95526, net95528, net95530, net95540,
         net95557, net95493, net98500, net98509, net95345, net95344, net78582,
         net78580, net78572, net78571, net78569, net78570, net78568, net78576,
         net78575, net78574, net78573, net78567, net78579, net78577, n1, n6,
         n7, n8, n9, n10, n11, n12, n14, n15, n16, n17, n18, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54;

  DFF_X1 \RS1_DX_reg[4]  ( .D(N17), .CK(CLK), .QN(n19) );
  DFF_X1 \RS1_DX_reg[3]  ( .D(N16), .CK(CLK), .QN(n20) );
  DFF_X1 \RS1_DX_reg[2]  ( .D(N15), .CK(CLK), .QN(n21) );
  DFF_X1 \RS1_DX_reg[1]  ( .D(N14), .CK(CLK), .QN(net78482) );
  DFF_X1 \RS1_DX_reg[0]  ( .D(N13), .CK(CLK), .QN(net78481) );
  DFF_X1 \RS2_DX_reg[2]  ( .D(N20), .CK(CLK), .QN(net78478) );
  DFF_X1 \RS2_DX_reg[1]  ( .D(N19), .CK(CLK), .QN(net78477) );
  DFF_X1 \RS2_DX_reg[0]  ( .D(N18), .CK(CLK), .QN(net78476) );
  DFF_X1 \RS2_DX_reg[4]  ( .D(n9), .CK(CLK), .Q(net78559), .QN(net95493) );
  DFF_X1 \RS2_XM_reg[4]  ( .D(n65), .CK(CLK), .Q(net78558), .QN(net78475) );
  DFF_X1 \RS2_XM_reg[3]  ( .D(n64), .CK(CLK), .Q(n14), .QN(n51) );
  DFF_X1 \RS2_XM_reg[2]  ( .D(n63), .CK(CLK), .QN(net78473) );
  DFF_X1 \RS2_XM_reg[1]  ( .D(n62), .CK(CLK), .QN(net78472) );
  DFF_X1 \RS2_XM_reg[0]  ( .D(n61), .CK(CLK), .QN(net78471) );
  OR4_X1 U3 ( .A1(n35), .A2(net78592), .A3(net78608), .A4(n36), .ZN(n1) );
  INV_X2 U4 ( .A(n1), .ZN(ForwardC) );
  NAND4_X2 U5 ( .A1(n37), .A2(net78611), .A3(n38), .A4(n39), .ZN(n35) );
  NOR2_X1 U6 ( .A1(n6), .A2(net78579), .ZN(net78577) );
  NAND4_X1 U7 ( .A1(net78577), .A2(net78575), .A3(net78576), .A4(net78574), 
        .ZN(net78567) );
  XNOR2_X1 U8 ( .A(RD_XM[4]), .B(net95493), .ZN(net78579) );
  XOR2_X1 U9 ( .A(RD_XM[3]), .B(net95526), .Z(n6) );
  BUF_X1 U10 ( .A(RD_XM[4]), .Z(net95557) );
  XNOR2_X1 U11 ( .A(RD_XM[4]), .B(n19), .ZN(net78628) );
  XOR2_X1 U12 ( .A(net95493), .B(RD_MW[4]), .Z(net78580) );
  BUF_X1 U13 ( .A(RD_XM[3]), .Z(net95502) );
  NOR2_X1 U14 ( .A1(net78559), .A2(net95526), .ZN(net78573) );
  OAI21_X1 U15 ( .B1(net78567), .B2(net78565), .A(net78568), .ZN(net78570) );
  NOR2_X1 U16 ( .A1(net95388), .A2(net78567), .ZN(forwardB[1]) );
  XOR2_X1 U17 ( .A(net78476), .B(RD_XM[0]), .Z(net78574) );
  XOR2_X1 U18 ( .A(net78477), .B(RD_XM[1]), .Z(net78576) );
  XOR2_X1 U19 ( .A(net78478), .B(RD_XM[2]), .Z(net78575) );
  MUX2_X1 U20 ( .A(net78471), .B(net78476), .S(n53), .Z(net78564) );
  XNOR2_X1 U21 ( .A(RD_MW[0]), .B(net78476), .ZN(net78571) );
  NAND4_X1 U22 ( .A1(net78476), .A2(net78478), .A3(net78477), .A4(net78573), 
        .ZN(net78568) );
  CLKBUF_X1 U23 ( .A(RD_XM[0]), .Z(net95512) );
  MUX2_X1 U24 ( .A(net78472), .B(net78477), .S(n53), .Z(net78563) );
  XNOR2_X1 U25 ( .A(RD_MW[1]), .B(net78477), .ZN(net78572) );
  BUF_X1 U26 ( .A(RD_XM[1]), .Z(net95528) );
  MUX2_X1 U27 ( .A(net78473), .B(net78478), .S(n53), .Z(net78562) );
  XOR2_X1 U28 ( .A(net78478), .B(RD_MW[2]), .Z(net78582) );
  BUF_X1 U29 ( .A(RD_XM[2]), .Z(net95540) );
  NOR3_X2 U30 ( .A1(net78570), .A2(net78569), .A3(net95345), .ZN(forwardB[0])
         );
  INV_X2 U31 ( .A(REGWRITE_XM), .ZN(net78565) );
  INV_X1 U32 ( .A(net78568), .ZN(net78566) );
  MUX2_X1 U33 ( .A(net78558), .B(net78559), .S(n53), .Z(n65) );
  INV_X1 U34 ( .A(net95344), .ZN(net95345) );
  NOR2_X1 U35 ( .A1(net78572), .A2(net78571), .ZN(net95344) );
  NAND4_X1 U36 ( .A1(REGWRITE_MW), .A2(net78580), .A3(n7), .A4(net78582), .ZN(
        net78569) );
  XOR2_X1 U37 ( .A(net78479), .B(RD_MW[3]), .Z(n7) );
  CLKBUF_X1 U38 ( .A(RD_MW[0]), .Z(net98500) );
  XOR2_X1 U39 ( .A(RS1[0]), .B(RD_MW[0]), .Z(net78593) );
  BUF_X2 U40 ( .A(RD_MW[1]), .Z(net98509) );
  NAND4_X1 U41 ( .A1(REGWRITE_MW), .A2(net78629), .A3(net78630), .A4(n8), .ZN(
        net78618) );
  INV_X1 U42 ( .A(REGWRITE_MW), .ZN(net78592) );
  XOR2_X1 U43 ( .A(n21), .B(RD_MW[2]), .Z(n8) );
  INV_X1 U44 ( .A(RD_MW[2]), .ZN(net78606) );
  BUF_X1 U46 ( .A(RD_MW[3]), .Z(net95530) );
  BUF_X2 U47 ( .A(RD_MW[4]), .Z(net95508) );
  AND2_X1 U48 ( .A1(RS2[4]), .A2(n53), .ZN(n9) );
  XOR2_X1 U49 ( .A(net78471), .B(net98500), .Z(net78611) );
  XNOR2_X1 U50 ( .A(net78481), .B(net98500), .ZN(net78620) );
  XNOR2_X1 U51 ( .A(net98509), .B(RS1[1]), .ZN(net78605) );
  XNOR2_X1 U52 ( .A(net78472), .B(net98509), .ZN(net78608) );
  XNOR2_X1 U53 ( .A(net78482), .B(net98509), .ZN(net78621) );
  CLKBUF_X1 U54 ( .A(net95526), .Z(net95523) );
  CLKBUF_X1 U55 ( .A(net95530), .Z(net95500) );
  NAND2_X1 U56 ( .A1(n11), .A2(n12), .ZN(n10) );
  AND4_X1 U57 ( .A1(n32), .A2(n33), .A3(n34), .A4(net78605), .ZN(n11) );
  NOR2_X1 U58 ( .A1(net78566), .A2(net78565), .ZN(net95387) );
  INV_X1 U59 ( .A(net95387), .ZN(net95388) );
  NOR3_X1 U60 ( .A1(n18), .A2(n22), .A3(net78565), .ZN(ForwardD[1]) );
  NOR2_X2 U61 ( .A1(n24), .A2(n10), .ZN(ForwardD[0]) );
  NOR4_X4 U62 ( .A1(net78618), .A2(n44), .A3(net78620), .A4(net78621), .ZN(
        ForwardA[0]) );
  NOR2_X1 U63 ( .A1(net78593), .A2(net78592), .ZN(n12) );
  MUX2_X1 U67 ( .A(n14), .B(net95523), .S(n53), .Z(n64) );
  INV_X1 U68 ( .A(net78562), .ZN(n63) );
  INV_X1 U69 ( .A(net78563), .ZN(n62) );
  INV_X1 U70 ( .A(net78564), .ZN(n61) );
  AND2_X1 U71 ( .A1(RS2[2]), .A2(n53), .ZN(N20) );
  AND2_X1 U72 ( .A1(RS2[1]), .A2(n53), .ZN(N19) );
  AND2_X1 U73 ( .A1(RS2[0]), .A2(n53), .ZN(N18) );
  NOR2_X1 U74 ( .A1(n54), .A2(n15), .ZN(N17) );
  NOR2_X1 U75 ( .A1(n54), .A2(n16), .ZN(N16) );
  NOR2_X1 U76 ( .A1(n54), .A2(n17), .ZN(N15) );
  AND2_X1 U77 ( .A1(n53), .A2(RS1[1]), .ZN(N14) );
  AND2_X1 U78 ( .A1(n53), .A2(RS1[0]), .ZN(N13) );
  INV_X1 U79 ( .A(n23), .ZN(n22) );
  OAI21_X1 U80 ( .B1(net78565), .B2(n18), .A(n23), .ZN(n24) );
  NAND4_X1 U81 ( .A1(n16), .A2(n15), .A3(n17), .A4(n25), .ZN(n23) );
  NOR2_X1 U82 ( .A1(RS1[1]), .A2(RS1[0]), .ZN(n25) );
  INV_X1 U83 ( .A(RS1[2]), .ZN(n17) );
  NAND4_X1 U84 ( .A1(n29), .A2(n27), .A3(n28), .A4(n26), .ZN(n18) );
  NOR2_X1 U85 ( .A1(n30), .A2(n31), .ZN(n29) );
  XOR2_X1 U86 ( .A(RS1[4]), .B(net95557), .Z(n31) );
  XOR2_X1 U87 ( .A(RS1[3]), .B(net95502), .Z(n30) );
  XNOR2_X1 U88 ( .A(net95528), .B(RS1[1]), .ZN(n28) );
  XOR2_X1 U89 ( .A(net78601), .B(RS1[2]), .Z(n27) );
  INV_X1 U90 ( .A(net95540), .ZN(net78601) );
  XNOR2_X1 U91 ( .A(net95512), .B(RS1[0]), .ZN(n26) );
  XOR2_X1 U92 ( .A(net78606), .B(RS1[2]), .Z(n34) );
  XOR2_X1 U93 ( .A(net95530), .B(n16), .Z(n33) );
  INV_X1 U94 ( .A(RS1[3]), .ZN(n16) );
  XOR2_X1 U95 ( .A(net95508), .B(n15), .Z(n32) );
  INV_X1 U96 ( .A(RS1[4]), .ZN(n15) );
  XOR2_X1 U97 ( .A(net78473), .B(net78606), .Z(n36) );
  NAND4_X1 U98 ( .A1(net78472), .A2(net78471), .A3(net78473), .A4(n40), .ZN(
        n39) );
  NOR2_X1 U99 ( .A1(n14), .A2(net78558), .ZN(n40) );
  XOR2_X1 U100 ( .A(n51), .B(net95500), .Z(n38) );
  XOR2_X1 U101 ( .A(net78475), .B(net95508), .Z(n37) );
  NOR3_X1 U102 ( .A1(n41), .A2(n42), .A3(net78565), .ZN(ForwardA[1]) );
  INV_X1 U103 ( .A(n43), .ZN(n42) );
  OAI21_X1 U104 ( .B1(net78565), .B2(n41), .A(n43), .ZN(n44) );
  NAND4_X1 U105 ( .A1(net78481), .A2(n21), .A3(net78482), .A4(n45), .ZN(n43)
         );
  AND2_X1 U106 ( .A1(n20), .A2(n19), .ZN(n45) );
  NAND4_X1 U107 ( .A1(n46), .A2(n47), .A3(n48), .A4(n49), .ZN(n41) );
  NOR2_X1 U108 ( .A1(n50), .A2(net78628), .ZN(n49) );
  XNOR2_X1 U109 ( .A(net95502), .B(n20), .ZN(n50) );
  XOR2_X1 U110 ( .A(net78482), .B(net95528), .Z(n48) );
  XOR2_X1 U111 ( .A(n21), .B(net95540), .Z(n47) );
  XOR2_X1 U112 ( .A(net78481), .B(net95512), .Z(n46) );
  XOR2_X1 U113 ( .A(n20), .B(net95530), .Z(net78630) );
  XOR2_X1 U114 ( .A(n19), .B(net95508), .Z(net78629) );
  DFF_X1 \RS2_DX_reg[3]  ( .D(n52), .CK(CLK), .Q(net95526), .QN(net78479) );
  AND2_X1 U45 ( .A1(RS2[3]), .A2(n53), .ZN(n52) );
  INV_X1 U64 ( .A(n54), .ZN(n53) );
  INV_X2 U65 ( .A(RST), .ZN(n54) );
endmodule


module MUX21_GENERIC_N5 ( A, B, SEL, Y );
  input [4:0] A;
  input [4:0] B;
  output [4:0] Y;
  input SEL;
  wire   n2, n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(n2), .ZN(Y[4]) );
  AOI22_X1 U2 ( .A1(SEL), .A2(A[4]), .B1(B[4]), .B2(n3), .ZN(n2) );
  INV_X1 U3 ( .A(n4), .ZN(Y[3]) );
  AOI22_X1 U4 ( .A1(A[3]), .A2(SEL), .B1(B[3]), .B2(n3), .ZN(n4) );
  INV_X1 U5 ( .A(n5), .ZN(Y[2]) );
  AOI22_X1 U6 ( .A1(A[2]), .A2(SEL), .B1(B[2]), .B2(n3), .ZN(n5) );
  INV_X1 U7 ( .A(n6), .ZN(Y[1]) );
  AOI22_X1 U8 ( .A1(A[1]), .A2(SEL), .B1(B[1]), .B2(n3), .ZN(n6) );
  INV_X1 U9 ( .A(n7), .ZN(Y[0]) );
  AOI22_X1 U10 ( .A1(A[0]), .A2(SEL), .B1(B[0]), .B2(n3), .ZN(n7) );
  INV_X1 U11 ( .A(SEL), .ZN(n3) );
endmodule


module MUX21 ( A, B, SEL, Y );
  input A, B, SEL;
  output Y;
  wire   n4, n2, n3;

  INV_X1 U3 ( .A(SEL), .ZN(n3) );
  BUF_X2 U1 ( .A(n4), .Z(Y) );
  INV_X1 U2 ( .A(n2), .ZN(n4) );
  AOI22_X1 U4 ( .A1(SEL), .A2(A), .B1(B), .B2(n3), .ZN(n2) );
endmodule


module BranchMgmt_NUMBIT32 ( Rin, Cond, Jump, Branch );
  input [31:0] Rin;
  input Cond, Jump;
  output Branch;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13;

  OR2_X1 U2 ( .A1(n2), .A2(Jump), .ZN(Branch) );
  XNOR2_X1 U3 ( .A(n3), .B(Cond), .ZN(n2) );
  NOR2_X1 U4 ( .A1(n4), .A2(n5), .ZN(n3) );
  NAND4_X1 U5 ( .A1(n6), .A2(n7), .A3(n8), .A4(n9), .ZN(n5) );
  NOR4_X1 U6 ( .A1(Rin[23]), .A2(Rin[22]), .A3(Rin[21]), .A4(Rin[20]), .ZN(n9)
         );
  NOR4_X1 U7 ( .A1(Rin[1]), .A2(Rin[19]), .A3(Rin[18]), .A4(Rin[17]), .ZN(n8)
         );
  NOR4_X1 U8 ( .A1(Rin[16]), .A2(Rin[15]), .A3(Rin[14]), .A4(Rin[13]), .ZN(n7)
         );
  NOR4_X1 U9 ( .A1(Rin[12]), .A2(Rin[11]), .A3(Rin[10]), .A4(Rin[0]), .ZN(n6)
         );
  NAND4_X1 U10 ( .A1(n12), .A2(n11), .A3(n10), .A4(n13), .ZN(n4) );
  NOR4_X1 U11 ( .A1(Rin[9]), .A2(Rin[8]), .A3(Rin[7]), .A4(Rin[6]), .ZN(n13)
         );
  NOR4_X1 U12 ( .A1(Rin[5]), .A2(Rin[4]), .A3(Rin[3]), .A4(Rin[31]), .ZN(n12)
         );
  NOR4_X1 U13 ( .A1(Rin[30]), .A2(Rin[2]), .A3(Rin[29]), .A4(Rin[28]), .ZN(n11) );
  NOR4_X1 U14 ( .A1(Rin[27]), .A2(Rin[26]), .A3(Rin[25]), .A4(Rin[24]), .ZN(
        n10) );
endmodule


module signExtend_NUMBIT_in26_NUMBIT_out32 ( in_s, sign_unsign, out_s );
  input [25:0] in_s;
  output [31:0] out_s;
  input sign_unsign;
  wire   out_s_31;
  assign out_s[31] = out_s_31;
  assign out_s[30] = out_s_31;
  assign out_s[29] = out_s_31;
  assign out_s[28] = out_s_31;
  assign out_s[27] = out_s_31;
  assign out_s[26] = out_s_31;
  assign out_s[25] = in_s[25];
  assign out_s[24] = in_s[24];
  assign out_s[23] = in_s[23];
  assign out_s[22] = in_s[22];
  assign out_s[21] = in_s[21];
  assign out_s[20] = in_s[20];
  assign out_s[19] = in_s[19];
  assign out_s[18] = in_s[18];
  assign out_s[17] = in_s[17];
  assign out_s[16] = in_s[16];
  assign out_s[15] = in_s[15];
  assign out_s[14] = in_s[14];
  assign out_s[13] = in_s[13];
  assign out_s[12] = in_s[12];
  assign out_s[11] = in_s[11];
  assign out_s[10] = in_s[10];
  assign out_s[9] = in_s[9];
  assign out_s[8] = in_s[8];
  assign out_s[7] = in_s[7];
  assign out_s[6] = in_s[6];
  assign out_s[5] = in_s[5];
  assign out_s[4] = in_s[4];
  assign out_s[3] = in_s[3];
  assign out_s[2] = in_s[2];
  assign out_s[1] = in_s[1];
  assign out_s[0] = in_s[0];

  AND2_X1 U1 ( .A1(sign_unsign), .A2(in_s[25]), .ZN(out_s_31) );
endmodule


module signExtend_NUMBIT_in16_NUMBIT_out32 ( in_s, sign_unsign, out_s );
  input [15:0] in_s;
  output [31:0] out_s;
  input sign_unsign;
  wire   out_s_31;
  assign out_s[31] = out_s_31;
  assign out_s[30] = out_s_31;
  assign out_s[29] = out_s_31;
  assign out_s[28] = out_s_31;
  assign out_s[27] = out_s_31;
  assign out_s[26] = out_s_31;
  assign out_s[25] = out_s_31;
  assign out_s[24] = out_s_31;
  assign out_s[23] = out_s_31;
  assign out_s[22] = out_s_31;
  assign out_s[21] = out_s_31;
  assign out_s[20] = out_s_31;
  assign out_s[19] = out_s_31;
  assign out_s[18] = out_s_31;
  assign out_s[17] = out_s_31;
  assign out_s[16] = out_s_31;
  assign out_s[15] = in_s[15];
  assign out_s[14] = in_s[14];
  assign out_s[13] = in_s[13];
  assign out_s[12] = in_s[12];
  assign out_s[11] = in_s[11];
  assign out_s[10] = in_s[10];
  assign out_s[9] = in_s[9];
  assign out_s[8] = in_s[8];
  assign out_s[7] = in_s[7];
  assign out_s[6] = in_s[6];
  assign out_s[5] = in_s[5];
  assign out_s[4] = in_s[4];
  assign out_s[3] = in_s[3];
  assign out_s[2] = in_s[2];
  assign out_s[1] = in_s[1];
  assign out_s[0] = in_s[0];

  AND2_X1 U1 ( .A1(sign_unsign), .A2(in_s[15]), .ZN(out_s_31) );
endmodule


module register_file_NUMBIT32_BITADDR5 ( CLK, RESET, ENABLE, RD1, RD2, WR, 
        ADD_WR, ADD_RD1, ADD_RD2, DATAIN, OUT1, OUT2 );
  input [4:0] ADD_WR;
  input [4:0] ADD_RD1;
  input [4:0] ADD_RD2;
  input [31:0] DATAIN;
  output [31:0] OUT1;
  output [31:0] OUT2;
  input CLK, RESET, ENABLE, RD1, RD2, WR;
  wire   \REGISTERS[1][31] , \REGISTERS[1][30] , \REGISTERS[1][29] ,
         \REGISTERS[1][28] , \REGISTERS[1][27] , \REGISTERS[1][26] ,
         \REGISTERS[1][25] , \REGISTERS[1][24] , \REGISTERS[1][23] ,
         \REGISTERS[1][22] , \REGISTERS[1][21] , \REGISTERS[1][20] ,
         \REGISTERS[1][19] , \REGISTERS[1][18] , \REGISTERS[1][17] ,
         \REGISTERS[1][16] , \REGISTERS[1][15] , \REGISTERS[1][14] ,
         \REGISTERS[1][13] , \REGISTERS[1][12] , \REGISTERS[1][11] ,
         \REGISTERS[1][10] , \REGISTERS[1][9] , \REGISTERS[1][8] ,
         \REGISTERS[1][7] , \REGISTERS[1][6] , \REGISTERS[1][5] ,
         \REGISTERS[1][4] , \REGISTERS[1][3] , \REGISTERS[1][2] ,
         \REGISTERS[1][1] , \REGISTERS[1][0] , \REGISTERS[2][31] ,
         \REGISTERS[2][30] , \REGISTERS[2][29] , \REGISTERS[2][28] ,
         \REGISTERS[2][27] , \REGISTERS[2][26] , \REGISTERS[2][25] ,
         \REGISTERS[2][24] , \REGISTERS[2][23] , \REGISTERS[2][22] ,
         \REGISTERS[2][21] , \REGISTERS[2][20] , \REGISTERS[2][19] ,
         \REGISTERS[2][18] , \REGISTERS[2][17] , \REGISTERS[2][16] ,
         \REGISTERS[2][15] , \REGISTERS[2][14] , \REGISTERS[2][13] ,
         \REGISTERS[2][12] , \REGISTERS[2][11] , \REGISTERS[2][10] ,
         \REGISTERS[2][9] , \REGISTERS[2][8] , \REGISTERS[2][7] ,
         \REGISTERS[2][6] , \REGISTERS[2][5] , \REGISTERS[2][4] ,
         \REGISTERS[2][3] , \REGISTERS[2][2] , \REGISTERS[2][1] ,
         \REGISTERS[2][0] , \REGISTERS[3][31] , \REGISTERS[3][30] ,
         \REGISTERS[3][29] , \REGISTERS[3][28] , \REGISTERS[3][27] ,
         \REGISTERS[3][26] , \REGISTERS[3][25] , \REGISTERS[3][24] ,
         \REGISTERS[3][23] , \REGISTERS[3][22] , \REGISTERS[3][21] ,
         \REGISTERS[3][20] , \REGISTERS[3][19] , \REGISTERS[3][18] ,
         \REGISTERS[3][17] , \REGISTERS[3][16] , \REGISTERS[3][15] ,
         \REGISTERS[3][14] , \REGISTERS[3][13] , \REGISTERS[3][12] ,
         \REGISTERS[3][11] , \REGISTERS[3][10] , \REGISTERS[3][9] ,
         \REGISTERS[3][8] , \REGISTERS[3][7] , \REGISTERS[3][6] ,
         \REGISTERS[3][5] , \REGISTERS[3][4] , \REGISTERS[3][3] ,
         \REGISTERS[3][2] , \REGISTERS[3][1] , \REGISTERS[3][0] ,
         \REGISTERS[4][31] , \REGISTERS[4][30] , \REGISTERS[4][29] ,
         \REGISTERS[4][28] , \REGISTERS[4][27] , \REGISTERS[4][26] ,
         \REGISTERS[4][25] , \REGISTERS[4][24] , \REGISTERS[4][23] ,
         \REGISTERS[4][22] , \REGISTERS[4][21] , \REGISTERS[4][20] ,
         \REGISTERS[4][19] , \REGISTERS[4][18] , \REGISTERS[4][17] ,
         \REGISTERS[4][16] , \REGISTERS[4][15] , \REGISTERS[4][14] ,
         \REGISTERS[4][13] , \REGISTERS[4][12] , \REGISTERS[4][11] ,
         \REGISTERS[4][10] , \REGISTERS[4][9] , \REGISTERS[4][8] ,
         \REGISTERS[4][7] , \REGISTERS[4][6] , \REGISTERS[4][5] ,
         \REGISTERS[4][4] , \REGISTERS[4][3] , \REGISTERS[4][2] ,
         \REGISTERS[4][1] , \REGISTERS[4][0] , \REGISTERS[5][31] ,
         \REGISTERS[5][30] , \REGISTERS[5][29] , \REGISTERS[5][28] ,
         \REGISTERS[5][27] , \REGISTERS[5][26] , \REGISTERS[5][25] ,
         \REGISTERS[5][24] , \REGISTERS[5][23] , \REGISTERS[5][22] ,
         \REGISTERS[5][21] , \REGISTERS[5][20] , \REGISTERS[5][19] ,
         \REGISTERS[5][18] , \REGISTERS[5][17] , \REGISTERS[5][16] ,
         \REGISTERS[5][15] , \REGISTERS[5][14] , \REGISTERS[5][13] ,
         \REGISTERS[5][12] , \REGISTERS[5][11] , \REGISTERS[5][10] ,
         \REGISTERS[5][9] , \REGISTERS[5][8] , \REGISTERS[5][7] ,
         \REGISTERS[5][6] , \REGISTERS[5][5] , \REGISTERS[5][4] ,
         \REGISTERS[5][3] , \REGISTERS[5][2] , \REGISTERS[5][1] ,
         \REGISTERS[5][0] , \REGISTERS[6][31] , \REGISTERS[6][30] ,
         \REGISTERS[6][29] , \REGISTERS[6][28] , \REGISTERS[6][27] ,
         \REGISTERS[6][26] , \REGISTERS[6][25] , \REGISTERS[6][24] ,
         \REGISTERS[6][23] , \REGISTERS[6][22] , \REGISTERS[6][21] ,
         \REGISTERS[6][20] , \REGISTERS[6][19] , \REGISTERS[6][18] ,
         \REGISTERS[6][17] , \REGISTERS[6][16] , \REGISTERS[6][15] ,
         \REGISTERS[6][14] , \REGISTERS[6][13] , \REGISTERS[6][12] ,
         \REGISTERS[6][11] , \REGISTERS[6][10] , \REGISTERS[6][9] ,
         \REGISTERS[6][8] , \REGISTERS[6][7] , \REGISTERS[6][6] ,
         \REGISTERS[6][5] , \REGISTERS[6][4] , \REGISTERS[6][3] ,
         \REGISTERS[6][2] , \REGISTERS[6][1] , \REGISTERS[6][0] ,
         \REGISTERS[7][31] , \REGISTERS[7][30] , \REGISTERS[7][29] ,
         \REGISTERS[7][28] , \REGISTERS[7][27] , \REGISTERS[7][26] ,
         \REGISTERS[7][25] , \REGISTERS[7][24] , \REGISTERS[7][23] ,
         \REGISTERS[7][22] , \REGISTERS[7][21] , \REGISTERS[7][20] ,
         \REGISTERS[7][19] , \REGISTERS[7][18] , \REGISTERS[7][17] ,
         \REGISTERS[7][16] , \REGISTERS[7][15] , \REGISTERS[7][14] ,
         \REGISTERS[7][13] , \REGISTERS[7][12] , \REGISTERS[7][11] ,
         \REGISTERS[7][10] , \REGISTERS[7][9] , \REGISTERS[7][8] ,
         \REGISTERS[7][7] , \REGISTERS[7][6] , \REGISTERS[7][5] ,
         \REGISTERS[7][4] , \REGISTERS[7][3] , \REGISTERS[7][2] ,
         \REGISTERS[7][1] , \REGISTERS[7][0] , \REGISTERS[8][31] ,
         \REGISTERS[8][30] , \REGISTERS[8][29] , \REGISTERS[8][28] ,
         \REGISTERS[8][27] , \REGISTERS[8][26] , \REGISTERS[8][25] ,
         \REGISTERS[8][24] , \REGISTERS[8][23] , \REGISTERS[8][22] ,
         \REGISTERS[8][21] , \REGISTERS[8][20] , \REGISTERS[8][19] ,
         \REGISTERS[8][18] , \REGISTERS[8][17] , \REGISTERS[8][16] ,
         \REGISTERS[8][15] , \REGISTERS[8][14] , \REGISTERS[8][13] ,
         \REGISTERS[8][12] , \REGISTERS[8][11] , \REGISTERS[8][10] ,
         \REGISTERS[8][9] , \REGISTERS[8][8] , \REGISTERS[8][7] ,
         \REGISTERS[8][6] , \REGISTERS[8][5] , \REGISTERS[8][4] ,
         \REGISTERS[8][3] , \REGISTERS[8][2] , \REGISTERS[8][1] ,
         \REGISTERS[8][0] , \REGISTERS[9][31] , \REGISTERS[9][30] ,
         \REGISTERS[9][29] , \REGISTERS[9][28] , \REGISTERS[9][27] ,
         \REGISTERS[9][26] , \REGISTERS[9][25] , \REGISTERS[9][24] ,
         \REGISTERS[9][23] , \REGISTERS[9][22] , \REGISTERS[9][21] ,
         \REGISTERS[9][20] , \REGISTERS[9][19] , \REGISTERS[9][18] ,
         \REGISTERS[9][17] , \REGISTERS[9][16] , \REGISTERS[9][15] ,
         \REGISTERS[9][14] , \REGISTERS[9][13] , \REGISTERS[9][12] ,
         \REGISTERS[9][11] , \REGISTERS[9][10] , \REGISTERS[9][9] ,
         \REGISTERS[9][8] , \REGISTERS[9][7] , \REGISTERS[9][6] ,
         \REGISTERS[9][5] , \REGISTERS[9][4] , \REGISTERS[9][3] ,
         \REGISTERS[9][2] , \REGISTERS[9][1] , \REGISTERS[9][0] ,
         \REGISTERS[10][31] , \REGISTERS[10][30] , \REGISTERS[10][29] ,
         \REGISTERS[10][28] , \REGISTERS[10][27] , \REGISTERS[10][26] ,
         \REGISTERS[10][25] , \REGISTERS[10][24] , \REGISTERS[10][23] ,
         \REGISTERS[10][22] , \REGISTERS[10][21] , \REGISTERS[10][20] ,
         \REGISTERS[10][19] , \REGISTERS[10][18] , \REGISTERS[10][17] ,
         \REGISTERS[10][16] , \REGISTERS[10][15] , \REGISTERS[10][14] ,
         \REGISTERS[10][13] , \REGISTERS[10][12] , \REGISTERS[10][11] ,
         \REGISTERS[10][10] , \REGISTERS[10][9] , \REGISTERS[10][8] ,
         \REGISTERS[10][7] , \REGISTERS[10][6] , \REGISTERS[10][5] ,
         \REGISTERS[10][4] , \REGISTERS[10][3] , \REGISTERS[10][2] ,
         \REGISTERS[10][1] , \REGISTERS[10][0] , \REGISTERS[11][31] ,
         \REGISTERS[11][30] , \REGISTERS[11][29] , \REGISTERS[11][28] ,
         \REGISTERS[11][27] , \REGISTERS[11][26] , \REGISTERS[11][25] ,
         \REGISTERS[11][24] , \REGISTERS[11][23] , \REGISTERS[11][22] ,
         \REGISTERS[11][21] , \REGISTERS[11][20] , \REGISTERS[11][19] ,
         \REGISTERS[11][18] , \REGISTERS[11][17] , \REGISTERS[11][16] ,
         \REGISTERS[11][15] , \REGISTERS[11][14] , \REGISTERS[11][13] ,
         \REGISTERS[11][12] , \REGISTERS[11][11] , \REGISTERS[11][10] ,
         \REGISTERS[11][9] , \REGISTERS[11][8] , \REGISTERS[11][7] ,
         \REGISTERS[11][6] , \REGISTERS[11][5] , \REGISTERS[11][4] ,
         \REGISTERS[11][3] , \REGISTERS[11][2] , \REGISTERS[11][1] ,
         \REGISTERS[11][0] , \REGISTERS[12][31] , \REGISTERS[12][30] ,
         \REGISTERS[12][29] , \REGISTERS[12][28] , \REGISTERS[12][27] ,
         \REGISTERS[12][26] , \REGISTERS[12][25] , \REGISTERS[12][24] ,
         \REGISTERS[12][23] , \REGISTERS[12][22] , \REGISTERS[12][21] ,
         \REGISTERS[12][20] , \REGISTERS[12][19] , \REGISTERS[12][18] ,
         \REGISTERS[12][17] , \REGISTERS[12][16] , \REGISTERS[12][15] ,
         \REGISTERS[12][14] , \REGISTERS[12][13] , \REGISTERS[12][12] ,
         \REGISTERS[12][11] , \REGISTERS[12][10] , \REGISTERS[12][9] ,
         \REGISTERS[12][8] , \REGISTERS[12][7] , \REGISTERS[12][6] ,
         \REGISTERS[12][5] , \REGISTERS[12][4] , \REGISTERS[12][3] ,
         \REGISTERS[12][2] , \REGISTERS[12][1] , \REGISTERS[12][0] ,
         \REGISTERS[13][31] , \REGISTERS[13][30] , \REGISTERS[13][29] ,
         \REGISTERS[13][28] , \REGISTERS[13][27] , \REGISTERS[13][26] ,
         \REGISTERS[13][25] , \REGISTERS[13][24] , \REGISTERS[13][23] ,
         \REGISTERS[13][22] , \REGISTERS[13][21] , \REGISTERS[13][20] ,
         \REGISTERS[13][19] , \REGISTERS[13][18] , \REGISTERS[13][17] ,
         \REGISTERS[13][16] , \REGISTERS[13][15] , \REGISTERS[13][14] ,
         \REGISTERS[13][13] , \REGISTERS[13][12] , \REGISTERS[13][11] ,
         \REGISTERS[13][10] , \REGISTERS[13][9] , \REGISTERS[13][8] ,
         \REGISTERS[13][7] , \REGISTERS[13][6] , \REGISTERS[13][5] ,
         \REGISTERS[13][4] , \REGISTERS[13][3] , \REGISTERS[13][2] ,
         \REGISTERS[13][1] , \REGISTERS[13][0] , \REGISTERS[14][31] ,
         \REGISTERS[14][30] , \REGISTERS[14][29] , \REGISTERS[14][28] ,
         \REGISTERS[14][27] , \REGISTERS[14][26] , \REGISTERS[14][25] ,
         \REGISTERS[14][24] , \REGISTERS[14][23] , \REGISTERS[14][22] ,
         \REGISTERS[14][21] , \REGISTERS[14][20] , \REGISTERS[14][19] ,
         \REGISTERS[14][18] , \REGISTERS[14][17] , \REGISTERS[14][16] ,
         \REGISTERS[14][15] , \REGISTERS[14][14] , \REGISTERS[14][13] ,
         \REGISTERS[14][12] , \REGISTERS[14][11] , \REGISTERS[14][10] ,
         \REGISTERS[14][9] , \REGISTERS[14][8] , \REGISTERS[14][7] ,
         \REGISTERS[14][6] , \REGISTERS[14][5] , \REGISTERS[14][4] ,
         \REGISTERS[14][3] , \REGISTERS[14][2] , \REGISTERS[14][1] ,
         \REGISTERS[14][0] , \REGISTERS[15][31] , \REGISTERS[15][30] ,
         \REGISTERS[15][29] , \REGISTERS[15][28] , \REGISTERS[15][27] ,
         \REGISTERS[15][26] , \REGISTERS[15][25] , \REGISTERS[15][24] ,
         \REGISTERS[15][23] , \REGISTERS[15][22] , \REGISTERS[15][21] ,
         \REGISTERS[15][20] , \REGISTERS[15][19] , \REGISTERS[15][18] ,
         \REGISTERS[15][17] , \REGISTERS[15][16] , \REGISTERS[15][15] ,
         \REGISTERS[15][14] , \REGISTERS[15][13] , \REGISTERS[15][12] ,
         \REGISTERS[15][11] , \REGISTERS[15][10] , \REGISTERS[15][9] ,
         \REGISTERS[15][8] , \REGISTERS[15][7] , \REGISTERS[15][6] ,
         \REGISTERS[15][5] , \REGISTERS[15][4] , \REGISTERS[15][3] ,
         \REGISTERS[15][2] , \REGISTERS[15][1] , \REGISTERS[15][0] ,
         \REGISTERS[16][31] , \REGISTERS[16][30] , \REGISTERS[16][29] ,
         \REGISTERS[16][28] , \REGISTERS[16][27] , \REGISTERS[16][26] ,
         \REGISTERS[16][25] , \REGISTERS[16][24] , \REGISTERS[16][23] ,
         \REGISTERS[16][22] , \REGISTERS[16][21] , \REGISTERS[16][20] ,
         \REGISTERS[16][19] , \REGISTERS[16][18] , \REGISTERS[16][17] ,
         \REGISTERS[16][16] , \REGISTERS[16][15] , \REGISTERS[16][14] ,
         \REGISTERS[16][13] , \REGISTERS[16][12] , \REGISTERS[16][11] ,
         \REGISTERS[16][10] , \REGISTERS[16][9] , \REGISTERS[16][8] ,
         \REGISTERS[16][7] , \REGISTERS[16][6] , \REGISTERS[16][5] ,
         \REGISTERS[16][4] , \REGISTERS[16][3] , \REGISTERS[16][2] ,
         \REGISTERS[16][1] , \REGISTERS[16][0] , \REGISTERS[17][31] ,
         \REGISTERS[17][30] , \REGISTERS[17][29] , \REGISTERS[17][28] ,
         \REGISTERS[17][27] , \REGISTERS[17][26] , \REGISTERS[17][25] ,
         \REGISTERS[17][24] , \REGISTERS[17][23] , \REGISTERS[17][22] ,
         \REGISTERS[17][21] , \REGISTERS[17][20] , \REGISTERS[17][19] ,
         \REGISTERS[17][18] , \REGISTERS[17][17] , \REGISTERS[17][16] ,
         \REGISTERS[17][15] , \REGISTERS[17][14] , \REGISTERS[17][13] ,
         \REGISTERS[17][12] , \REGISTERS[17][11] , \REGISTERS[17][10] ,
         \REGISTERS[17][9] , \REGISTERS[17][8] , \REGISTERS[17][7] ,
         \REGISTERS[17][6] , \REGISTERS[17][5] , \REGISTERS[17][4] ,
         \REGISTERS[17][3] , \REGISTERS[17][2] , \REGISTERS[17][1] ,
         \REGISTERS[17][0] , \REGISTERS[18][31] , \REGISTERS[18][30] ,
         \REGISTERS[18][29] , \REGISTERS[18][28] , \REGISTERS[18][27] ,
         \REGISTERS[18][26] , \REGISTERS[18][25] , \REGISTERS[18][24] ,
         \REGISTERS[18][23] , \REGISTERS[18][22] , \REGISTERS[18][21] ,
         \REGISTERS[18][20] , \REGISTERS[18][19] , \REGISTERS[18][18] ,
         \REGISTERS[18][17] , \REGISTERS[18][16] , \REGISTERS[18][15] ,
         \REGISTERS[18][14] , \REGISTERS[18][13] , \REGISTERS[18][12] ,
         \REGISTERS[18][11] , \REGISTERS[18][10] , \REGISTERS[18][9] ,
         \REGISTERS[18][8] , \REGISTERS[18][7] , \REGISTERS[18][6] ,
         \REGISTERS[18][5] , \REGISTERS[18][4] , \REGISTERS[18][3] ,
         \REGISTERS[18][2] , \REGISTERS[18][1] , \REGISTERS[18][0] ,
         \REGISTERS[19][31] , \REGISTERS[19][30] , \REGISTERS[19][29] ,
         \REGISTERS[19][28] , \REGISTERS[19][27] , \REGISTERS[19][26] ,
         \REGISTERS[19][25] , \REGISTERS[19][24] , \REGISTERS[19][23] ,
         \REGISTERS[19][22] , \REGISTERS[19][21] , \REGISTERS[19][20] ,
         \REGISTERS[19][19] , \REGISTERS[19][18] , \REGISTERS[19][17] ,
         \REGISTERS[19][16] , \REGISTERS[19][15] , \REGISTERS[19][14] ,
         \REGISTERS[19][13] , \REGISTERS[19][12] , \REGISTERS[19][11] ,
         \REGISTERS[19][10] , \REGISTERS[19][9] , \REGISTERS[19][8] ,
         \REGISTERS[19][7] , \REGISTERS[19][6] , \REGISTERS[19][5] ,
         \REGISTERS[19][4] , \REGISTERS[19][3] , \REGISTERS[19][2] ,
         \REGISTERS[19][1] , \REGISTERS[19][0] , \REGISTERS[20][31] ,
         \REGISTERS[20][30] , \REGISTERS[20][29] , \REGISTERS[20][28] ,
         \REGISTERS[20][27] , \REGISTERS[20][26] , \REGISTERS[20][25] ,
         \REGISTERS[20][24] , \REGISTERS[20][23] , \REGISTERS[20][22] ,
         \REGISTERS[20][21] , \REGISTERS[20][20] , \REGISTERS[20][19] ,
         \REGISTERS[20][18] , \REGISTERS[20][17] , \REGISTERS[20][16] ,
         \REGISTERS[20][15] , \REGISTERS[20][14] , \REGISTERS[20][13] ,
         \REGISTERS[20][12] , \REGISTERS[20][11] , \REGISTERS[20][10] ,
         \REGISTERS[20][9] , \REGISTERS[20][8] , \REGISTERS[20][7] ,
         \REGISTERS[20][6] , \REGISTERS[20][5] , \REGISTERS[20][4] ,
         \REGISTERS[20][3] , \REGISTERS[20][2] , \REGISTERS[20][1] ,
         \REGISTERS[20][0] , \REGISTERS[21][31] , \REGISTERS[21][30] ,
         \REGISTERS[21][29] , \REGISTERS[21][28] , \REGISTERS[21][27] ,
         \REGISTERS[21][26] , \REGISTERS[21][25] , \REGISTERS[21][24] ,
         \REGISTERS[21][23] , \REGISTERS[21][22] , \REGISTERS[21][21] ,
         \REGISTERS[21][20] , \REGISTERS[21][19] , \REGISTERS[21][18] ,
         \REGISTERS[21][17] , \REGISTERS[21][16] , \REGISTERS[21][15] ,
         \REGISTERS[21][14] , \REGISTERS[21][13] , \REGISTERS[21][12] ,
         \REGISTERS[21][11] , \REGISTERS[21][10] , \REGISTERS[21][9] ,
         \REGISTERS[21][8] , \REGISTERS[21][7] , \REGISTERS[21][6] ,
         \REGISTERS[21][5] , \REGISTERS[21][4] , \REGISTERS[21][3] ,
         \REGISTERS[21][2] , \REGISTERS[21][1] , \REGISTERS[21][0] ,
         \REGISTERS[22][31] , \REGISTERS[22][30] , \REGISTERS[22][29] ,
         \REGISTERS[22][28] , \REGISTERS[22][27] , \REGISTERS[22][26] ,
         \REGISTERS[22][25] , \REGISTERS[22][24] , \REGISTERS[22][23] ,
         \REGISTERS[22][22] , \REGISTERS[22][21] , \REGISTERS[22][20] ,
         \REGISTERS[22][19] , \REGISTERS[22][18] , \REGISTERS[22][17] ,
         \REGISTERS[22][16] , \REGISTERS[22][15] , \REGISTERS[22][14] ,
         \REGISTERS[22][13] , \REGISTERS[22][12] , \REGISTERS[22][11] ,
         \REGISTERS[22][10] , \REGISTERS[22][9] , \REGISTERS[22][8] ,
         \REGISTERS[22][7] , \REGISTERS[22][6] , \REGISTERS[22][5] ,
         \REGISTERS[22][4] , \REGISTERS[22][3] , \REGISTERS[22][2] ,
         \REGISTERS[22][1] , \REGISTERS[22][0] , \REGISTERS[23][31] ,
         \REGISTERS[23][30] , \REGISTERS[23][29] , \REGISTERS[23][28] ,
         \REGISTERS[23][27] , \REGISTERS[23][26] , \REGISTERS[23][25] ,
         \REGISTERS[23][24] , \REGISTERS[23][23] , \REGISTERS[23][22] ,
         \REGISTERS[23][21] , \REGISTERS[23][20] , \REGISTERS[23][19] ,
         \REGISTERS[23][18] , \REGISTERS[23][17] , \REGISTERS[23][16] ,
         \REGISTERS[23][15] , \REGISTERS[23][14] , \REGISTERS[23][13] ,
         \REGISTERS[23][12] , \REGISTERS[23][11] , \REGISTERS[23][10] ,
         \REGISTERS[23][9] , \REGISTERS[23][8] , \REGISTERS[23][7] ,
         \REGISTERS[23][6] , \REGISTERS[23][5] , \REGISTERS[23][4] ,
         \REGISTERS[23][3] , \REGISTERS[23][2] , \REGISTERS[23][1] ,
         \REGISTERS[23][0] , \REGISTERS[24][31] , \REGISTERS[24][30] ,
         \REGISTERS[24][29] , \REGISTERS[24][28] , \REGISTERS[24][27] ,
         \REGISTERS[24][26] , \REGISTERS[24][25] , \REGISTERS[24][24] ,
         \REGISTERS[24][23] , \REGISTERS[24][22] , \REGISTERS[24][21] ,
         \REGISTERS[24][20] , \REGISTERS[24][19] , \REGISTERS[24][18] ,
         \REGISTERS[24][17] , \REGISTERS[24][16] , \REGISTERS[24][15] ,
         \REGISTERS[24][14] , \REGISTERS[24][13] , \REGISTERS[24][12] ,
         \REGISTERS[24][11] , \REGISTERS[24][10] , \REGISTERS[24][9] ,
         \REGISTERS[24][8] , \REGISTERS[24][7] , \REGISTERS[24][6] ,
         \REGISTERS[24][5] , \REGISTERS[24][4] , \REGISTERS[24][3] ,
         \REGISTERS[24][2] , \REGISTERS[24][1] , \REGISTERS[24][0] ,
         \REGISTERS[25][31] , \REGISTERS[25][30] , \REGISTERS[25][29] ,
         \REGISTERS[25][28] , \REGISTERS[25][27] , \REGISTERS[25][26] ,
         \REGISTERS[25][25] , \REGISTERS[25][24] , \REGISTERS[25][23] ,
         \REGISTERS[25][22] , \REGISTERS[25][21] , \REGISTERS[25][20] ,
         \REGISTERS[25][19] , \REGISTERS[25][18] , \REGISTERS[25][17] ,
         \REGISTERS[25][16] , \REGISTERS[25][15] , \REGISTERS[25][14] ,
         \REGISTERS[25][13] , \REGISTERS[25][12] , \REGISTERS[25][11] ,
         \REGISTERS[25][10] , \REGISTERS[25][9] , \REGISTERS[25][8] ,
         \REGISTERS[25][7] , \REGISTERS[25][6] , \REGISTERS[25][5] ,
         \REGISTERS[25][4] , \REGISTERS[25][3] , \REGISTERS[25][2] ,
         \REGISTERS[25][1] , \REGISTERS[25][0] , \REGISTERS[26][31] ,
         \REGISTERS[26][30] , \REGISTERS[26][29] , \REGISTERS[26][28] ,
         \REGISTERS[26][27] , \REGISTERS[26][26] , \REGISTERS[26][25] ,
         \REGISTERS[26][24] , \REGISTERS[26][23] , \REGISTERS[26][22] ,
         \REGISTERS[26][21] , \REGISTERS[26][20] , \REGISTERS[26][19] ,
         \REGISTERS[26][18] , \REGISTERS[26][17] , \REGISTERS[26][16] ,
         \REGISTERS[26][15] , \REGISTERS[26][14] , \REGISTERS[26][13] ,
         \REGISTERS[26][12] , \REGISTERS[26][11] , \REGISTERS[26][10] ,
         \REGISTERS[26][9] , \REGISTERS[26][8] , \REGISTERS[26][7] ,
         \REGISTERS[26][6] , \REGISTERS[26][5] , \REGISTERS[26][4] ,
         \REGISTERS[26][3] , \REGISTERS[26][2] , \REGISTERS[26][1] ,
         \REGISTERS[26][0] , \REGISTERS[27][31] , \REGISTERS[27][30] ,
         \REGISTERS[27][29] , \REGISTERS[27][28] , \REGISTERS[27][27] ,
         \REGISTERS[27][26] , \REGISTERS[27][25] , \REGISTERS[27][24] ,
         \REGISTERS[27][23] , \REGISTERS[27][22] , \REGISTERS[27][21] ,
         \REGISTERS[27][20] , \REGISTERS[27][19] , \REGISTERS[27][18] ,
         \REGISTERS[27][17] , \REGISTERS[27][16] , \REGISTERS[27][15] ,
         \REGISTERS[27][14] , \REGISTERS[27][13] , \REGISTERS[27][12] ,
         \REGISTERS[27][11] , \REGISTERS[27][10] , \REGISTERS[27][9] ,
         \REGISTERS[27][8] , \REGISTERS[27][7] , \REGISTERS[27][6] ,
         \REGISTERS[27][5] , \REGISTERS[27][4] , \REGISTERS[27][3] ,
         \REGISTERS[27][2] , \REGISTERS[27][1] , \REGISTERS[27][0] ,
         \REGISTERS[28][31] , \REGISTERS[28][30] , \REGISTERS[28][29] ,
         \REGISTERS[28][28] , \REGISTERS[28][27] , \REGISTERS[28][26] ,
         \REGISTERS[28][25] , \REGISTERS[28][24] , \REGISTERS[28][23] ,
         \REGISTERS[28][22] , \REGISTERS[28][21] , \REGISTERS[28][20] ,
         \REGISTERS[28][19] , \REGISTERS[28][18] , \REGISTERS[28][17] ,
         \REGISTERS[28][16] , \REGISTERS[28][15] , \REGISTERS[28][14] ,
         \REGISTERS[28][13] , \REGISTERS[28][12] , \REGISTERS[28][11] ,
         \REGISTERS[28][10] , \REGISTERS[28][9] , \REGISTERS[28][8] ,
         \REGISTERS[28][7] , \REGISTERS[28][6] , \REGISTERS[28][5] ,
         \REGISTERS[28][4] , \REGISTERS[28][3] , \REGISTERS[28][2] ,
         \REGISTERS[28][1] , \REGISTERS[28][0] , \REGISTERS[29][31] ,
         \REGISTERS[29][30] , \REGISTERS[29][29] , \REGISTERS[29][28] ,
         \REGISTERS[29][27] , \REGISTERS[29][26] , \REGISTERS[29][25] ,
         \REGISTERS[29][24] , \REGISTERS[29][23] , \REGISTERS[29][22] ,
         \REGISTERS[29][21] , \REGISTERS[29][20] , \REGISTERS[29][19] ,
         \REGISTERS[29][18] , \REGISTERS[29][17] , \REGISTERS[29][16] ,
         \REGISTERS[29][15] , \REGISTERS[29][14] , \REGISTERS[29][13] ,
         \REGISTERS[29][12] , \REGISTERS[29][11] , \REGISTERS[29][10] ,
         \REGISTERS[29][9] , \REGISTERS[29][8] , \REGISTERS[29][7] ,
         \REGISTERS[29][6] , \REGISTERS[29][5] , \REGISTERS[29][4] ,
         \REGISTERS[29][3] , \REGISTERS[29][2] , \REGISTERS[29][1] ,
         \REGISTERS[29][0] , \REGISTERS[30][31] , \REGISTERS[30][30] ,
         \REGISTERS[30][29] , \REGISTERS[30][28] , \REGISTERS[30][27] ,
         \REGISTERS[30][26] , \REGISTERS[30][25] , \REGISTERS[30][24] ,
         \REGISTERS[30][23] , \REGISTERS[30][22] , \REGISTERS[30][21] ,
         \REGISTERS[30][20] , \REGISTERS[30][19] , \REGISTERS[30][18] ,
         \REGISTERS[30][17] , \REGISTERS[30][16] , \REGISTERS[30][15] ,
         \REGISTERS[30][14] , \REGISTERS[30][13] , \REGISTERS[30][12] ,
         \REGISTERS[30][11] , \REGISTERS[30][10] , \REGISTERS[30][9] ,
         \REGISTERS[30][8] , \REGISTERS[30][7] , \REGISTERS[30][6] ,
         \REGISTERS[30][5] , \REGISTERS[30][4] , \REGISTERS[30][3] ,
         \REGISTERS[30][2] , \REGISTERS[30][1] , \REGISTERS[30][0] ,
         \REGISTERS[31][31] , \REGISTERS[31][30] , \REGISTERS[31][29] ,
         \REGISTERS[31][28] , \REGISTERS[31][27] , \REGISTERS[31][26] ,
         \REGISTERS[31][25] , \REGISTERS[31][24] , \REGISTERS[31][23] ,
         \REGISTERS[31][22] , \REGISTERS[31][21] , \REGISTERS[31][20] ,
         \REGISTERS[31][19] , \REGISTERS[31][18] , \REGISTERS[31][17] ,
         \REGISTERS[31][16] , \REGISTERS[31][15] , \REGISTERS[31][14] ,
         \REGISTERS[31][13] , \REGISTERS[31][12] , \REGISTERS[31][11] ,
         \REGISTERS[31][10] , \REGISTERS[31][9] , \REGISTERS[31][8] ,
         \REGISTERS[31][7] , \REGISTERS[31][6] , \REGISTERS[31][5] ,
         \REGISTERS[31][4] , \REGISTERS[31][3] , \REGISTERS[31][2] ,
         \REGISTERS[31][1] , \REGISTERS[31][0] , N2163, N2227, N2291, N2355,
         N2419, N2483, N2547, N2611, N2675, N2739, N2803, N2867, N2931, N2995,
         N3059, N3123, N3187, N3251, N3315, N3379, N3443, N3507, N3571, N3635,
         N3699, N3763, N3827, N3891, N3955, N4019, N4083, N4086, N4088, N4090,
         N4092, N4094, N4096, N4098, N4100, N4102, N4104, N4106, N4108, N4110,
         N4112, N4114, N4116, N4118, N4120, N4122, N4124, N4126, N4128, N4130,
         N4132, N4134, N4136, N4138, N4140, N4142, N4144, N4146, N4148, N4215,
         N4216, N4217, N4218, N4219, N4220, N4221, N4222, N4223, N4224, N4225,
         N4226, N4227, N4228, N4229, N4230, N4231, N4232, N4233, N4234, N4235,
         N4236, N4237, N4238, N4239, N4240, N4241, N4242, N4243, N4244, N4245,
         N4246, N4278, N4344, N4345, N4346, N4347, N4348, N4349, N4350, N4351,
         N4352, N4353, N4354, N4355, N4356, N4357, N4358, N4359, N4360, N4361,
         N4362, N4363, N4364, N4365, N4366, N4367, N4368, N4369, N4370, N4371,
         N4372, N4373, N4374, N4375, N4407, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1,
         n193, n227, n261, n295, n329;

  DLH_X1 \REGISTERS_reg[1][31]  ( .G(N4083), .D(N4148), .Q(\REGISTERS[1][31] )
         );
  DLH_X1 \REGISTERS_reg[1][30]  ( .G(N4083), .D(N4146), .Q(\REGISTERS[1][30] )
         );
  DLH_X1 \REGISTERS_reg[1][29]  ( .G(N4083), .D(N4144), .Q(\REGISTERS[1][29] )
         );
  DLH_X1 \REGISTERS_reg[1][28]  ( .G(N4083), .D(N4142), .Q(\REGISTERS[1][28] )
         );
  DLH_X1 \REGISTERS_reg[1][27]  ( .G(N4083), .D(N4140), .Q(\REGISTERS[1][27] )
         );
  DLH_X1 \REGISTERS_reg[1][26]  ( .G(N4083), .D(N4138), .Q(\REGISTERS[1][26] )
         );
  DLH_X1 \REGISTERS_reg[1][25]  ( .G(N4083), .D(N4136), .Q(\REGISTERS[1][25] )
         );
  DLH_X1 \REGISTERS_reg[1][24]  ( .G(N4083), .D(N4134), .Q(\REGISTERS[1][24] )
         );
  DLH_X1 \REGISTERS_reg[1][23]  ( .G(N4083), .D(N4132), .Q(\REGISTERS[1][23] )
         );
  DLH_X1 \REGISTERS_reg[1][22]  ( .G(N4083), .D(N4130), .Q(\REGISTERS[1][22] )
         );
  DLH_X1 \REGISTERS_reg[1][21]  ( .G(N4083), .D(N4128), .Q(\REGISTERS[1][21] )
         );
  DLH_X1 \REGISTERS_reg[1][20]  ( .G(N4083), .D(N4126), .Q(\REGISTERS[1][20] )
         );
  DLH_X1 \REGISTERS_reg[1][19]  ( .G(N4083), .D(N4124), .Q(\REGISTERS[1][19] )
         );
  DLH_X1 \REGISTERS_reg[1][18]  ( .G(N4083), .D(N4122), .Q(\REGISTERS[1][18] )
         );
  DLH_X1 \REGISTERS_reg[1][17]  ( .G(N4083), .D(N4120), .Q(\REGISTERS[1][17] )
         );
  DLH_X1 \REGISTERS_reg[1][16]  ( .G(N4083), .D(N4118), .Q(\REGISTERS[1][16] )
         );
  DLH_X1 \REGISTERS_reg[1][15]  ( .G(N4083), .D(N4116), .Q(\REGISTERS[1][15] )
         );
  DLH_X1 \REGISTERS_reg[1][14]  ( .G(N4083), .D(N4114), .Q(\REGISTERS[1][14] )
         );
  DLH_X1 \REGISTERS_reg[1][13]  ( .G(N4083), .D(N4112), .Q(\REGISTERS[1][13] )
         );
  DLH_X1 \REGISTERS_reg[1][12]  ( .G(N4083), .D(N4110), .Q(\REGISTERS[1][12] )
         );
  DLH_X1 \REGISTERS_reg[1][11]  ( .G(N4083), .D(N4108), .Q(\REGISTERS[1][11] )
         );
  DLH_X1 \REGISTERS_reg[1][10]  ( .G(N4083), .D(N4106), .Q(\REGISTERS[1][10] )
         );
  DLH_X1 \REGISTERS_reg[1][9]  ( .G(N4083), .D(N4104), .Q(\REGISTERS[1][9] )
         );
  DLH_X1 \REGISTERS_reg[1][8]  ( .G(N4083), .D(N4102), .Q(\REGISTERS[1][8] )
         );
  DLH_X1 \REGISTERS_reg[1][7]  ( .G(N4083), .D(N4100), .Q(\REGISTERS[1][7] )
         );
  DLH_X1 \REGISTERS_reg[1][6]  ( .G(N4083), .D(N4098), .Q(\REGISTERS[1][6] )
         );
  DLH_X1 \REGISTERS_reg[1][5]  ( .G(N4083), .D(N4096), .Q(\REGISTERS[1][5] )
         );
  DLH_X1 \REGISTERS_reg[1][4]  ( .G(N4083), .D(N4094), .Q(\REGISTERS[1][4] )
         );
  DLH_X1 \REGISTERS_reg[1][3]  ( .G(N4083), .D(N4092), .Q(\REGISTERS[1][3] )
         );
  DLH_X1 \REGISTERS_reg[1][2]  ( .G(N4083), .D(N4090), .Q(\REGISTERS[1][2] )
         );
  DLH_X1 \REGISTERS_reg[1][1]  ( .G(N4083), .D(N4088), .Q(\REGISTERS[1][1] )
         );
  DLH_X1 \REGISTERS_reg[1][0]  ( .G(N4083), .D(N4086), .Q(\REGISTERS[1][0] )
         );
  DLH_X1 \REGISTERS_reg[2][31]  ( .G(N4019), .D(N4148), .Q(\REGISTERS[2][31] )
         );
  DLH_X1 \REGISTERS_reg[2][30]  ( .G(N4019), .D(N4146), .Q(\REGISTERS[2][30] )
         );
  DLH_X1 \REGISTERS_reg[2][29]  ( .G(N4019), .D(N4144), .Q(\REGISTERS[2][29] )
         );
  DLH_X1 \REGISTERS_reg[2][28]  ( .G(N4019), .D(N4142), .Q(\REGISTERS[2][28] )
         );
  DLH_X1 \REGISTERS_reg[2][27]  ( .G(N4019), .D(N4140), .Q(\REGISTERS[2][27] )
         );
  DLH_X1 \REGISTERS_reg[2][26]  ( .G(N4019), .D(N4138), .Q(\REGISTERS[2][26] )
         );
  DLH_X1 \REGISTERS_reg[2][25]  ( .G(N4019), .D(N4136), .Q(\REGISTERS[2][25] )
         );
  DLH_X1 \REGISTERS_reg[2][24]  ( .G(N4019), .D(N4134), .Q(\REGISTERS[2][24] )
         );
  DLH_X1 \REGISTERS_reg[2][23]  ( .G(N4019), .D(N4132), .Q(\REGISTERS[2][23] )
         );
  DLH_X1 \REGISTERS_reg[2][22]  ( .G(N4019), .D(N4130), .Q(\REGISTERS[2][22] )
         );
  DLH_X1 \REGISTERS_reg[2][21]  ( .G(N4019), .D(N4128), .Q(\REGISTERS[2][21] )
         );
  DLH_X1 \REGISTERS_reg[2][20]  ( .G(N4019), .D(N4126), .Q(\REGISTERS[2][20] )
         );
  DLH_X1 \REGISTERS_reg[2][19]  ( .G(N4019), .D(N4124), .Q(\REGISTERS[2][19] )
         );
  DLH_X1 \REGISTERS_reg[2][18]  ( .G(N4019), .D(N4122), .Q(\REGISTERS[2][18] )
         );
  DLH_X1 \REGISTERS_reg[2][17]  ( .G(N4019), .D(N4120), .Q(\REGISTERS[2][17] )
         );
  DLH_X1 \REGISTERS_reg[2][16]  ( .G(N4019), .D(N4118), .Q(\REGISTERS[2][16] )
         );
  DLH_X1 \REGISTERS_reg[2][15]  ( .G(N4019), .D(N4116), .Q(\REGISTERS[2][15] )
         );
  DLH_X1 \REGISTERS_reg[2][14]  ( .G(N4019), .D(N4114), .Q(\REGISTERS[2][14] )
         );
  DLH_X1 \REGISTERS_reg[2][13]  ( .G(N4019), .D(N4112), .Q(\REGISTERS[2][13] )
         );
  DLH_X1 \REGISTERS_reg[2][12]  ( .G(N4019), .D(N4110), .Q(\REGISTERS[2][12] )
         );
  DLH_X1 \REGISTERS_reg[2][11]  ( .G(N4019), .D(N4108), .Q(\REGISTERS[2][11] )
         );
  DLH_X1 \REGISTERS_reg[2][10]  ( .G(N4019), .D(N4106), .Q(\REGISTERS[2][10] )
         );
  DLH_X1 \REGISTERS_reg[2][9]  ( .G(N4019), .D(N4104), .Q(\REGISTERS[2][9] )
         );
  DLH_X1 \REGISTERS_reg[2][8]  ( .G(N4019), .D(N4102), .Q(\REGISTERS[2][8] )
         );
  DLH_X1 \REGISTERS_reg[2][7]  ( .G(N4019), .D(N4100), .Q(\REGISTERS[2][7] )
         );
  DLH_X1 \REGISTERS_reg[2][6]  ( .G(N4019), .D(N4098), .Q(\REGISTERS[2][6] )
         );
  DLH_X1 \REGISTERS_reg[2][5]  ( .G(N4019), .D(N4096), .Q(\REGISTERS[2][5] )
         );
  DLH_X1 \REGISTERS_reg[2][4]  ( .G(N4019), .D(N4094), .Q(\REGISTERS[2][4] )
         );
  DLH_X1 \REGISTERS_reg[2][3]  ( .G(N4019), .D(N4092), .Q(\REGISTERS[2][3] )
         );
  DLH_X1 \REGISTERS_reg[2][2]  ( .G(N4019), .D(N4090), .Q(\REGISTERS[2][2] )
         );
  DLH_X1 \REGISTERS_reg[2][1]  ( .G(N4019), .D(N4088), .Q(\REGISTERS[2][1] )
         );
  DLH_X1 \REGISTERS_reg[2][0]  ( .G(N4019), .D(N4086), .Q(\REGISTERS[2][0] )
         );
  DLH_X1 \REGISTERS_reg[3][31]  ( .G(N3955), .D(N4148), .Q(\REGISTERS[3][31] )
         );
  DLH_X1 \REGISTERS_reg[3][30]  ( .G(N3955), .D(N4146), .Q(\REGISTERS[3][30] )
         );
  DLH_X1 \REGISTERS_reg[3][29]  ( .G(N3955), .D(N4144), .Q(\REGISTERS[3][29] )
         );
  DLH_X1 \REGISTERS_reg[3][28]  ( .G(N3955), .D(N4142), .Q(\REGISTERS[3][28] )
         );
  DLH_X1 \REGISTERS_reg[3][27]  ( .G(N3955), .D(N4140), .Q(\REGISTERS[3][27] )
         );
  DLH_X1 \REGISTERS_reg[3][26]  ( .G(N3955), .D(N4138), .Q(\REGISTERS[3][26] )
         );
  DLH_X1 \REGISTERS_reg[3][25]  ( .G(N3955), .D(N4136), .Q(\REGISTERS[3][25] )
         );
  DLH_X1 \REGISTERS_reg[3][24]  ( .G(N3955), .D(N4134), .Q(\REGISTERS[3][24] )
         );
  DLH_X1 \REGISTERS_reg[3][23]  ( .G(N3955), .D(N4132), .Q(\REGISTERS[3][23] )
         );
  DLH_X1 \REGISTERS_reg[3][22]  ( .G(N3955), .D(N4130), .Q(\REGISTERS[3][22] )
         );
  DLH_X1 \REGISTERS_reg[3][21]  ( .G(N3955), .D(N4128), .Q(\REGISTERS[3][21] )
         );
  DLH_X1 \REGISTERS_reg[3][20]  ( .G(N3955), .D(N4126), .Q(\REGISTERS[3][20] )
         );
  DLH_X1 \REGISTERS_reg[3][19]  ( .G(N3955), .D(N4124), .Q(\REGISTERS[3][19] )
         );
  DLH_X1 \REGISTERS_reg[3][18]  ( .G(N3955), .D(N4122), .Q(\REGISTERS[3][18] )
         );
  DLH_X1 \REGISTERS_reg[3][17]  ( .G(N3955), .D(N4120), .Q(\REGISTERS[3][17] )
         );
  DLH_X1 \REGISTERS_reg[3][16]  ( .G(N3955), .D(N4118), .Q(\REGISTERS[3][16] )
         );
  DLH_X1 \REGISTERS_reg[3][15]  ( .G(N3955), .D(N4116), .Q(\REGISTERS[3][15] )
         );
  DLH_X1 \REGISTERS_reg[3][14]  ( .G(N3955), .D(N4114), .Q(\REGISTERS[3][14] )
         );
  DLH_X1 \REGISTERS_reg[3][13]  ( .G(N3955), .D(N4112), .Q(\REGISTERS[3][13] )
         );
  DLH_X1 \REGISTERS_reg[3][12]  ( .G(N3955), .D(N4110), .Q(\REGISTERS[3][12] )
         );
  DLH_X1 \REGISTERS_reg[3][11]  ( .G(N3955), .D(N4108), .Q(\REGISTERS[3][11] )
         );
  DLH_X1 \REGISTERS_reg[3][10]  ( .G(N3955), .D(N4106), .Q(\REGISTERS[3][10] )
         );
  DLH_X1 \REGISTERS_reg[3][9]  ( .G(N3955), .D(N4104), .Q(\REGISTERS[3][9] )
         );
  DLH_X1 \REGISTERS_reg[3][8]  ( .G(N3955), .D(N4102), .Q(\REGISTERS[3][8] )
         );
  DLH_X1 \REGISTERS_reg[3][7]  ( .G(N3955), .D(N4100), .Q(\REGISTERS[3][7] )
         );
  DLH_X1 \REGISTERS_reg[3][6]  ( .G(N3955), .D(N4098), .Q(\REGISTERS[3][6] )
         );
  DLH_X1 \REGISTERS_reg[3][5]  ( .G(N3955), .D(N4096), .Q(\REGISTERS[3][5] )
         );
  DLH_X1 \REGISTERS_reg[3][4]  ( .G(N3955), .D(N4094), .Q(\REGISTERS[3][4] )
         );
  DLH_X1 \REGISTERS_reg[3][3]  ( .G(N3955), .D(N4092), .Q(\REGISTERS[3][3] )
         );
  DLH_X1 \REGISTERS_reg[3][2]  ( .G(N3955), .D(N4090), .Q(\REGISTERS[3][2] )
         );
  DLH_X1 \REGISTERS_reg[3][1]  ( .G(N3955), .D(N4088), .Q(\REGISTERS[3][1] )
         );
  DLH_X1 \REGISTERS_reg[3][0]  ( .G(N3955), .D(N4086), .Q(\REGISTERS[3][0] )
         );
  DLH_X1 \REGISTERS_reg[4][31]  ( .G(N3891), .D(N4148), .Q(\REGISTERS[4][31] )
         );
  DLH_X1 \REGISTERS_reg[4][30]  ( .G(N3891), .D(N4146), .Q(\REGISTERS[4][30] )
         );
  DLH_X1 \REGISTERS_reg[4][29]  ( .G(N3891), .D(N4144), .Q(\REGISTERS[4][29] )
         );
  DLH_X1 \REGISTERS_reg[4][28]  ( .G(N3891), .D(N4142), .Q(\REGISTERS[4][28] )
         );
  DLH_X1 \REGISTERS_reg[4][27]  ( .G(N3891), .D(N4140), .Q(\REGISTERS[4][27] )
         );
  DLH_X1 \REGISTERS_reg[4][26]  ( .G(N3891), .D(N4138), .Q(\REGISTERS[4][26] )
         );
  DLH_X1 \REGISTERS_reg[4][25]  ( .G(N3891), .D(N4136), .Q(\REGISTERS[4][25] )
         );
  DLH_X1 \REGISTERS_reg[4][24]  ( .G(N3891), .D(N4134), .Q(\REGISTERS[4][24] )
         );
  DLH_X1 \REGISTERS_reg[4][23]  ( .G(N3891), .D(N4132), .Q(\REGISTERS[4][23] )
         );
  DLH_X1 \REGISTERS_reg[4][22]  ( .G(N3891), .D(N4130), .Q(\REGISTERS[4][22] )
         );
  DLH_X1 \REGISTERS_reg[4][21]  ( .G(N3891), .D(N4128), .Q(\REGISTERS[4][21] )
         );
  DLH_X1 \REGISTERS_reg[4][20]  ( .G(N3891), .D(N4126), .Q(\REGISTERS[4][20] )
         );
  DLH_X1 \REGISTERS_reg[4][19]  ( .G(N3891), .D(N4124), .Q(\REGISTERS[4][19] )
         );
  DLH_X1 \REGISTERS_reg[4][18]  ( .G(N3891), .D(N4122), .Q(\REGISTERS[4][18] )
         );
  DLH_X1 \REGISTERS_reg[4][17]  ( .G(N3891), .D(N4120), .Q(\REGISTERS[4][17] )
         );
  DLH_X1 \REGISTERS_reg[4][16]  ( .G(N3891), .D(N4118), .Q(\REGISTERS[4][16] )
         );
  DLH_X1 \REGISTERS_reg[4][15]  ( .G(N3891), .D(N4116), .Q(\REGISTERS[4][15] )
         );
  DLH_X1 \REGISTERS_reg[4][14]  ( .G(N3891), .D(N4114), .Q(\REGISTERS[4][14] )
         );
  DLH_X1 \REGISTERS_reg[4][13]  ( .G(N3891), .D(N4112), .Q(\REGISTERS[4][13] )
         );
  DLH_X1 \REGISTERS_reg[4][12]  ( .G(N3891), .D(N4110), .Q(\REGISTERS[4][12] )
         );
  DLH_X1 \REGISTERS_reg[4][11]  ( .G(N3891), .D(N4108), .Q(\REGISTERS[4][11] )
         );
  DLH_X1 \REGISTERS_reg[4][10]  ( .G(N3891), .D(N4106), .Q(\REGISTERS[4][10] )
         );
  DLH_X1 \REGISTERS_reg[4][9]  ( .G(N3891), .D(N4104), .Q(\REGISTERS[4][9] )
         );
  DLH_X1 \REGISTERS_reg[4][8]  ( .G(N3891), .D(N4102), .Q(\REGISTERS[4][8] )
         );
  DLH_X1 \REGISTERS_reg[4][7]  ( .G(N3891), .D(N4100), .Q(\REGISTERS[4][7] )
         );
  DLH_X1 \REGISTERS_reg[4][6]  ( .G(N3891), .D(N4098), .Q(\REGISTERS[4][6] )
         );
  DLH_X1 \REGISTERS_reg[4][5]  ( .G(N3891), .D(N4096), .Q(\REGISTERS[4][5] )
         );
  DLH_X1 \REGISTERS_reg[4][4]  ( .G(N3891), .D(N4094), .Q(\REGISTERS[4][4] )
         );
  DLH_X1 \REGISTERS_reg[4][3]  ( .G(N3891), .D(N4092), .Q(\REGISTERS[4][3] )
         );
  DLH_X1 \REGISTERS_reg[4][2]  ( .G(N3891), .D(N4090), .Q(\REGISTERS[4][2] )
         );
  DLH_X1 \REGISTERS_reg[4][1]  ( .G(N3891), .D(N4088), .Q(\REGISTERS[4][1] )
         );
  DLH_X1 \REGISTERS_reg[4][0]  ( .G(N3891), .D(N4086), .Q(\REGISTERS[4][0] )
         );
  DLH_X1 \REGISTERS_reg[5][31]  ( .G(N3827), .D(N4148), .Q(\REGISTERS[5][31] )
         );
  DLH_X1 \REGISTERS_reg[5][30]  ( .G(N3827), .D(N4146), .Q(\REGISTERS[5][30] )
         );
  DLH_X1 \REGISTERS_reg[5][29]  ( .G(N3827), .D(N4144), .Q(\REGISTERS[5][29] )
         );
  DLH_X1 \REGISTERS_reg[5][28]  ( .G(N3827), .D(N4142), .Q(\REGISTERS[5][28] )
         );
  DLH_X1 \REGISTERS_reg[5][27]  ( .G(N3827), .D(N4140), .Q(\REGISTERS[5][27] )
         );
  DLH_X1 \REGISTERS_reg[5][26]  ( .G(N3827), .D(N4138), .Q(\REGISTERS[5][26] )
         );
  DLH_X1 \REGISTERS_reg[5][25]  ( .G(N3827), .D(N4136), .Q(\REGISTERS[5][25] )
         );
  DLH_X1 \REGISTERS_reg[5][24]  ( .G(N3827), .D(N4134), .Q(\REGISTERS[5][24] )
         );
  DLH_X1 \REGISTERS_reg[5][23]  ( .G(N3827), .D(N4132), .Q(\REGISTERS[5][23] )
         );
  DLH_X1 \REGISTERS_reg[5][22]  ( .G(N3827), .D(N4130), .Q(\REGISTERS[5][22] )
         );
  DLH_X1 \REGISTERS_reg[5][21]  ( .G(N3827), .D(N4128), .Q(\REGISTERS[5][21] )
         );
  DLH_X1 \REGISTERS_reg[5][20]  ( .G(N3827), .D(N4126), .Q(\REGISTERS[5][20] )
         );
  DLH_X1 \REGISTERS_reg[5][19]  ( .G(N3827), .D(N4124), .Q(\REGISTERS[5][19] )
         );
  DLH_X1 \REGISTERS_reg[5][18]  ( .G(N3827), .D(N4122), .Q(\REGISTERS[5][18] )
         );
  DLH_X1 \REGISTERS_reg[5][17]  ( .G(N3827), .D(N4120), .Q(\REGISTERS[5][17] )
         );
  DLH_X1 \REGISTERS_reg[5][16]  ( .G(N3827), .D(N4118), .Q(\REGISTERS[5][16] )
         );
  DLH_X1 \REGISTERS_reg[5][15]  ( .G(N3827), .D(N4116), .Q(\REGISTERS[5][15] )
         );
  DLH_X1 \REGISTERS_reg[5][14]  ( .G(N3827), .D(N4114), .Q(\REGISTERS[5][14] )
         );
  DLH_X1 \REGISTERS_reg[5][13]  ( .G(N3827), .D(N4112), .Q(\REGISTERS[5][13] )
         );
  DLH_X1 \REGISTERS_reg[5][12]  ( .G(N3827), .D(N4110), .Q(\REGISTERS[5][12] )
         );
  DLH_X1 \REGISTERS_reg[5][11]  ( .G(N3827), .D(N4108), .Q(\REGISTERS[5][11] )
         );
  DLH_X1 \REGISTERS_reg[5][10]  ( .G(N3827), .D(N4106), .Q(\REGISTERS[5][10] )
         );
  DLH_X1 \REGISTERS_reg[5][9]  ( .G(N3827), .D(N4104), .Q(\REGISTERS[5][9] )
         );
  DLH_X1 \REGISTERS_reg[5][8]  ( .G(N3827), .D(N4102), .Q(\REGISTERS[5][8] )
         );
  DLH_X1 \REGISTERS_reg[5][7]  ( .G(N3827), .D(N4100), .Q(\REGISTERS[5][7] )
         );
  DLH_X1 \REGISTERS_reg[5][6]  ( .G(N3827), .D(N4098), .Q(\REGISTERS[5][6] )
         );
  DLH_X1 \REGISTERS_reg[5][5]  ( .G(N3827), .D(N4096), .Q(\REGISTERS[5][5] )
         );
  DLH_X1 \REGISTERS_reg[5][4]  ( .G(N3827), .D(N4094), .Q(\REGISTERS[5][4] )
         );
  DLH_X1 \REGISTERS_reg[5][3]  ( .G(N3827), .D(N4092), .Q(\REGISTERS[5][3] )
         );
  DLH_X1 \REGISTERS_reg[5][2]  ( .G(N3827), .D(N4090), .Q(\REGISTERS[5][2] )
         );
  DLH_X1 \REGISTERS_reg[5][1]  ( .G(N3827), .D(N4088), .Q(\REGISTERS[5][1] )
         );
  DLH_X1 \REGISTERS_reg[5][0]  ( .G(N3827), .D(N4086), .Q(\REGISTERS[5][0] )
         );
  DLH_X1 \REGISTERS_reg[6][31]  ( .G(N3763), .D(N4148), .Q(\REGISTERS[6][31] )
         );
  DLH_X1 \REGISTERS_reg[6][30]  ( .G(N3763), .D(N4146), .Q(\REGISTERS[6][30] )
         );
  DLH_X1 \REGISTERS_reg[6][29]  ( .G(N3763), .D(N4144), .Q(\REGISTERS[6][29] )
         );
  DLH_X1 \REGISTERS_reg[6][28]  ( .G(N3763), .D(N4142), .Q(\REGISTERS[6][28] )
         );
  DLH_X1 \REGISTERS_reg[6][27]  ( .G(N3763), .D(N4140), .Q(\REGISTERS[6][27] )
         );
  DLH_X1 \REGISTERS_reg[6][26]  ( .G(N3763), .D(N4138), .Q(\REGISTERS[6][26] )
         );
  DLH_X1 \REGISTERS_reg[6][25]  ( .G(N3763), .D(N4136), .Q(\REGISTERS[6][25] )
         );
  DLH_X1 \REGISTERS_reg[6][24]  ( .G(N3763), .D(N4134), .Q(\REGISTERS[6][24] )
         );
  DLH_X1 \REGISTERS_reg[6][23]  ( .G(N3763), .D(N4132), .Q(\REGISTERS[6][23] )
         );
  DLH_X1 \REGISTERS_reg[6][22]  ( .G(N3763), .D(N4130), .Q(\REGISTERS[6][22] )
         );
  DLH_X1 \REGISTERS_reg[6][21]  ( .G(N3763), .D(N4128), .Q(\REGISTERS[6][21] )
         );
  DLH_X1 \REGISTERS_reg[6][20]  ( .G(N3763), .D(N4126), .Q(\REGISTERS[6][20] )
         );
  DLH_X1 \REGISTERS_reg[6][19]  ( .G(N3763), .D(N4124), .Q(\REGISTERS[6][19] )
         );
  DLH_X1 \REGISTERS_reg[6][18]  ( .G(N3763), .D(N4122), .Q(\REGISTERS[6][18] )
         );
  DLH_X1 \REGISTERS_reg[6][17]  ( .G(N3763), .D(N4120), .Q(\REGISTERS[6][17] )
         );
  DLH_X1 \REGISTERS_reg[6][16]  ( .G(N3763), .D(N4118), .Q(\REGISTERS[6][16] )
         );
  DLH_X1 \REGISTERS_reg[6][15]  ( .G(N3763), .D(N4116), .Q(\REGISTERS[6][15] )
         );
  DLH_X1 \REGISTERS_reg[6][14]  ( .G(N3763), .D(N4114), .Q(\REGISTERS[6][14] )
         );
  DLH_X1 \REGISTERS_reg[6][13]  ( .G(N3763), .D(N4112), .Q(\REGISTERS[6][13] )
         );
  DLH_X1 \REGISTERS_reg[6][12]  ( .G(N3763), .D(N4110), .Q(\REGISTERS[6][12] )
         );
  DLH_X1 \REGISTERS_reg[6][11]  ( .G(N3763), .D(N4108), .Q(\REGISTERS[6][11] )
         );
  DLH_X1 \REGISTERS_reg[6][10]  ( .G(N3763), .D(N4106), .Q(\REGISTERS[6][10] )
         );
  DLH_X1 \REGISTERS_reg[6][9]  ( .G(N3763), .D(N4104), .Q(\REGISTERS[6][9] )
         );
  DLH_X1 \REGISTERS_reg[6][8]  ( .G(N3763), .D(N4102), .Q(\REGISTERS[6][8] )
         );
  DLH_X1 \REGISTERS_reg[6][7]  ( .G(N3763), .D(N4100), .Q(\REGISTERS[6][7] )
         );
  DLH_X1 \REGISTERS_reg[6][6]  ( .G(N3763), .D(N4098), .Q(\REGISTERS[6][6] )
         );
  DLH_X1 \REGISTERS_reg[6][5]  ( .G(N3763), .D(N4096), .Q(\REGISTERS[6][5] )
         );
  DLH_X1 \REGISTERS_reg[6][4]  ( .G(N3763), .D(N4094), .Q(\REGISTERS[6][4] )
         );
  DLH_X1 \REGISTERS_reg[6][3]  ( .G(N3763), .D(N4092), .Q(\REGISTERS[6][3] )
         );
  DLH_X1 \REGISTERS_reg[6][2]  ( .G(N3763), .D(N4090), .Q(\REGISTERS[6][2] )
         );
  DLH_X1 \REGISTERS_reg[6][1]  ( .G(N3763), .D(N4088), .Q(\REGISTERS[6][1] )
         );
  DLH_X1 \REGISTERS_reg[6][0]  ( .G(N3763), .D(N4086), .Q(\REGISTERS[6][0] )
         );
  DLH_X1 \REGISTERS_reg[7][31]  ( .G(N3699), .D(N4148), .Q(\REGISTERS[7][31] )
         );
  DLH_X1 \REGISTERS_reg[7][30]  ( .G(N3699), .D(N4146), .Q(\REGISTERS[7][30] )
         );
  DLH_X1 \REGISTERS_reg[7][29]  ( .G(N3699), .D(N4144), .Q(\REGISTERS[7][29] )
         );
  DLH_X1 \REGISTERS_reg[7][28]  ( .G(N3699), .D(N4142), .Q(\REGISTERS[7][28] )
         );
  DLH_X1 \REGISTERS_reg[7][27]  ( .G(N3699), .D(N4140), .Q(\REGISTERS[7][27] )
         );
  DLH_X1 \REGISTERS_reg[7][26]  ( .G(N3699), .D(N4138), .Q(\REGISTERS[7][26] )
         );
  DLH_X1 \REGISTERS_reg[7][25]  ( .G(N3699), .D(N4136), .Q(\REGISTERS[7][25] )
         );
  DLH_X1 \REGISTERS_reg[7][24]  ( .G(N3699), .D(N4134), .Q(\REGISTERS[7][24] )
         );
  DLH_X1 \REGISTERS_reg[7][23]  ( .G(N3699), .D(N4132), .Q(\REGISTERS[7][23] )
         );
  DLH_X1 \REGISTERS_reg[7][22]  ( .G(N3699), .D(N4130), .Q(\REGISTERS[7][22] )
         );
  DLH_X1 \REGISTERS_reg[7][21]  ( .G(N3699), .D(N4128), .Q(\REGISTERS[7][21] )
         );
  DLH_X1 \REGISTERS_reg[7][20]  ( .G(N3699), .D(N4126), .Q(\REGISTERS[7][20] )
         );
  DLH_X1 \REGISTERS_reg[7][19]  ( .G(N3699), .D(N4124), .Q(\REGISTERS[7][19] )
         );
  DLH_X1 \REGISTERS_reg[7][18]  ( .G(N3699), .D(N4122), .Q(\REGISTERS[7][18] )
         );
  DLH_X1 \REGISTERS_reg[7][17]  ( .G(N3699), .D(N4120), .Q(\REGISTERS[7][17] )
         );
  DLH_X1 \REGISTERS_reg[7][16]  ( .G(N3699), .D(N4118), .Q(\REGISTERS[7][16] )
         );
  DLH_X1 \REGISTERS_reg[7][15]  ( .G(N3699), .D(N4116), .Q(\REGISTERS[7][15] )
         );
  DLH_X1 \REGISTERS_reg[7][14]  ( .G(N3699), .D(N4114), .Q(\REGISTERS[7][14] )
         );
  DLH_X1 \REGISTERS_reg[7][13]  ( .G(N3699), .D(N4112), .Q(\REGISTERS[7][13] )
         );
  DLH_X1 \REGISTERS_reg[7][12]  ( .G(N3699), .D(N4110), .Q(\REGISTERS[7][12] )
         );
  DLH_X1 \REGISTERS_reg[7][11]  ( .G(N3699), .D(N4108), .Q(\REGISTERS[7][11] )
         );
  DLH_X1 \REGISTERS_reg[7][10]  ( .G(N3699), .D(N4106), .Q(\REGISTERS[7][10] )
         );
  DLH_X1 \REGISTERS_reg[7][9]  ( .G(N3699), .D(N4104), .Q(\REGISTERS[7][9] )
         );
  DLH_X1 \REGISTERS_reg[7][8]  ( .G(N3699), .D(N4102), .Q(\REGISTERS[7][8] )
         );
  DLH_X1 \REGISTERS_reg[7][7]  ( .G(N3699), .D(N4100), .Q(\REGISTERS[7][7] )
         );
  DLH_X1 \REGISTERS_reg[7][6]  ( .G(N3699), .D(N4098), .Q(\REGISTERS[7][6] )
         );
  DLH_X1 \REGISTERS_reg[7][5]  ( .G(N3699), .D(N4096), .Q(\REGISTERS[7][5] )
         );
  DLH_X1 \REGISTERS_reg[7][4]  ( .G(N3699), .D(N4094), .Q(\REGISTERS[7][4] )
         );
  DLH_X1 \REGISTERS_reg[7][3]  ( .G(N3699), .D(N4092), .Q(\REGISTERS[7][3] )
         );
  DLH_X1 \REGISTERS_reg[7][2]  ( .G(N3699), .D(N4090), .Q(\REGISTERS[7][2] )
         );
  DLH_X1 \REGISTERS_reg[7][1]  ( .G(N3699), .D(N4088), .Q(\REGISTERS[7][1] )
         );
  DLH_X1 \REGISTERS_reg[7][0]  ( .G(N3699), .D(N4086), .Q(\REGISTERS[7][0] )
         );
  DLH_X1 \REGISTERS_reg[8][31]  ( .G(N3635), .D(N4148), .Q(\REGISTERS[8][31] )
         );
  DLH_X1 \REGISTERS_reg[8][30]  ( .G(N3635), .D(N4146), .Q(\REGISTERS[8][30] )
         );
  DLH_X1 \REGISTERS_reg[8][29]  ( .G(N3635), .D(N4144), .Q(\REGISTERS[8][29] )
         );
  DLH_X1 \REGISTERS_reg[8][28]  ( .G(N3635), .D(N4142), .Q(\REGISTERS[8][28] )
         );
  DLH_X1 \REGISTERS_reg[8][27]  ( .G(N3635), .D(N4140), .Q(\REGISTERS[8][27] )
         );
  DLH_X1 \REGISTERS_reg[8][26]  ( .G(N3635), .D(N4138), .Q(\REGISTERS[8][26] )
         );
  DLH_X1 \REGISTERS_reg[8][25]  ( .G(N3635), .D(N4136), .Q(\REGISTERS[8][25] )
         );
  DLH_X1 \REGISTERS_reg[8][24]  ( .G(N3635), .D(N4134), .Q(\REGISTERS[8][24] )
         );
  DLH_X1 \REGISTERS_reg[8][23]  ( .G(N3635), .D(N4132), .Q(\REGISTERS[8][23] )
         );
  DLH_X1 \REGISTERS_reg[8][22]  ( .G(N3635), .D(N4130), .Q(\REGISTERS[8][22] )
         );
  DLH_X1 \REGISTERS_reg[8][21]  ( .G(N3635), .D(N4128), .Q(\REGISTERS[8][21] )
         );
  DLH_X1 \REGISTERS_reg[8][20]  ( .G(N3635), .D(N4126), .Q(\REGISTERS[8][20] )
         );
  DLH_X1 \REGISTERS_reg[8][19]  ( .G(N3635), .D(N4124), .Q(\REGISTERS[8][19] )
         );
  DLH_X1 \REGISTERS_reg[8][18]  ( .G(N3635), .D(N4122), .Q(\REGISTERS[8][18] )
         );
  DLH_X1 \REGISTERS_reg[8][17]  ( .G(N3635), .D(N4120), .Q(\REGISTERS[8][17] )
         );
  DLH_X1 \REGISTERS_reg[8][16]  ( .G(N3635), .D(N4118), .Q(\REGISTERS[8][16] )
         );
  DLH_X1 \REGISTERS_reg[8][15]  ( .G(N3635), .D(N4116), .Q(\REGISTERS[8][15] )
         );
  DLH_X1 \REGISTERS_reg[8][14]  ( .G(N3635), .D(N4114), .Q(\REGISTERS[8][14] )
         );
  DLH_X1 \REGISTERS_reg[8][13]  ( .G(N3635), .D(N4112), .Q(\REGISTERS[8][13] )
         );
  DLH_X1 \REGISTERS_reg[8][12]  ( .G(N3635), .D(N4110), .Q(\REGISTERS[8][12] )
         );
  DLH_X1 \REGISTERS_reg[8][11]  ( .G(N3635), .D(N4108), .Q(\REGISTERS[8][11] )
         );
  DLH_X1 \REGISTERS_reg[8][10]  ( .G(N3635), .D(N4106), .Q(\REGISTERS[8][10] )
         );
  DLH_X1 \REGISTERS_reg[8][9]  ( .G(N3635), .D(N4104), .Q(\REGISTERS[8][9] )
         );
  DLH_X1 \REGISTERS_reg[8][8]  ( .G(N3635), .D(N4102), .Q(\REGISTERS[8][8] )
         );
  DLH_X1 \REGISTERS_reg[8][7]  ( .G(N3635), .D(N4100), .Q(\REGISTERS[8][7] )
         );
  DLH_X1 \REGISTERS_reg[8][6]  ( .G(N3635), .D(N4098), .Q(\REGISTERS[8][6] )
         );
  DLH_X1 \REGISTERS_reg[8][5]  ( .G(N3635), .D(N4096), .Q(\REGISTERS[8][5] )
         );
  DLH_X1 \REGISTERS_reg[8][4]  ( .G(N3635), .D(N4094), .Q(\REGISTERS[8][4] )
         );
  DLH_X1 \REGISTERS_reg[8][3]  ( .G(N3635), .D(N4092), .Q(\REGISTERS[8][3] )
         );
  DLH_X1 \REGISTERS_reg[8][2]  ( .G(N3635), .D(N4090), .Q(\REGISTERS[8][2] )
         );
  DLH_X1 \REGISTERS_reg[8][1]  ( .G(N3635), .D(N4088), .Q(\REGISTERS[8][1] )
         );
  DLH_X1 \REGISTERS_reg[8][0]  ( .G(N3635), .D(N4086), .Q(\REGISTERS[8][0] )
         );
  DLH_X1 \REGISTERS_reg[9][31]  ( .G(N3571), .D(N4148), .Q(\REGISTERS[9][31] )
         );
  DLH_X1 \REGISTERS_reg[9][30]  ( .G(N3571), .D(N4146), .Q(\REGISTERS[9][30] )
         );
  DLH_X1 \REGISTERS_reg[9][29]  ( .G(N3571), .D(N4144), .Q(\REGISTERS[9][29] )
         );
  DLH_X1 \REGISTERS_reg[9][28]  ( .G(N3571), .D(N4142), .Q(\REGISTERS[9][28] )
         );
  DLH_X1 \REGISTERS_reg[9][27]  ( .G(N3571), .D(N4140), .Q(\REGISTERS[9][27] )
         );
  DLH_X1 \REGISTERS_reg[9][26]  ( .G(N3571), .D(N4138), .Q(\REGISTERS[9][26] )
         );
  DLH_X1 \REGISTERS_reg[9][25]  ( .G(N3571), .D(N4136), .Q(\REGISTERS[9][25] )
         );
  DLH_X1 \REGISTERS_reg[9][24]  ( .G(N3571), .D(N4134), .Q(\REGISTERS[9][24] )
         );
  DLH_X1 \REGISTERS_reg[9][23]  ( .G(N3571), .D(N4132), .Q(\REGISTERS[9][23] )
         );
  DLH_X1 \REGISTERS_reg[9][22]  ( .G(N3571), .D(N4130), .Q(\REGISTERS[9][22] )
         );
  DLH_X1 \REGISTERS_reg[9][21]  ( .G(N3571), .D(N4128), .Q(\REGISTERS[9][21] )
         );
  DLH_X1 \REGISTERS_reg[9][20]  ( .G(N3571), .D(N4126), .Q(\REGISTERS[9][20] )
         );
  DLH_X1 \REGISTERS_reg[9][19]  ( .G(N3571), .D(N4124), .Q(\REGISTERS[9][19] )
         );
  DLH_X1 \REGISTERS_reg[9][18]  ( .G(N3571), .D(N4122), .Q(\REGISTERS[9][18] )
         );
  DLH_X1 \REGISTERS_reg[9][17]  ( .G(N3571), .D(N4120), .Q(\REGISTERS[9][17] )
         );
  DLH_X1 \REGISTERS_reg[9][16]  ( .G(N3571), .D(N4118), .Q(\REGISTERS[9][16] )
         );
  DLH_X1 \REGISTERS_reg[9][15]  ( .G(N3571), .D(N4116), .Q(\REGISTERS[9][15] )
         );
  DLH_X1 \REGISTERS_reg[9][14]  ( .G(N3571), .D(N4114), .Q(\REGISTERS[9][14] )
         );
  DLH_X1 \REGISTERS_reg[9][13]  ( .G(N3571), .D(N4112), .Q(\REGISTERS[9][13] )
         );
  DLH_X1 \REGISTERS_reg[9][12]  ( .G(N3571), .D(N4110), .Q(\REGISTERS[9][12] )
         );
  DLH_X1 \REGISTERS_reg[9][11]  ( .G(N3571), .D(N4108), .Q(\REGISTERS[9][11] )
         );
  DLH_X1 \REGISTERS_reg[9][10]  ( .G(N3571), .D(N4106), .Q(\REGISTERS[9][10] )
         );
  DLH_X1 \REGISTERS_reg[9][9]  ( .G(N3571), .D(N4104), .Q(\REGISTERS[9][9] )
         );
  DLH_X1 \REGISTERS_reg[9][8]  ( .G(N3571), .D(N4102), .Q(\REGISTERS[9][8] )
         );
  DLH_X1 \REGISTERS_reg[9][7]  ( .G(N3571), .D(N4100), .Q(\REGISTERS[9][7] )
         );
  DLH_X1 \REGISTERS_reg[9][6]  ( .G(N3571), .D(N4098), .Q(\REGISTERS[9][6] )
         );
  DLH_X1 \REGISTERS_reg[9][5]  ( .G(N3571), .D(N4096), .Q(\REGISTERS[9][5] )
         );
  DLH_X1 \REGISTERS_reg[9][4]  ( .G(N3571), .D(N4094), .Q(\REGISTERS[9][4] )
         );
  DLH_X1 \REGISTERS_reg[9][3]  ( .G(N3571), .D(N4092), .Q(\REGISTERS[9][3] )
         );
  DLH_X1 \REGISTERS_reg[9][2]  ( .G(N3571), .D(N4090), .Q(\REGISTERS[9][2] )
         );
  DLH_X1 \REGISTERS_reg[9][1]  ( .G(N3571), .D(N4088), .Q(\REGISTERS[9][1] )
         );
  DLH_X1 \REGISTERS_reg[9][0]  ( .G(N3571), .D(N4086), .Q(\REGISTERS[9][0] )
         );
  DLH_X1 \REGISTERS_reg[10][31]  ( .G(N3507), .D(N4148), .Q(
        \REGISTERS[10][31] ) );
  DLH_X1 \REGISTERS_reg[10][30]  ( .G(N3507), .D(N4146), .Q(
        \REGISTERS[10][30] ) );
  DLH_X1 \REGISTERS_reg[10][29]  ( .G(N3507), .D(N4144), .Q(
        \REGISTERS[10][29] ) );
  DLH_X1 \REGISTERS_reg[10][28]  ( .G(N3507), .D(N4142), .Q(
        \REGISTERS[10][28] ) );
  DLH_X1 \REGISTERS_reg[10][27]  ( .G(N3507), .D(N4140), .Q(
        \REGISTERS[10][27] ) );
  DLH_X1 \REGISTERS_reg[10][26]  ( .G(N3507), .D(N4138), .Q(
        \REGISTERS[10][26] ) );
  DLH_X1 \REGISTERS_reg[10][25]  ( .G(N3507), .D(N4136), .Q(
        \REGISTERS[10][25] ) );
  DLH_X1 \REGISTERS_reg[10][24]  ( .G(N3507), .D(N4134), .Q(
        \REGISTERS[10][24] ) );
  DLH_X1 \REGISTERS_reg[10][23]  ( .G(N3507), .D(N4132), .Q(
        \REGISTERS[10][23] ) );
  DLH_X1 \REGISTERS_reg[10][22]  ( .G(N3507), .D(N4130), .Q(
        \REGISTERS[10][22] ) );
  DLH_X1 \REGISTERS_reg[10][21]  ( .G(N3507), .D(N4128), .Q(
        \REGISTERS[10][21] ) );
  DLH_X1 \REGISTERS_reg[10][20]  ( .G(N3507), .D(N4126), .Q(
        \REGISTERS[10][20] ) );
  DLH_X1 \REGISTERS_reg[10][19]  ( .G(N3507), .D(N4124), .Q(
        \REGISTERS[10][19] ) );
  DLH_X1 \REGISTERS_reg[10][18]  ( .G(N3507), .D(N4122), .Q(
        \REGISTERS[10][18] ) );
  DLH_X1 \REGISTERS_reg[10][17]  ( .G(N3507), .D(N4120), .Q(
        \REGISTERS[10][17] ) );
  DLH_X1 \REGISTERS_reg[10][16]  ( .G(N3507), .D(N4118), .Q(
        \REGISTERS[10][16] ) );
  DLH_X1 \REGISTERS_reg[10][15]  ( .G(N3507), .D(N4116), .Q(
        \REGISTERS[10][15] ) );
  DLH_X1 \REGISTERS_reg[10][14]  ( .G(N3507), .D(N4114), .Q(
        \REGISTERS[10][14] ) );
  DLH_X1 \REGISTERS_reg[10][13]  ( .G(N3507), .D(N4112), .Q(
        \REGISTERS[10][13] ) );
  DLH_X1 \REGISTERS_reg[10][12]  ( .G(N3507), .D(N4110), .Q(
        \REGISTERS[10][12] ) );
  DLH_X1 \REGISTERS_reg[10][11]  ( .G(N3507), .D(N4108), .Q(
        \REGISTERS[10][11] ) );
  DLH_X1 \REGISTERS_reg[10][10]  ( .G(N3507), .D(N4106), .Q(
        \REGISTERS[10][10] ) );
  DLH_X1 \REGISTERS_reg[10][9]  ( .G(N3507), .D(N4104), .Q(\REGISTERS[10][9] )
         );
  DLH_X1 \REGISTERS_reg[10][8]  ( .G(N3507), .D(N4102), .Q(\REGISTERS[10][8] )
         );
  DLH_X1 \REGISTERS_reg[10][7]  ( .G(N3507), .D(N4100), .Q(\REGISTERS[10][7] )
         );
  DLH_X1 \REGISTERS_reg[10][6]  ( .G(N3507), .D(N4098), .Q(\REGISTERS[10][6] )
         );
  DLH_X1 \REGISTERS_reg[10][5]  ( .G(N3507), .D(N4096), .Q(\REGISTERS[10][5] )
         );
  DLH_X1 \REGISTERS_reg[10][4]  ( .G(N3507), .D(N4094), .Q(\REGISTERS[10][4] )
         );
  DLH_X1 \REGISTERS_reg[10][3]  ( .G(N3507), .D(N4092), .Q(\REGISTERS[10][3] )
         );
  DLH_X1 \REGISTERS_reg[10][2]  ( .G(N3507), .D(N4090), .Q(\REGISTERS[10][2] )
         );
  DLH_X1 \REGISTERS_reg[10][1]  ( .G(N3507), .D(N4088), .Q(\REGISTERS[10][1] )
         );
  DLH_X1 \REGISTERS_reg[10][0]  ( .G(N3507), .D(N4086), .Q(\REGISTERS[10][0] )
         );
  DLH_X1 \REGISTERS_reg[11][31]  ( .G(N3443), .D(N4148), .Q(
        \REGISTERS[11][31] ) );
  DLH_X1 \REGISTERS_reg[11][30]  ( .G(N3443), .D(N4146), .Q(
        \REGISTERS[11][30] ) );
  DLH_X1 \REGISTERS_reg[11][29]  ( .G(N3443), .D(N4144), .Q(
        \REGISTERS[11][29] ) );
  DLH_X1 \REGISTERS_reg[11][28]  ( .G(N3443), .D(N4142), .Q(
        \REGISTERS[11][28] ) );
  DLH_X1 \REGISTERS_reg[11][27]  ( .G(N3443), .D(N4140), .Q(
        \REGISTERS[11][27] ) );
  DLH_X1 \REGISTERS_reg[11][26]  ( .G(N3443), .D(N4138), .Q(
        \REGISTERS[11][26] ) );
  DLH_X1 \REGISTERS_reg[11][25]  ( .G(N3443), .D(N4136), .Q(
        \REGISTERS[11][25] ) );
  DLH_X1 \REGISTERS_reg[11][24]  ( .G(N3443), .D(N4134), .Q(
        \REGISTERS[11][24] ) );
  DLH_X1 \REGISTERS_reg[11][23]  ( .G(N3443), .D(N4132), .Q(
        \REGISTERS[11][23] ) );
  DLH_X1 \REGISTERS_reg[11][22]  ( .G(N3443), .D(N4130), .Q(
        \REGISTERS[11][22] ) );
  DLH_X1 \REGISTERS_reg[11][21]  ( .G(N3443), .D(N4128), .Q(
        \REGISTERS[11][21] ) );
  DLH_X1 \REGISTERS_reg[11][20]  ( .G(N3443), .D(N4126), .Q(
        \REGISTERS[11][20] ) );
  DLH_X1 \REGISTERS_reg[11][19]  ( .G(N3443), .D(N4124), .Q(
        \REGISTERS[11][19] ) );
  DLH_X1 \REGISTERS_reg[11][18]  ( .G(N3443), .D(N4122), .Q(
        \REGISTERS[11][18] ) );
  DLH_X1 \REGISTERS_reg[11][17]  ( .G(N3443), .D(N4120), .Q(
        \REGISTERS[11][17] ) );
  DLH_X1 \REGISTERS_reg[11][16]  ( .G(N3443), .D(N4118), .Q(
        \REGISTERS[11][16] ) );
  DLH_X1 \REGISTERS_reg[11][15]  ( .G(N3443), .D(N4116), .Q(
        \REGISTERS[11][15] ) );
  DLH_X1 \REGISTERS_reg[11][14]  ( .G(N3443), .D(N4114), .Q(
        \REGISTERS[11][14] ) );
  DLH_X1 \REGISTERS_reg[11][13]  ( .G(N3443), .D(N4112), .Q(
        \REGISTERS[11][13] ) );
  DLH_X1 \REGISTERS_reg[11][12]  ( .G(N3443), .D(N4110), .Q(
        \REGISTERS[11][12] ) );
  DLH_X1 \REGISTERS_reg[11][11]  ( .G(N3443), .D(N4108), .Q(
        \REGISTERS[11][11] ) );
  DLH_X1 \REGISTERS_reg[11][10]  ( .G(N3443), .D(N4106), .Q(
        \REGISTERS[11][10] ) );
  DLH_X1 \REGISTERS_reg[11][9]  ( .G(N3443), .D(N4104), .Q(\REGISTERS[11][9] )
         );
  DLH_X1 \REGISTERS_reg[11][8]  ( .G(N3443), .D(N4102), .Q(\REGISTERS[11][8] )
         );
  DLH_X1 \REGISTERS_reg[11][7]  ( .G(N3443), .D(N4100), .Q(\REGISTERS[11][7] )
         );
  DLH_X1 \REGISTERS_reg[11][6]  ( .G(N3443), .D(N4098), .Q(\REGISTERS[11][6] )
         );
  DLH_X1 \REGISTERS_reg[11][5]  ( .G(N3443), .D(N4096), .Q(\REGISTERS[11][5] )
         );
  DLH_X1 \REGISTERS_reg[11][4]  ( .G(N3443), .D(N4094), .Q(\REGISTERS[11][4] )
         );
  DLH_X1 \REGISTERS_reg[11][3]  ( .G(N3443), .D(N4092), .Q(\REGISTERS[11][3] )
         );
  DLH_X1 \REGISTERS_reg[11][2]  ( .G(N3443), .D(N4090), .Q(\REGISTERS[11][2] )
         );
  DLH_X1 \REGISTERS_reg[11][1]  ( .G(N3443), .D(N4088), .Q(\REGISTERS[11][1] )
         );
  DLH_X1 \REGISTERS_reg[11][0]  ( .G(N3443), .D(N4086), .Q(\REGISTERS[11][0] )
         );
  DLH_X1 \REGISTERS_reg[12][31]  ( .G(N3379), .D(N4148), .Q(
        \REGISTERS[12][31] ) );
  DLH_X1 \REGISTERS_reg[12][30]  ( .G(N3379), .D(N4146), .Q(
        \REGISTERS[12][30] ) );
  DLH_X1 \REGISTERS_reg[12][29]  ( .G(N3379), .D(N4144), .Q(
        \REGISTERS[12][29] ) );
  DLH_X1 \REGISTERS_reg[12][28]  ( .G(N3379), .D(N4142), .Q(
        \REGISTERS[12][28] ) );
  DLH_X1 \REGISTERS_reg[12][27]  ( .G(N3379), .D(N4140), .Q(
        \REGISTERS[12][27] ) );
  DLH_X1 \REGISTERS_reg[12][26]  ( .G(N3379), .D(N4138), .Q(
        \REGISTERS[12][26] ) );
  DLH_X1 \REGISTERS_reg[12][25]  ( .G(N3379), .D(N4136), .Q(
        \REGISTERS[12][25] ) );
  DLH_X1 \REGISTERS_reg[12][24]  ( .G(N3379), .D(N4134), .Q(
        \REGISTERS[12][24] ) );
  DLH_X1 \REGISTERS_reg[12][23]  ( .G(N3379), .D(N4132), .Q(
        \REGISTERS[12][23] ) );
  DLH_X1 \REGISTERS_reg[12][22]  ( .G(N3379), .D(N4130), .Q(
        \REGISTERS[12][22] ) );
  DLH_X1 \REGISTERS_reg[12][21]  ( .G(N3379), .D(N4128), .Q(
        \REGISTERS[12][21] ) );
  DLH_X1 \REGISTERS_reg[12][20]  ( .G(N3379), .D(N4126), .Q(
        \REGISTERS[12][20] ) );
  DLH_X1 \REGISTERS_reg[12][19]  ( .G(N3379), .D(N4124), .Q(
        \REGISTERS[12][19] ) );
  DLH_X1 \REGISTERS_reg[12][18]  ( .G(N3379), .D(N4122), .Q(
        \REGISTERS[12][18] ) );
  DLH_X1 \REGISTERS_reg[12][17]  ( .G(N3379), .D(N4120), .Q(
        \REGISTERS[12][17] ) );
  DLH_X1 \REGISTERS_reg[12][16]  ( .G(N3379), .D(N4118), .Q(
        \REGISTERS[12][16] ) );
  DLH_X1 \REGISTERS_reg[12][15]  ( .G(N3379), .D(N4116), .Q(
        \REGISTERS[12][15] ) );
  DLH_X1 \REGISTERS_reg[12][14]  ( .G(N3379), .D(N4114), .Q(
        \REGISTERS[12][14] ) );
  DLH_X1 \REGISTERS_reg[12][13]  ( .G(N3379), .D(N4112), .Q(
        \REGISTERS[12][13] ) );
  DLH_X1 \REGISTERS_reg[12][12]  ( .G(N3379), .D(N4110), .Q(
        \REGISTERS[12][12] ) );
  DLH_X1 \REGISTERS_reg[12][11]  ( .G(N3379), .D(N4108), .Q(
        \REGISTERS[12][11] ) );
  DLH_X1 \REGISTERS_reg[12][10]  ( .G(N3379), .D(N4106), .Q(
        \REGISTERS[12][10] ) );
  DLH_X1 \REGISTERS_reg[12][9]  ( .G(N3379), .D(N4104), .Q(\REGISTERS[12][9] )
         );
  DLH_X1 \REGISTERS_reg[12][8]  ( .G(N3379), .D(N4102), .Q(\REGISTERS[12][8] )
         );
  DLH_X1 \REGISTERS_reg[12][7]  ( .G(N3379), .D(N4100), .Q(\REGISTERS[12][7] )
         );
  DLH_X1 \REGISTERS_reg[12][6]  ( .G(N3379), .D(N4098), .Q(\REGISTERS[12][6] )
         );
  DLH_X1 \REGISTERS_reg[12][5]  ( .G(N3379), .D(N4096), .Q(\REGISTERS[12][5] )
         );
  DLH_X1 \REGISTERS_reg[12][4]  ( .G(N3379), .D(N4094), .Q(\REGISTERS[12][4] )
         );
  DLH_X1 \REGISTERS_reg[12][3]  ( .G(N3379), .D(N4092), .Q(\REGISTERS[12][3] )
         );
  DLH_X1 \REGISTERS_reg[12][2]  ( .G(N3379), .D(N4090), .Q(\REGISTERS[12][2] )
         );
  DLH_X1 \REGISTERS_reg[12][1]  ( .G(N3379), .D(N4088), .Q(\REGISTERS[12][1] )
         );
  DLH_X1 \REGISTERS_reg[12][0]  ( .G(N3379), .D(N4086), .Q(\REGISTERS[12][0] )
         );
  DLH_X1 \REGISTERS_reg[13][31]  ( .G(N3315), .D(N4148), .Q(
        \REGISTERS[13][31] ) );
  DLH_X1 \REGISTERS_reg[13][30]  ( .G(N3315), .D(N4146), .Q(
        \REGISTERS[13][30] ) );
  DLH_X1 \REGISTERS_reg[13][29]  ( .G(N3315), .D(N4144), .Q(
        \REGISTERS[13][29] ) );
  DLH_X1 \REGISTERS_reg[13][28]  ( .G(N3315), .D(N4142), .Q(
        \REGISTERS[13][28] ) );
  DLH_X1 \REGISTERS_reg[13][27]  ( .G(N3315), .D(N4140), .Q(
        \REGISTERS[13][27] ) );
  DLH_X1 \REGISTERS_reg[13][26]  ( .G(N3315), .D(N4138), .Q(
        \REGISTERS[13][26] ) );
  DLH_X1 \REGISTERS_reg[13][25]  ( .G(N3315), .D(N4136), .Q(
        \REGISTERS[13][25] ) );
  DLH_X1 \REGISTERS_reg[13][24]  ( .G(N3315), .D(N4134), .Q(
        \REGISTERS[13][24] ) );
  DLH_X1 \REGISTERS_reg[13][23]  ( .G(N3315), .D(N4132), .Q(
        \REGISTERS[13][23] ) );
  DLH_X1 \REGISTERS_reg[13][22]  ( .G(N3315), .D(N4130), .Q(
        \REGISTERS[13][22] ) );
  DLH_X1 \REGISTERS_reg[13][21]  ( .G(N3315), .D(N4128), .Q(
        \REGISTERS[13][21] ) );
  DLH_X1 \REGISTERS_reg[13][20]  ( .G(N3315), .D(N4126), .Q(
        \REGISTERS[13][20] ) );
  DLH_X1 \REGISTERS_reg[13][19]  ( .G(N3315), .D(N4124), .Q(
        \REGISTERS[13][19] ) );
  DLH_X1 \REGISTERS_reg[13][18]  ( .G(N3315), .D(N4122), .Q(
        \REGISTERS[13][18] ) );
  DLH_X1 \REGISTERS_reg[13][17]  ( .G(N3315), .D(N4120), .Q(
        \REGISTERS[13][17] ) );
  DLH_X1 \REGISTERS_reg[13][16]  ( .G(N3315), .D(N4118), .Q(
        \REGISTERS[13][16] ) );
  DLH_X1 \REGISTERS_reg[13][15]  ( .G(N3315), .D(N4116), .Q(
        \REGISTERS[13][15] ) );
  DLH_X1 \REGISTERS_reg[13][14]  ( .G(N3315), .D(N4114), .Q(
        \REGISTERS[13][14] ) );
  DLH_X1 \REGISTERS_reg[13][13]  ( .G(N3315), .D(N4112), .Q(
        \REGISTERS[13][13] ) );
  DLH_X1 \REGISTERS_reg[13][12]  ( .G(N3315), .D(N4110), .Q(
        \REGISTERS[13][12] ) );
  DLH_X1 \REGISTERS_reg[13][11]  ( .G(N3315), .D(N4108), .Q(
        \REGISTERS[13][11] ) );
  DLH_X1 \REGISTERS_reg[13][10]  ( .G(N3315), .D(N4106), .Q(
        \REGISTERS[13][10] ) );
  DLH_X1 \REGISTERS_reg[13][9]  ( .G(N3315), .D(N4104), .Q(\REGISTERS[13][9] )
         );
  DLH_X1 \REGISTERS_reg[13][8]  ( .G(N3315), .D(N4102), .Q(\REGISTERS[13][8] )
         );
  DLH_X1 \REGISTERS_reg[13][7]  ( .G(N3315), .D(N4100), .Q(\REGISTERS[13][7] )
         );
  DLH_X1 \REGISTERS_reg[13][6]  ( .G(N3315), .D(N4098), .Q(\REGISTERS[13][6] )
         );
  DLH_X1 \REGISTERS_reg[13][5]  ( .G(N3315), .D(N4096), .Q(\REGISTERS[13][5] )
         );
  DLH_X1 \REGISTERS_reg[13][4]  ( .G(N3315), .D(N4094), .Q(\REGISTERS[13][4] )
         );
  DLH_X1 \REGISTERS_reg[13][3]  ( .G(N3315), .D(N4092), .Q(\REGISTERS[13][3] )
         );
  DLH_X1 \REGISTERS_reg[13][2]  ( .G(N3315), .D(N4090), .Q(\REGISTERS[13][2] )
         );
  DLH_X1 \REGISTERS_reg[13][1]  ( .G(N3315), .D(N4088), .Q(\REGISTERS[13][1] )
         );
  DLH_X1 \REGISTERS_reg[13][0]  ( .G(N3315), .D(N4086), .Q(\REGISTERS[13][0] )
         );
  DLH_X1 \REGISTERS_reg[14][31]  ( .G(N3251), .D(N4148), .Q(
        \REGISTERS[14][31] ) );
  DLH_X1 \REGISTERS_reg[14][30]  ( .G(N3251), .D(N4146), .Q(
        \REGISTERS[14][30] ) );
  DLH_X1 \REGISTERS_reg[14][29]  ( .G(N3251), .D(N4144), .Q(
        \REGISTERS[14][29] ) );
  DLH_X1 \REGISTERS_reg[14][28]  ( .G(N3251), .D(N4142), .Q(
        \REGISTERS[14][28] ) );
  DLH_X1 \REGISTERS_reg[14][27]  ( .G(N3251), .D(N4140), .Q(
        \REGISTERS[14][27] ) );
  DLH_X1 \REGISTERS_reg[14][26]  ( .G(N3251), .D(N4138), .Q(
        \REGISTERS[14][26] ) );
  DLH_X1 \REGISTERS_reg[14][25]  ( .G(N3251), .D(N4136), .Q(
        \REGISTERS[14][25] ) );
  DLH_X1 \REGISTERS_reg[14][24]  ( .G(N3251), .D(N4134), .Q(
        \REGISTERS[14][24] ) );
  DLH_X1 \REGISTERS_reg[14][23]  ( .G(N3251), .D(N4132), .Q(
        \REGISTERS[14][23] ) );
  DLH_X1 \REGISTERS_reg[14][22]  ( .G(N3251), .D(N4130), .Q(
        \REGISTERS[14][22] ) );
  DLH_X1 \REGISTERS_reg[14][21]  ( .G(N3251), .D(N4128), .Q(
        \REGISTERS[14][21] ) );
  DLH_X1 \REGISTERS_reg[14][20]  ( .G(N3251), .D(N4126), .Q(
        \REGISTERS[14][20] ) );
  DLH_X1 \REGISTERS_reg[14][19]  ( .G(N3251), .D(N4124), .Q(
        \REGISTERS[14][19] ) );
  DLH_X1 \REGISTERS_reg[14][18]  ( .G(N3251), .D(N4122), .Q(
        \REGISTERS[14][18] ) );
  DLH_X1 \REGISTERS_reg[14][17]  ( .G(N3251), .D(N4120), .Q(
        \REGISTERS[14][17] ) );
  DLH_X1 \REGISTERS_reg[14][16]  ( .G(N3251), .D(N4118), .Q(
        \REGISTERS[14][16] ) );
  DLH_X1 \REGISTERS_reg[14][15]  ( .G(N3251), .D(N4116), .Q(
        \REGISTERS[14][15] ) );
  DLH_X1 \REGISTERS_reg[14][14]  ( .G(N3251), .D(N4114), .Q(
        \REGISTERS[14][14] ) );
  DLH_X1 \REGISTERS_reg[14][13]  ( .G(N3251), .D(N4112), .Q(
        \REGISTERS[14][13] ) );
  DLH_X1 \REGISTERS_reg[14][12]  ( .G(N3251), .D(N4110), .Q(
        \REGISTERS[14][12] ) );
  DLH_X1 \REGISTERS_reg[14][11]  ( .G(N3251), .D(N4108), .Q(
        \REGISTERS[14][11] ) );
  DLH_X1 \REGISTERS_reg[14][10]  ( .G(N3251), .D(N4106), .Q(
        \REGISTERS[14][10] ) );
  DLH_X1 \REGISTERS_reg[14][9]  ( .G(N3251), .D(N4104), .Q(\REGISTERS[14][9] )
         );
  DLH_X1 \REGISTERS_reg[14][8]  ( .G(N3251), .D(N4102), .Q(\REGISTERS[14][8] )
         );
  DLH_X1 \REGISTERS_reg[14][7]  ( .G(N3251), .D(N4100), .Q(\REGISTERS[14][7] )
         );
  DLH_X1 \REGISTERS_reg[14][6]  ( .G(N3251), .D(N4098), .Q(\REGISTERS[14][6] )
         );
  DLH_X1 \REGISTERS_reg[14][5]  ( .G(N3251), .D(N4096), .Q(\REGISTERS[14][5] )
         );
  DLH_X1 \REGISTERS_reg[14][4]  ( .G(N3251), .D(N4094), .Q(\REGISTERS[14][4] )
         );
  DLH_X1 \REGISTERS_reg[14][3]  ( .G(N3251), .D(N4092), .Q(\REGISTERS[14][3] )
         );
  DLH_X1 \REGISTERS_reg[14][2]  ( .G(N3251), .D(N4090), .Q(\REGISTERS[14][2] )
         );
  DLH_X1 \REGISTERS_reg[14][1]  ( .G(N3251), .D(N4088), .Q(\REGISTERS[14][1] )
         );
  DLH_X1 \REGISTERS_reg[14][0]  ( .G(N3251), .D(N4086), .Q(\REGISTERS[14][0] )
         );
  DLH_X1 \REGISTERS_reg[15][31]  ( .G(N3187), .D(N4148), .Q(
        \REGISTERS[15][31] ) );
  DLH_X1 \REGISTERS_reg[15][30]  ( .G(N3187), .D(N4146), .Q(
        \REGISTERS[15][30] ) );
  DLH_X1 \REGISTERS_reg[15][29]  ( .G(N3187), .D(N4144), .Q(
        \REGISTERS[15][29] ) );
  DLH_X1 \REGISTERS_reg[15][28]  ( .G(N3187), .D(N4142), .Q(
        \REGISTERS[15][28] ) );
  DLH_X1 \REGISTERS_reg[15][27]  ( .G(N3187), .D(N4140), .Q(
        \REGISTERS[15][27] ) );
  DLH_X1 \REGISTERS_reg[15][26]  ( .G(N3187), .D(N4138), .Q(
        \REGISTERS[15][26] ) );
  DLH_X1 \REGISTERS_reg[15][25]  ( .G(N3187), .D(N4136), .Q(
        \REGISTERS[15][25] ) );
  DLH_X1 \REGISTERS_reg[15][24]  ( .G(N3187), .D(N4134), .Q(
        \REGISTERS[15][24] ) );
  DLH_X1 \REGISTERS_reg[15][23]  ( .G(N3187), .D(N4132), .Q(
        \REGISTERS[15][23] ) );
  DLH_X1 \REGISTERS_reg[15][22]  ( .G(N3187), .D(N4130), .Q(
        \REGISTERS[15][22] ) );
  DLH_X1 \REGISTERS_reg[15][21]  ( .G(N3187), .D(N4128), .Q(
        \REGISTERS[15][21] ) );
  DLH_X1 \REGISTERS_reg[15][20]  ( .G(N3187), .D(N4126), .Q(
        \REGISTERS[15][20] ) );
  DLH_X1 \REGISTERS_reg[15][19]  ( .G(N3187), .D(N4124), .Q(
        \REGISTERS[15][19] ) );
  DLH_X1 \REGISTERS_reg[15][18]  ( .G(N3187), .D(N4122), .Q(
        \REGISTERS[15][18] ) );
  DLH_X1 \REGISTERS_reg[15][17]  ( .G(N3187), .D(N4120), .Q(
        \REGISTERS[15][17] ) );
  DLH_X1 \REGISTERS_reg[15][16]  ( .G(N3187), .D(N4118), .Q(
        \REGISTERS[15][16] ) );
  DLH_X1 \REGISTERS_reg[15][15]  ( .G(N3187), .D(N4116), .Q(
        \REGISTERS[15][15] ) );
  DLH_X1 \REGISTERS_reg[15][14]  ( .G(N3187), .D(N4114), .Q(
        \REGISTERS[15][14] ) );
  DLH_X1 \REGISTERS_reg[15][13]  ( .G(N3187), .D(N4112), .Q(
        \REGISTERS[15][13] ) );
  DLH_X1 \REGISTERS_reg[15][12]  ( .G(N3187), .D(N4110), .Q(
        \REGISTERS[15][12] ) );
  DLH_X1 \REGISTERS_reg[15][11]  ( .G(N3187), .D(N4108), .Q(
        \REGISTERS[15][11] ) );
  DLH_X1 \REGISTERS_reg[15][10]  ( .G(N3187), .D(N4106), .Q(
        \REGISTERS[15][10] ) );
  DLH_X1 \REGISTERS_reg[15][9]  ( .G(N3187), .D(N4104), .Q(\REGISTERS[15][9] )
         );
  DLH_X1 \REGISTERS_reg[15][8]  ( .G(N3187), .D(N4102), .Q(\REGISTERS[15][8] )
         );
  DLH_X1 \REGISTERS_reg[15][7]  ( .G(N3187), .D(N4100), .Q(\REGISTERS[15][7] )
         );
  DLH_X1 \REGISTERS_reg[15][6]  ( .G(N3187), .D(N4098), .Q(\REGISTERS[15][6] )
         );
  DLH_X1 \REGISTERS_reg[15][5]  ( .G(N3187), .D(N4096), .Q(\REGISTERS[15][5] )
         );
  DLH_X1 \REGISTERS_reg[15][4]  ( .G(N3187), .D(N4094), .Q(\REGISTERS[15][4] )
         );
  DLH_X1 \REGISTERS_reg[15][3]  ( .G(N3187), .D(N4092), .Q(\REGISTERS[15][3] )
         );
  DLH_X1 \REGISTERS_reg[15][2]  ( .G(N3187), .D(N4090), .Q(\REGISTERS[15][2] )
         );
  DLH_X1 \REGISTERS_reg[15][1]  ( .G(N3187), .D(N4088), .Q(\REGISTERS[15][1] )
         );
  DLH_X1 \REGISTERS_reg[15][0]  ( .G(N3187), .D(N4086), .Q(\REGISTERS[15][0] )
         );
  DLH_X1 \REGISTERS_reg[16][31]  ( .G(N3123), .D(N4148), .Q(
        \REGISTERS[16][31] ) );
  DLH_X1 \REGISTERS_reg[16][30]  ( .G(N3123), .D(N4146), .Q(
        \REGISTERS[16][30] ) );
  DLH_X1 \REGISTERS_reg[16][29]  ( .G(N3123), .D(N4144), .Q(
        \REGISTERS[16][29] ) );
  DLH_X1 \REGISTERS_reg[16][28]  ( .G(N3123), .D(N4142), .Q(
        \REGISTERS[16][28] ) );
  DLH_X1 \REGISTERS_reg[16][27]  ( .G(N3123), .D(N4140), .Q(
        \REGISTERS[16][27] ) );
  DLH_X1 \REGISTERS_reg[16][26]  ( .G(N3123), .D(N4138), .Q(
        \REGISTERS[16][26] ) );
  DLH_X1 \REGISTERS_reg[16][25]  ( .G(N3123), .D(N4136), .Q(
        \REGISTERS[16][25] ) );
  DLH_X1 \REGISTERS_reg[16][24]  ( .G(N3123), .D(N4134), .Q(
        \REGISTERS[16][24] ) );
  DLH_X1 \REGISTERS_reg[16][23]  ( .G(N3123), .D(N4132), .Q(
        \REGISTERS[16][23] ) );
  DLH_X1 \REGISTERS_reg[16][22]  ( .G(N3123), .D(N4130), .Q(
        \REGISTERS[16][22] ) );
  DLH_X1 \REGISTERS_reg[16][21]  ( .G(N3123), .D(N4128), .Q(
        \REGISTERS[16][21] ) );
  DLH_X1 \REGISTERS_reg[16][20]  ( .G(N3123), .D(N4126), .Q(
        \REGISTERS[16][20] ) );
  DLH_X1 \REGISTERS_reg[16][19]  ( .G(N3123), .D(N4124), .Q(
        \REGISTERS[16][19] ) );
  DLH_X1 \REGISTERS_reg[16][18]  ( .G(N3123), .D(N4122), .Q(
        \REGISTERS[16][18] ) );
  DLH_X1 \REGISTERS_reg[16][17]  ( .G(N3123), .D(N4120), .Q(
        \REGISTERS[16][17] ) );
  DLH_X1 \REGISTERS_reg[16][16]  ( .G(N3123), .D(N4118), .Q(
        \REGISTERS[16][16] ) );
  DLH_X1 \REGISTERS_reg[16][15]  ( .G(N3123), .D(N4116), .Q(
        \REGISTERS[16][15] ) );
  DLH_X1 \REGISTERS_reg[16][14]  ( .G(N3123), .D(N4114), .Q(
        \REGISTERS[16][14] ) );
  DLH_X1 \REGISTERS_reg[16][13]  ( .G(N3123), .D(N4112), .Q(
        \REGISTERS[16][13] ) );
  DLH_X1 \REGISTERS_reg[16][12]  ( .G(N3123), .D(N4110), .Q(
        \REGISTERS[16][12] ) );
  DLH_X1 \REGISTERS_reg[16][11]  ( .G(N3123), .D(N4108), .Q(
        \REGISTERS[16][11] ) );
  DLH_X1 \REGISTERS_reg[16][10]  ( .G(N3123), .D(N4106), .Q(
        \REGISTERS[16][10] ) );
  DLH_X1 \REGISTERS_reg[16][9]  ( .G(N3123), .D(N4104), .Q(\REGISTERS[16][9] )
         );
  DLH_X1 \REGISTERS_reg[16][8]  ( .G(N3123), .D(N4102), .Q(\REGISTERS[16][8] )
         );
  DLH_X1 \REGISTERS_reg[16][7]  ( .G(N3123), .D(N4100), .Q(\REGISTERS[16][7] )
         );
  DLH_X1 \REGISTERS_reg[16][6]  ( .G(N3123), .D(N4098), .Q(\REGISTERS[16][6] )
         );
  DLH_X1 \REGISTERS_reg[16][5]  ( .G(N3123), .D(N4096), .Q(\REGISTERS[16][5] )
         );
  DLH_X1 \REGISTERS_reg[16][4]  ( .G(N3123), .D(N4094), .Q(\REGISTERS[16][4] )
         );
  DLH_X1 \REGISTERS_reg[16][3]  ( .G(N3123), .D(N4092), .Q(\REGISTERS[16][3] )
         );
  DLH_X1 \REGISTERS_reg[16][2]  ( .G(N3123), .D(N4090), .Q(\REGISTERS[16][2] )
         );
  DLH_X1 \REGISTERS_reg[16][1]  ( .G(N3123), .D(N4088), .Q(\REGISTERS[16][1] )
         );
  DLH_X1 \REGISTERS_reg[16][0]  ( .G(N3123), .D(N4086), .Q(\REGISTERS[16][0] )
         );
  DLH_X1 \REGISTERS_reg[17][31]  ( .G(N3059), .D(N4148), .Q(
        \REGISTERS[17][31] ) );
  DLH_X1 \REGISTERS_reg[17][30]  ( .G(N3059), .D(N4146), .Q(
        \REGISTERS[17][30] ) );
  DLH_X1 \REGISTERS_reg[17][29]  ( .G(N3059), .D(N4144), .Q(
        \REGISTERS[17][29] ) );
  DLH_X1 \REGISTERS_reg[17][28]  ( .G(N3059), .D(N4142), .Q(
        \REGISTERS[17][28] ) );
  DLH_X1 \REGISTERS_reg[17][27]  ( .G(N3059), .D(N4140), .Q(
        \REGISTERS[17][27] ) );
  DLH_X1 \REGISTERS_reg[17][26]  ( .G(N3059), .D(N4138), .Q(
        \REGISTERS[17][26] ) );
  DLH_X1 \REGISTERS_reg[17][25]  ( .G(N3059), .D(N4136), .Q(
        \REGISTERS[17][25] ) );
  DLH_X1 \REGISTERS_reg[17][24]  ( .G(N3059), .D(N4134), .Q(
        \REGISTERS[17][24] ) );
  DLH_X1 \REGISTERS_reg[17][23]  ( .G(N3059), .D(N4132), .Q(
        \REGISTERS[17][23] ) );
  DLH_X1 \REGISTERS_reg[17][22]  ( .G(N3059), .D(N4130), .Q(
        \REGISTERS[17][22] ) );
  DLH_X1 \REGISTERS_reg[17][21]  ( .G(N3059), .D(N4128), .Q(
        \REGISTERS[17][21] ) );
  DLH_X1 \REGISTERS_reg[17][20]  ( .G(N3059), .D(N4126), .Q(
        \REGISTERS[17][20] ) );
  DLH_X1 \REGISTERS_reg[17][19]  ( .G(N3059), .D(N4124), .Q(
        \REGISTERS[17][19] ) );
  DLH_X1 \REGISTERS_reg[17][18]  ( .G(N3059), .D(N4122), .Q(
        \REGISTERS[17][18] ) );
  DLH_X1 \REGISTERS_reg[17][17]  ( .G(N3059), .D(N4120), .Q(
        \REGISTERS[17][17] ) );
  DLH_X1 \REGISTERS_reg[17][16]  ( .G(N3059), .D(N4118), .Q(
        \REGISTERS[17][16] ) );
  DLH_X1 \REGISTERS_reg[17][15]  ( .G(N3059), .D(N4116), .Q(
        \REGISTERS[17][15] ) );
  DLH_X1 \REGISTERS_reg[17][14]  ( .G(N3059), .D(N4114), .Q(
        \REGISTERS[17][14] ) );
  DLH_X1 \REGISTERS_reg[17][13]  ( .G(N3059), .D(N4112), .Q(
        \REGISTERS[17][13] ) );
  DLH_X1 \REGISTERS_reg[17][12]  ( .G(N3059), .D(N4110), .Q(
        \REGISTERS[17][12] ) );
  DLH_X1 \REGISTERS_reg[17][11]  ( .G(N3059), .D(N4108), .Q(
        \REGISTERS[17][11] ) );
  DLH_X1 \REGISTERS_reg[17][10]  ( .G(N3059), .D(N4106), .Q(
        \REGISTERS[17][10] ) );
  DLH_X1 \REGISTERS_reg[17][9]  ( .G(N3059), .D(N4104), .Q(\REGISTERS[17][9] )
         );
  DLH_X1 \REGISTERS_reg[17][8]  ( .G(N3059), .D(N4102), .Q(\REGISTERS[17][8] )
         );
  DLH_X1 \REGISTERS_reg[17][7]  ( .G(N3059), .D(N4100), .Q(\REGISTERS[17][7] )
         );
  DLH_X1 \REGISTERS_reg[17][6]  ( .G(N3059), .D(N4098), .Q(\REGISTERS[17][6] )
         );
  DLH_X1 \REGISTERS_reg[17][5]  ( .G(N3059), .D(N4096), .Q(\REGISTERS[17][5] )
         );
  DLH_X1 \REGISTERS_reg[17][4]  ( .G(N3059), .D(N4094), .Q(\REGISTERS[17][4] )
         );
  DLH_X1 \REGISTERS_reg[17][3]  ( .G(N3059), .D(N4092), .Q(\REGISTERS[17][3] )
         );
  DLH_X1 \REGISTERS_reg[17][2]  ( .G(N3059), .D(N4090), .Q(\REGISTERS[17][2] )
         );
  DLH_X1 \REGISTERS_reg[17][1]  ( .G(N3059), .D(N4088), .Q(\REGISTERS[17][1] )
         );
  DLH_X1 \REGISTERS_reg[17][0]  ( .G(N3059), .D(N4086), .Q(\REGISTERS[17][0] )
         );
  DLH_X1 \REGISTERS_reg[18][31]  ( .G(N2995), .D(N4148), .Q(
        \REGISTERS[18][31] ) );
  DLH_X1 \REGISTERS_reg[18][30]  ( .G(N2995), .D(N4146), .Q(
        \REGISTERS[18][30] ) );
  DLH_X1 \REGISTERS_reg[18][29]  ( .G(N2995), .D(N4144), .Q(
        \REGISTERS[18][29] ) );
  DLH_X1 \REGISTERS_reg[18][28]  ( .G(N2995), .D(N4142), .Q(
        \REGISTERS[18][28] ) );
  DLH_X1 \REGISTERS_reg[18][27]  ( .G(N2995), .D(N4140), .Q(
        \REGISTERS[18][27] ) );
  DLH_X1 \REGISTERS_reg[18][26]  ( .G(N2995), .D(N4138), .Q(
        \REGISTERS[18][26] ) );
  DLH_X1 \REGISTERS_reg[18][25]  ( .G(N2995), .D(N4136), .Q(
        \REGISTERS[18][25] ) );
  DLH_X1 \REGISTERS_reg[18][24]  ( .G(N2995), .D(N4134), .Q(
        \REGISTERS[18][24] ) );
  DLH_X1 \REGISTERS_reg[18][23]  ( .G(N2995), .D(N4132), .Q(
        \REGISTERS[18][23] ) );
  DLH_X1 \REGISTERS_reg[18][22]  ( .G(N2995), .D(N4130), .Q(
        \REGISTERS[18][22] ) );
  DLH_X1 \REGISTERS_reg[18][21]  ( .G(N2995), .D(N4128), .Q(
        \REGISTERS[18][21] ) );
  DLH_X1 \REGISTERS_reg[18][20]  ( .G(N2995), .D(N4126), .Q(
        \REGISTERS[18][20] ) );
  DLH_X1 \REGISTERS_reg[18][19]  ( .G(N2995), .D(N4124), .Q(
        \REGISTERS[18][19] ) );
  DLH_X1 \REGISTERS_reg[18][18]  ( .G(N2995), .D(N4122), .Q(
        \REGISTERS[18][18] ) );
  DLH_X1 \REGISTERS_reg[18][17]  ( .G(N2995), .D(N4120), .Q(
        \REGISTERS[18][17] ) );
  DLH_X1 \REGISTERS_reg[18][16]  ( .G(N2995), .D(N4118), .Q(
        \REGISTERS[18][16] ) );
  DLH_X1 \REGISTERS_reg[18][15]  ( .G(N2995), .D(N4116), .Q(
        \REGISTERS[18][15] ) );
  DLH_X1 \REGISTERS_reg[18][14]  ( .G(N2995), .D(N4114), .Q(
        \REGISTERS[18][14] ) );
  DLH_X1 \REGISTERS_reg[18][13]  ( .G(N2995), .D(N4112), .Q(
        \REGISTERS[18][13] ) );
  DLH_X1 \REGISTERS_reg[18][12]  ( .G(N2995), .D(N4110), .Q(
        \REGISTERS[18][12] ) );
  DLH_X1 \REGISTERS_reg[18][11]  ( .G(N2995), .D(N4108), .Q(
        \REGISTERS[18][11] ) );
  DLH_X1 \REGISTERS_reg[18][10]  ( .G(N2995), .D(N4106), .Q(
        \REGISTERS[18][10] ) );
  DLH_X1 \REGISTERS_reg[18][9]  ( .G(N2995), .D(N4104), .Q(\REGISTERS[18][9] )
         );
  DLH_X1 \REGISTERS_reg[18][8]  ( .G(N2995), .D(N4102), .Q(\REGISTERS[18][8] )
         );
  DLH_X1 \REGISTERS_reg[18][7]  ( .G(N2995), .D(N4100), .Q(\REGISTERS[18][7] )
         );
  DLH_X1 \REGISTERS_reg[18][6]  ( .G(N2995), .D(N4098), .Q(\REGISTERS[18][6] )
         );
  DLH_X1 \REGISTERS_reg[18][5]  ( .G(N2995), .D(N4096), .Q(\REGISTERS[18][5] )
         );
  DLH_X1 \REGISTERS_reg[18][4]  ( .G(N2995), .D(N4094), .Q(\REGISTERS[18][4] )
         );
  DLH_X1 \REGISTERS_reg[18][3]  ( .G(N2995), .D(N4092), .Q(\REGISTERS[18][3] )
         );
  DLH_X1 \REGISTERS_reg[18][2]  ( .G(N2995), .D(N4090), .Q(\REGISTERS[18][2] )
         );
  DLH_X1 \REGISTERS_reg[18][1]  ( .G(N2995), .D(N4088), .Q(\REGISTERS[18][1] )
         );
  DLH_X1 \REGISTERS_reg[18][0]  ( .G(N2995), .D(N4086), .Q(\REGISTERS[18][0] )
         );
  DLH_X1 \REGISTERS_reg[19][31]  ( .G(N2931), .D(N4148), .Q(
        \REGISTERS[19][31] ) );
  DLH_X1 \REGISTERS_reg[19][30]  ( .G(N2931), .D(N4146), .Q(
        \REGISTERS[19][30] ) );
  DLH_X1 \REGISTERS_reg[19][29]  ( .G(N2931), .D(N4144), .Q(
        \REGISTERS[19][29] ) );
  DLH_X1 \REGISTERS_reg[19][28]  ( .G(N2931), .D(N4142), .Q(
        \REGISTERS[19][28] ) );
  DLH_X1 \REGISTERS_reg[19][27]  ( .G(N2931), .D(N4140), .Q(
        \REGISTERS[19][27] ) );
  DLH_X1 \REGISTERS_reg[19][26]  ( .G(N2931), .D(N4138), .Q(
        \REGISTERS[19][26] ) );
  DLH_X1 \REGISTERS_reg[19][25]  ( .G(N2931), .D(N4136), .Q(
        \REGISTERS[19][25] ) );
  DLH_X1 \REGISTERS_reg[19][24]  ( .G(N2931), .D(N4134), .Q(
        \REGISTERS[19][24] ) );
  DLH_X1 \REGISTERS_reg[19][23]  ( .G(N2931), .D(N4132), .Q(
        \REGISTERS[19][23] ) );
  DLH_X1 \REGISTERS_reg[19][22]  ( .G(N2931), .D(N4130), .Q(
        \REGISTERS[19][22] ) );
  DLH_X1 \REGISTERS_reg[19][21]  ( .G(N2931), .D(N4128), .Q(
        \REGISTERS[19][21] ) );
  DLH_X1 \REGISTERS_reg[19][20]  ( .G(N2931), .D(N4126), .Q(
        \REGISTERS[19][20] ) );
  DLH_X1 \REGISTERS_reg[19][19]  ( .G(N2931), .D(N4124), .Q(
        \REGISTERS[19][19] ) );
  DLH_X1 \REGISTERS_reg[19][18]  ( .G(N2931), .D(N4122), .Q(
        \REGISTERS[19][18] ) );
  DLH_X1 \REGISTERS_reg[19][17]  ( .G(N2931), .D(N4120), .Q(
        \REGISTERS[19][17] ) );
  DLH_X1 \REGISTERS_reg[19][16]  ( .G(N2931), .D(N4118), .Q(
        \REGISTERS[19][16] ) );
  DLH_X1 \REGISTERS_reg[19][15]  ( .G(N2931), .D(N4116), .Q(
        \REGISTERS[19][15] ) );
  DLH_X1 \REGISTERS_reg[19][14]  ( .G(N2931), .D(N4114), .Q(
        \REGISTERS[19][14] ) );
  DLH_X1 \REGISTERS_reg[19][13]  ( .G(N2931), .D(N4112), .Q(
        \REGISTERS[19][13] ) );
  DLH_X1 \REGISTERS_reg[19][12]  ( .G(N2931), .D(N4110), .Q(
        \REGISTERS[19][12] ) );
  DLH_X1 \REGISTERS_reg[19][11]  ( .G(N2931), .D(N4108), .Q(
        \REGISTERS[19][11] ) );
  DLH_X1 \REGISTERS_reg[19][10]  ( .G(N2931), .D(N4106), .Q(
        \REGISTERS[19][10] ) );
  DLH_X1 \REGISTERS_reg[19][9]  ( .G(N2931), .D(N4104), .Q(\REGISTERS[19][9] )
         );
  DLH_X1 \REGISTERS_reg[19][8]  ( .G(N2931), .D(N4102), .Q(\REGISTERS[19][8] )
         );
  DLH_X1 \REGISTERS_reg[19][7]  ( .G(N2931), .D(N4100), .Q(\REGISTERS[19][7] )
         );
  DLH_X1 \REGISTERS_reg[19][6]  ( .G(N2931), .D(N4098), .Q(\REGISTERS[19][6] )
         );
  DLH_X1 \REGISTERS_reg[19][5]  ( .G(N2931), .D(N4096), .Q(\REGISTERS[19][5] )
         );
  DLH_X1 \REGISTERS_reg[19][4]  ( .G(N2931), .D(N4094), .Q(\REGISTERS[19][4] )
         );
  DLH_X1 \REGISTERS_reg[19][3]  ( .G(N2931), .D(N4092), .Q(\REGISTERS[19][3] )
         );
  DLH_X1 \REGISTERS_reg[19][2]  ( .G(N2931), .D(N4090), .Q(\REGISTERS[19][2] )
         );
  DLH_X1 \REGISTERS_reg[19][1]  ( .G(N2931), .D(N4088), .Q(\REGISTERS[19][1] )
         );
  DLH_X1 \REGISTERS_reg[19][0]  ( .G(N2931), .D(N4086), .Q(\REGISTERS[19][0] )
         );
  DLH_X1 \REGISTERS_reg[20][31]  ( .G(N2867), .D(N4148), .Q(
        \REGISTERS[20][31] ) );
  DLH_X1 \REGISTERS_reg[20][30]  ( .G(N2867), .D(N4146), .Q(
        \REGISTERS[20][30] ) );
  DLH_X1 \REGISTERS_reg[20][29]  ( .G(N2867), .D(N4144), .Q(
        \REGISTERS[20][29] ) );
  DLH_X1 \REGISTERS_reg[20][28]  ( .G(N2867), .D(N4142), .Q(
        \REGISTERS[20][28] ) );
  DLH_X1 \REGISTERS_reg[20][27]  ( .G(N2867), .D(N4140), .Q(
        \REGISTERS[20][27] ) );
  DLH_X1 \REGISTERS_reg[20][26]  ( .G(N2867), .D(N4138), .Q(
        \REGISTERS[20][26] ) );
  DLH_X1 \REGISTERS_reg[20][25]  ( .G(N2867), .D(N4136), .Q(
        \REGISTERS[20][25] ) );
  DLH_X1 \REGISTERS_reg[20][24]  ( .G(N2867), .D(N4134), .Q(
        \REGISTERS[20][24] ) );
  DLH_X1 \REGISTERS_reg[20][23]  ( .G(N2867), .D(N4132), .Q(
        \REGISTERS[20][23] ) );
  DLH_X1 \REGISTERS_reg[20][22]  ( .G(N2867), .D(N4130), .Q(
        \REGISTERS[20][22] ) );
  DLH_X1 \REGISTERS_reg[20][21]  ( .G(N2867), .D(N4128), .Q(
        \REGISTERS[20][21] ) );
  DLH_X1 \REGISTERS_reg[20][20]  ( .G(N2867), .D(N4126), .Q(
        \REGISTERS[20][20] ) );
  DLH_X1 \REGISTERS_reg[20][19]  ( .G(N2867), .D(N4124), .Q(
        \REGISTERS[20][19] ) );
  DLH_X1 \REGISTERS_reg[20][18]  ( .G(N2867), .D(N4122), .Q(
        \REGISTERS[20][18] ) );
  DLH_X1 \REGISTERS_reg[20][17]  ( .G(N2867), .D(N4120), .Q(
        \REGISTERS[20][17] ) );
  DLH_X1 \REGISTERS_reg[20][16]  ( .G(N2867), .D(N4118), .Q(
        \REGISTERS[20][16] ) );
  DLH_X1 \REGISTERS_reg[20][15]  ( .G(N2867), .D(N4116), .Q(
        \REGISTERS[20][15] ) );
  DLH_X1 \REGISTERS_reg[20][14]  ( .G(N2867), .D(N4114), .Q(
        \REGISTERS[20][14] ) );
  DLH_X1 \REGISTERS_reg[20][13]  ( .G(N2867), .D(N4112), .Q(
        \REGISTERS[20][13] ) );
  DLH_X1 \REGISTERS_reg[20][12]  ( .G(N2867), .D(N4110), .Q(
        \REGISTERS[20][12] ) );
  DLH_X1 \REGISTERS_reg[20][11]  ( .G(N2867), .D(N4108), .Q(
        \REGISTERS[20][11] ) );
  DLH_X1 \REGISTERS_reg[20][10]  ( .G(N2867), .D(N4106), .Q(
        \REGISTERS[20][10] ) );
  DLH_X1 \REGISTERS_reg[20][9]  ( .G(N2867), .D(N4104), .Q(\REGISTERS[20][9] )
         );
  DLH_X1 \REGISTERS_reg[20][8]  ( .G(N2867), .D(N4102), .Q(\REGISTERS[20][8] )
         );
  DLH_X1 \REGISTERS_reg[20][7]  ( .G(N2867), .D(N4100), .Q(\REGISTERS[20][7] )
         );
  DLH_X1 \REGISTERS_reg[20][6]  ( .G(N2867), .D(N4098), .Q(\REGISTERS[20][6] )
         );
  DLH_X1 \REGISTERS_reg[20][5]  ( .G(N2867), .D(N4096), .Q(\REGISTERS[20][5] )
         );
  DLH_X1 \REGISTERS_reg[20][4]  ( .G(N2867), .D(N4094), .Q(\REGISTERS[20][4] )
         );
  DLH_X1 \REGISTERS_reg[20][3]  ( .G(N2867), .D(N4092), .Q(\REGISTERS[20][3] )
         );
  DLH_X1 \REGISTERS_reg[20][2]  ( .G(N2867), .D(N4090), .Q(\REGISTERS[20][2] )
         );
  DLH_X1 \REGISTERS_reg[20][1]  ( .G(N2867), .D(N4088), .Q(\REGISTERS[20][1] )
         );
  DLH_X1 \REGISTERS_reg[20][0]  ( .G(N2867), .D(N4086), .Q(\REGISTERS[20][0] )
         );
  DLH_X1 \REGISTERS_reg[21][31]  ( .G(N2803), .D(N4148), .Q(
        \REGISTERS[21][31] ) );
  DLH_X1 \REGISTERS_reg[21][30]  ( .G(N2803), .D(N4146), .Q(
        \REGISTERS[21][30] ) );
  DLH_X1 \REGISTERS_reg[21][29]  ( .G(N2803), .D(N4144), .Q(
        \REGISTERS[21][29] ) );
  DLH_X1 \REGISTERS_reg[21][28]  ( .G(N2803), .D(N4142), .Q(
        \REGISTERS[21][28] ) );
  DLH_X1 \REGISTERS_reg[21][27]  ( .G(N2803), .D(N4140), .Q(
        \REGISTERS[21][27] ) );
  DLH_X1 \REGISTERS_reg[21][26]  ( .G(N2803), .D(N4138), .Q(
        \REGISTERS[21][26] ) );
  DLH_X1 \REGISTERS_reg[21][25]  ( .G(N2803), .D(N4136), .Q(
        \REGISTERS[21][25] ) );
  DLH_X1 \REGISTERS_reg[21][24]  ( .G(N2803), .D(N4134), .Q(
        \REGISTERS[21][24] ) );
  DLH_X1 \REGISTERS_reg[21][23]  ( .G(N2803), .D(N4132), .Q(
        \REGISTERS[21][23] ) );
  DLH_X1 \REGISTERS_reg[21][22]  ( .G(N2803), .D(N4130), .Q(
        \REGISTERS[21][22] ) );
  DLH_X1 \REGISTERS_reg[21][21]  ( .G(N2803), .D(N4128), .Q(
        \REGISTERS[21][21] ) );
  DLH_X1 \REGISTERS_reg[21][20]  ( .G(N2803), .D(N4126), .Q(
        \REGISTERS[21][20] ) );
  DLH_X1 \REGISTERS_reg[21][19]  ( .G(N2803), .D(N4124), .Q(
        \REGISTERS[21][19] ) );
  DLH_X1 \REGISTERS_reg[21][18]  ( .G(N2803), .D(N4122), .Q(
        \REGISTERS[21][18] ) );
  DLH_X1 \REGISTERS_reg[21][17]  ( .G(N2803), .D(N4120), .Q(
        \REGISTERS[21][17] ) );
  DLH_X1 \REGISTERS_reg[21][16]  ( .G(N2803), .D(N4118), .Q(
        \REGISTERS[21][16] ) );
  DLH_X1 \REGISTERS_reg[21][15]  ( .G(N2803), .D(N4116), .Q(
        \REGISTERS[21][15] ) );
  DLH_X1 \REGISTERS_reg[21][14]  ( .G(N2803), .D(N4114), .Q(
        \REGISTERS[21][14] ) );
  DLH_X1 \REGISTERS_reg[21][13]  ( .G(N2803), .D(N4112), .Q(
        \REGISTERS[21][13] ) );
  DLH_X1 \REGISTERS_reg[21][12]  ( .G(N2803), .D(N4110), .Q(
        \REGISTERS[21][12] ) );
  DLH_X1 \REGISTERS_reg[21][11]  ( .G(N2803), .D(N4108), .Q(
        \REGISTERS[21][11] ) );
  DLH_X1 \REGISTERS_reg[21][10]  ( .G(N2803), .D(N4106), .Q(
        \REGISTERS[21][10] ) );
  DLH_X1 \REGISTERS_reg[21][9]  ( .G(N2803), .D(N4104), .Q(\REGISTERS[21][9] )
         );
  DLH_X1 \REGISTERS_reg[21][8]  ( .G(N2803), .D(N4102), .Q(\REGISTERS[21][8] )
         );
  DLH_X1 \REGISTERS_reg[21][7]  ( .G(N2803), .D(N4100), .Q(\REGISTERS[21][7] )
         );
  DLH_X1 \REGISTERS_reg[21][6]  ( .G(N2803), .D(N4098), .Q(\REGISTERS[21][6] )
         );
  DLH_X1 \REGISTERS_reg[21][5]  ( .G(N2803), .D(N4096), .Q(\REGISTERS[21][5] )
         );
  DLH_X1 \REGISTERS_reg[21][4]  ( .G(N2803), .D(N4094), .Q(\REGISTERS[21][4] )
         );
  DLH_X1 \REGISTERS_reg[21][3]  ( .G(N2803), .D(N4092), .Q(\REGISTERS[21][3] )
         );
  DLH_X1 \REGISTERS_reg[21][2]  ( .G(N2803), .D(N4090), .Q(\REGISTERS[21][2] )
         );
  DLH_X1 \REGISTERS_reg[21][1]  ( .G(N2803), .D(N4088), .Q(\REGISTERS[21][1] )
         );
  DLH_X1 \REGISTERS_reg[21][0]  ( .G(N2803), .D(N4086), .Q(\REGISTERS[21][0] )
         );
  DLH_X1 \REGISTERS_reg[22][31]  ( .G(N2739), .D(N4148), .Q(
        \REGISTERS[22][31] ) );
  DLH_X1 \REGISTERS_reg[22][30]  ( .G(N2739), .D(N4146), .Q(
        \REGISTERS[22][30] ) );
  DLH_X1 \REGISTERS_reg[22][29]  ( .G(N2739), .D(N4144), .Q(
        \REGISTERS[22][29] ) );
  DLH_X1 \REGISTERS_reg[22][28]  ( .G(N2739), .D(N4142), .Q(
        \REGISTERS[22][28] ) );
  DLH_X1 \REGISTERS_reg[22][27]  ( .G(N2739), .D(N4140), .Q(
        \REGISTERS[22][27] ) );
  DLH_X1 \REGISTERS_reg[22][26]  ( .G(N2739), .D(N4138), .Q(
        \REGISTERS[22][26] ) );
  DLH_X1 \REGISTERS_reg[22][25]  ( .G(N2739), .D(N4136), .Q(
        \REGISTERS[22][25] ) );
  DLH_X1 \REGISTERS_reg[22][24]  ( .G(N2739), .D(N4134), .Q(
        \REGISTERS[22][24] ) );
  DLH_X1 \REGISTERS_reg[22][23]  ( .G(N2739), .D(N4132), .Q(
        \REGISTERS[22][23] ) );
  DLH_X1 \REGISTERS_reg[22][22]  ( .G(N2739), .D(N4130), .Q(
        \REGISTERS[22][22] ) );
  DLH_X1 \REGISTERS_reg[22][21]  ( .G(N2739), .D(N4128), .Q(
        \REGISTERS[22][21] ) );
  DLH_X1 \REGISTERS_reg[22][20]  ( .G(N2739), .D(N4126), .Q(
        \REGISTERS[22][20] ) );
  DLH_X1 \REGISTERS_reg[22][19]  ( .G(N2739), .D(N4124), .Q(
        \REGISTERS[22][19] ) );
  DLH_X1 \REGISTERS_reg[22][18]  ( .G(N2739), .D(N4122), .Q(
        \REGISTERS[22][18] ) );
  DLH_X1 \REGISTERS_reg[22][17]  ( .G(N2739), .D(N4120), .Q(
        \REGISTERS[22][17] ) );
  DLH_X1 \REGISTERS_reg[22][16]  ( .G(N2739), .D(N4118), .Q(
        \REGISTERS[22][16] ) );
  DLH_X1 \REGISTERS_reg[22][15]  ( .G(N2739), .D(N4116), .Q(
        \REGISTERS[22][15] ) );
  DLH_X1 \REGISTERS_reg[22][14]  ( .G(N2739), .D(N4114), .Q(
        \REGISTERS[22][14] ) );
  DLH_X1 \REGISTERS_reg[22][13]  ( .G(N2739), .D(N4112), .Q(
        \REGISTERS[22][13] ) );
  DLH_X1 \REGISTERS_reg[22][12]  ( .G(N2739), .D(N4110), .Q(
        \REGISTERS[22][12] ) );
  DLH_X1 \REGISTERS_reg[22][11]  ( .G(N2739), .D(N4108), .Q(
        \REGISTERS[22][11] ) );
  DLH_X1 \REGISTERS_reg[22][10]  ( .G(N2739), .D(N4106), .Q(
        \REGISTERS[22][10] ) );
  DLH_X1 \REGISTERS_reg[22][9]  ( .G(N2739), .D(N4104), .Q(\REGISTERS[22][9] )
         );
  DLH_X1 \REGISTERS_reg[22][8]  ( .G(N2739), .D(N4102), .Q(\REGISTERS[22][8] )
         );
  DLH_X1 \REGISTERS_reg[22][7]  ( .G(N2739), .D(N4100), .Q(\REGISTERS[22][7] )
         );
  DLH_X1 \REGISTERS_reg[22][6]  ( .G(N2739), .D(N4098), .Q(\REGISTERS[22][6] )
         );
  DLH_X1 \REGISTERS_reg[22][5]  ( .G(N2739), .D(N4096), .Q(\REGISTERS[22][5] )
         );
  DLH_X1 \REGISTERS_reg[22][4]  ( .G(N2739), .D(N4094), .Q(\REGISTERS[22][4] )
         );
  DLH_X1 \REGISTERS_reg[22][3]  ( .G(N2739), .D(N4092), .Q(\REGISTERS[22][3] )
         );
  DLH_X1 \REGISTERS_reg[22][2]  ( .G(N2739), .D(N4090), .Q(\REGISTERS[22][2] )
         );
  DLH_X1 \REGISTERS_reg[22][1]  ( .G(N2739), .D(N4088), .Q(\REGISTERS[22][1] )
         );
  DLH_X1 \REGISTERS_reg[22][0]  ( .G(N2739), .D(N4086), .Q(\REGISTERS[22][0] )
         );
  DLH_X1 \REGISTERS_reg[23][31]  ( .G(N2675), .D(N4148), .Q(
        \REGISTERS[23][31] ) );
  DLH_X1 \REGISTERS_reg[23][30]  ( .G(N2675), .D(N4146), .Q(
        \REGISTERS[23][30] ) );
  DLH_X1 \REGISTERS_reg[23][29]  ( .G(N2675), .D(N4144), .Q(
        \REGISTERS[23][29] ) );
  DLH_X1 \REGISTERS_reg[23][28]  ( .G(N2675), .D(N4142), .Q(
        \REGISTERS[23][28] ) );
  DLH_X1 \REGISTERS_reg[23][27]  ( .G(N2675), .D(N4140), .Q(
        \REGISTERS[23][27] ) );
  DLH_X1 \REGISTERS_reg[23][26]  ( .G(N2675), .D(N4138), .Q(
        \REGISTERS[23][26] ) );
  DLH_X1 \REGISTERS_reg[23][25]  ( .G(N2675), .D(N4136), .Q(
        \REGISTERS[23][25] ) );
  DLH_X1 \REGISTERS_reg[23][24]  ( .G(N2675), .D(N4134), .Q(
        \REGISTERS[23][24] ) );
  DLH_X1 \REGISTERS_reg[23][23]  ( .G(N2675), .D(N4132), .Q(
        \REGISTERS[23][23] ) );
  DLH_X1 \REGISTERS_reg[23][22]  ( .G(N2675), .D(N4130), .Q(
        \REGISTERS[23][22] ) );
  DLH_X1 \REGISTERS_reg[23][21]  ( .G(N2675), .D(N4128), .Q(
        \REGISTERS[23][21] ) );
  DLH_X1 \REGISTERS_reg[23][20]  ( .G(N2675), .D(N4126), .Q(
        \REGISTERS[23][20] ) );
  DLH_X1 \REGISTERS_reg[23][19]  ( .G(N2675), .D(N4124), .Q(
        \REGISTERS[23][19] ) );
  DLH_X1 \REGISTERS_reg[23][18]  ( .G(N2675), .D(N4122), .Q(
        \REGISTERS[23][18] ) );
  DLH_X1 \REGISTERS_reg[23][17]  ( .G(N2675), .D(N4120), .Q(
        \REGISTERS[23][17] ) );
  DLH_X1 \REGISTERS_reg[23][16]  ( .G(N2675), .D(N4118), .Q(
        \REGISTERS[23][16] ) );
  DLH_X1 \REGISTERS_reg[23][15]  ( .G(N2675), .D(N4116), .Q(
        \REGISTERS[23][15] ) );
  DLH_X1 \REGISTERS_reg[23][14]  ( .G(N2675), .D(N4114), .Q(
        \REGISTERS[23][14] ) );
  DLH_X1 \REGISTERS_reg[23][13]  ( .G(N2675), .D(N4112), .Q(
        \REGISTERS[23][13] ) );
  DLH_X1 \REGISTERS_reg[23][12]  ( .G(N2675), .D(N4110), .Q(
        \REGISTERS[23][12] ) );
  DLH_X1 \REGISTERS_reg[23][11]  ( .G(N2675), .D(N4108), .Q(
        \REGISTERS[23][11] ) );
  DLH_X1 \REGISTERS_reg[23][10]  ( .G(N2675), .D(N4106), .Q(
        \REGISTERS[23][10] ) );
  DLH_X1 \REGISTERS_reg[23][9]  ( .G(N2675), .D(N4104), .Q(\REGISTERS[23][9] )
         );
  DLH_X1 \REGISTERS_reg[23][8]  ( .G(N2675), .D(N4102), .Q(\REGISTERS[23][8] )
         );
  DLH_X1 \REGISTERS_reg[23][7]  ( .G(N2675), .D(N4100), .Q(\REGISTERS[23][7] )
         );
  DLH_X1 \REGISTERS_reg[23][6]  ( .G(N2675), .D(N4098), .Q(\REGISTERS[23][6] )
         );
  DLH_X1 \REGISTERS_reg[23][5]  ( .G(N2675), .D(N4096), .Q(\REGISTERS[23][5] )
         );
  DLH_X1 \REGISTERS_reg[23][4]  ( .G(N2675), .D(N4094), .Q(\REGISTERS[23][4] )
         );
  DLH_X1 \REGISTERS_reg[23][3]  ( .G(N2675), .D(N4092), .Q(\REGISTERS[23][3] )
         );
  DLH_X1 \REGISTERS_reg[23][2]  ( .G(N2675), .D(N4090), .Q(\REGISTERS[23][2] )
         );
  DLH_X1 \REGISTERS_reg[23][1]  ( .G(N2675), .D(N4088), .Q(\REGISTERS[23][1] )
         );
  DLH_X1 \REGISTERS_reg[23][0]  ( .G(N2675), .D(N4086), .Q(\REGISTERS[23][0] )
         );
  DLH_X1 \REGISTERS_reg[24][31]  ( .G(N2611), .D(N4148), .Q(
        \REGISTERS[24][31] ) );
  DLH_X1 \REGISTERS_reg[24][30]  ( .G(N2611), .D(N4146), .Q(
        \REGISTERS[24][30] ) );
  DLH_X1 \REGISTERS_reg[24][29]  ( .G(N2611), .D(N4144), .Q(
        \REGISTERS[24][29] ) );
  DLH_X1 \REGISTERS_reg[24][28]  ( .G(N2611), .D(N4142), .Q(
        \REGISTERS[24][28] ) );
  DLH_X1 \REGISTERS_reg[24][27]  ( .G(N2611), .D(N4140), .Q(
        \REGISTERS[24][27] ) );
  DLH_X1 \REGISTERS_reg[24][26]  ( .G(N2611), .D(N4138), .Q(
        \REGISTERS[24][26] ) );
  DLH_X1 \REGISTERS_reg[24][25]  ( .G(N2611), .D(N4136), .Q(
        \REGISTERS[24][25] ) );
  DLH_X1 \REGISTERS_reg[24][24]  ( .G(N2611), .D(N4134), .Q(
        \REGISTERS[24][24] ) );
  DLH_X1 \REGISTERS_reg[24][23]  ( .G(N2611), .D(N4132), .Q(
        \REGISTERS[24][23] ) );
  DLH_X1 \REGISTERS_reg[24][22]  ( .G(N2611), .D(N4130), .Q(
        \REGISTERS[24][22] ) );
  DLH_X1 \REGISTERS_reg[24][21]  ( .G(N2611), .D(N4128), .Q(
        \REGISTERS[24][21] ) );
  DLH_X1 \REGISTERS_reg[24][20]  ( .G(N2611), .D(N4126), .Q(
        \REGISTERS[24][20] ) );
  DLH_X1 \REGISTERS_reg[24][19]  ( .G(N2611), .D(N4124), .Q(
        \REGISTERS[24][19] ) );
  DLH_X1 \REGISTERS_reg[24][18]  ( .G(N2611), .D(N4122), .Q(
        \REGISTERS[24][18] ) );
  DLH_X1 \REGISTERS_reg[24][17]  ( .G(N2611), .D(N4120), .Q(
        \REGISTERS[24][17] ) );
  DLH_X1 \REGISTERS_reg[24][16]  ( .G(N2611), .D(N4118), .Q(
        \REGISTERS[24][16] ) );
  DLH_X1 \REGISTERS_reg[24][15]  ( .G(N2611), .D(N4116), .Q(
        \REGISTERS[24][15] ) );
  DLH_X1 \REGISTERS_reg[24][14]  ( .G(N2611), .D(N4114), .Q(
        \REGISTERS[24][14] ) );
  DLH_X1 \REGISTERS_reg[24][13]  ( .G(N2611), .D(N4112), .Q(
        \REGISTERS[24][13] ) );
  DLH_X1 \REGISTERS_reg[24][12]  ( .G(N2611), .D(N4110), .Q(
        \REGISTERS[24][12] ) );
  DLH_X1 \REGISTERS_reg[24][11]  ( .G(N2611), .D(N4108), .Q(
        \REGISTERS[24][11] ) );
  DLH_X1 \REGISTERS_reg[24][10]  ( .G(N2611), .D(N4106), .Q(
        \REGISTERS[24][10] ) );
  DLH_X1 \REGISTERS_reg[24][9]  ( .G(N2611), .D(N4104), .Q(\REGISTERS[24][9] )
         );
  DLH_X1 \REGISTERS_reg[24][8]  ( .G(N2611), .D(N4102), .Q(\REGISTERS[24][8] )
         );
  DLH_X1 \REGISTERS_reg[24][7]  ( .G(N2611), .D(N4100), .Q(\REGISTERS[24][7] )
         );
  DLH_X1 \REGISTERS_reg[24][6]  ( .G(N2611), .D(N4098), .Q(\REGISTERS[24][6] )
         );
  DLH_X1 \REGISTERS_reg[24][5]  ( .G(N2611), .D(N4096), .Q(\REGISTERS[24][5] )
         );
  DLH_X1 \REGISTERS_reg[24][4]  ( .G(N2611), .D(N4094), .Q(\REGISTERS[24][4] )
         );
  DLH_X1 \REGISTERS_reg[24][3]  ( .G(N2611), .D(N4092), .Q(\REGISTERS[24][3] )
         );
  DLH_X1 \REGISTERS_reg[24][2]  ( .G(N2611), .D(N4090), .Q(\REGISTERS[24][2] )
         );
  DLH_X1 \REGISTERS_reg[24][1]  ( .G(N2611), .D(N4088), .Q(\REGISTERS[24][1] )
         );
  DLH_X1 \REGISTERS_reg[24][0]  ( .G(N2611), .D(N4086), .Q(\REGISTERS[24][0] )
         );
  DLH_X1 \REGISTERS_reg[25][31]  ( .G(N2547), .D(N4148), .Q(
        \REGISTERS[25][31] ) );
  DLH_X1 \REGISTERS_reg[25][30]  ( .G(N2547), .D(N4146), .Q(
        \REGISTERS[25][30] ) );
  DLH_X1 \REGISTERS_reg[25][29]  ( .G(N2547), .D(N4144), .Q(
        \REGISTERS[25][29] ) );
  DLH_X1 \REGISTERS_reg[25][28]  ( .G(N2547), .D(N4142), .Q(
        \REGISTERS[25][28] ) );
  DLH_X1 \REGISTERS_reg[25][27]  ( .G(N2547), .D(N4140), .Q(
        \REGISTERS[25][27] ) );
  DLH_X1 \REGISTERS_reg[25][26]  ( .G(N2547), .D(N4138), .Q(
        \REGISTERS[25][26] ) );
  DLH_X1 \REGISTERS_reg[25][25]  ( .G(N2547), .D(N4136), .Q(
        \REGISTERS[25][25] ) );
  DLH_X1 \REGISTERS_reg[25][24]  ( .G(N2547), .D(N4134), .Q(
        \REGISTERS[25][24] ) );
  DLH_X1 \REGISTERS_reg[25][23]  ( .G(N2547), .D(N4132), .Q(
        \REGISTERS[25][23] ) );
  DLH_X1 \REGISTERS_reg[25][22]  ( .G(N2547), .D(N4130), .Q(
        \REGISTERS[25][22] ) );
  DLH_X1 \REGISTERS_reg[25][21]  ( .G(N2547), .D(N4128), .Q(
        \REGISTERS[25][21] ) );
  DLH_X1 \REGISTERS_reg[25][20]  ( .G(N2547), .D(N4126), .Q(
        \REGISTERS[25][20] ) );
  DLH_X1 \REGISTERS_reg[25][19]  ( .G(N2547), .D(N4124), .Q(
        \REGISTERS[25][19] ) );
  DLH_X1 \REGISTERS_reg[25][18]  ( .G(N2547), .D(N4122), .Q(
        \REGISTERS[25][18] ) );
  DLH_X1 \REGISTERS_reg[25][17]  ( .G(N2547), .D(N4120), .Q(
        \REGISTERS[25][17] ) );
  DLH_X1 \REGISTERS_reg[25][16]  ( .G(N2547), .D(N4118), .Q(
        \REGISTERS[25][16] ) );
  DLH_X1 \REGISTERS_reg[25][15]  ( .G(N2547), .D(N4116), .Q(
        \REGISTERS[25][15] ) );
  DLH_X1 \REGISTERS_reg[25][14]  ( .G(N2547), .D(N4114), .Q(
        \REGISTERS[25][14] ) );
  DLH_X1 \REGISTERS_reg[25][13]  ( .G(N2547), .D(N4112), .Q(
        \REGISTERS[25][13] ) );
  DLH_X1 \REGISTERS_reg[25][12]  ( .G(N2547), .D(N4110), .Q(
        \REGISTERS[25][12] ) );
  DLH_X1 \REGISTERS_reg[25][11]  ( .G(N2547), .D(N4108), .Q(
        \REGISTERS[25][11] ) );
  DLH_X1 \REGISTERS_reg[25][10]  ( .G(N2547), .D(N4106), .Q(
        \REGISTERS[25][10] ) );
  DLH_X1 \REGISTERS_reg[25][9]  ( .G(N2547), .D(N4104), .Q(\REGISTERS[25][9] )
         );
  DLH_X1 \REGISTERS_reg[25][8]  ( .G(N2547), .D(N4102), .Q(\REGISTERS[25][8] )
         );
  DLH_X1 \REGISTERS_reg[25][7]  ( .G(N2547), .D(N4100), .Q(\REGISTERS[25][7] )
         );
  DLH_X1 \REGISTERS_reg[25][6]  ( .G(N2547), .D(N4098), .Q(\REGISTERS[25][6] )
         );
  DLH_X1 \REGISTERS_reg[25][5]  ( .G(N2547), .D(N4096), .Q(\REGISTERS[25][5] )
         );
  DLH_X1 \REGISTERS_reg[25][4]  ( .G(N2547), .D(N4094), .Q(\REGISTERS[25][4] )
         );
  DLH_X1 \REGISTERS_reg[25][3]  ( .G(N2547), .D(N4092), .Q(\REGISTERS[25][3] )
         );
  DLH_X1 \REGISTERS_reg[25][2]  ( .G(N2547), .D(N4090), .Q(\REGISTERS[25][2] )
         );
  DLH_X1 \REGISTERS_reg[25][1]  ( .G(N2547), .D(N4088), .Q(\REGISTERS[25][1] )
         );
  DLH_X1 \REGISTERS_reg[25][0]  ( .G(N2547), .D(N4086), .Q(\REGISTERS[25][0] )
         );
  DLH_X1 \REGISTERS_reg[26][31]  ( .G(N2483), .D(N4148), .Q(
        \REGISTERS[26][31] ) );
  DLH_X1 \REGISTERS_reg[26][30]  ( .G(N2483), .D(N4146), .Q(
        \REGISTERS[26][30] ) );
  DLH_X1 \REGISTERS_reg[26][29]  ( .G(N2483), .D(N4144), .Q(
        \REGISTERS[26][29] ) );
  DLH_X1 \REGISTERS_reg[26][28]  ( .G(N2483), .D(N4142), .Q(
        \REGISTERS[26][28] ) );
  DLH_X1 \REGISTERS_reg[26][27]  ( .G(N2483), .D(N4140), .Q(
        \REGISTERS[26][27] ) );
  DLH_X1 \REGISTERS_reg[26][26]  ( .G(N2483), .D(N4138), .Q(
        \REGISTERS[26][26] ) );
  DLH_X1 \REGISTERS_reg[26][25]  ( .G(N2483), .D(N4136), .Q(
        \REGISTERS[26][25] ) );
  DLH_X1 \REGISTERS_reg[26][24]  ( .G(N2483), .D(N4134), .Q(
        \REGISTERS[26][24] ) );
  DLH_X1 \REGISTERS_reg[26][23]  ( .G(N2483), .D(N4132), .Q(
        \REGISTERS[26][23] ) );
  DLH_X1 \REGISTERS_reg[26][22]  ( .G(N2483), .D(N4130), .Q(
        \REGISTERS[26][22] ) );
  DLH_X1 \REGISTERS_reg[26][21]  ( .G(N2483), .D(N4128), .Q(
        \REGISTERS[26][21] ) );
  DLH_X1 \REGISTERS_reg[26][20]  ( .G(N2483), .D(N4126), .Q(
        \REGISTERS[26][20] ) );
  DLH_X1 \REGISTERS_reg[26][19]  ( .G(N2483), .D(N4124), .Q(
        \REGISTERS[26][19] ) );
  DLH_X1 \REGISTERS_reg[26][18]  ( .G(N2483), .D(N4122), .Q(
        \REGISTERS[26][18] ) );
  DLH_X1 \REGISTERS_reg[26][17]  ( .G(N2483), .D(N4120), .Q(
        \REGISTERS[26][17] ) );
  DLH_X1 \REGISTERS_reg[26][16]  ( .G(N2483), .D(N4118), .Q(
        \REGISTERS[26][16] ) );
  DLH_X1 \REGISTERS_reg[26][15]  ( .G(N2483), .D(N4116), .Q(
        \REGISTERS[26][15] ) );
  DLH_X1 \REGISTERS_reg[26][14]  ( .G(N2483), .D(N4114), .Q(
        \REGISTERS[26][14] ) );
  DLH_X1 \REGISTERS_reg[26][13]  ( .G(N2483), .D(N4112), .Q(
        \REGISTERS[26][13] ) );
  DLH_X1 \REGISTERS_reg[26][12]  ( .G(N2483), .D(N4110), .Q(
        \REGISTERS[26][12] ) );
  DLH_X1 \REGISTERS_reg[26][11]  ( .G(N2483), .D(N4108), .Q(
        \REGISTERS[26][11] ) );
  DLH_X1 \REGISTERS_reg[26][10]  ( .G(N2483), .D(N4106), .Q(
        \REGISTERS[26][10] ) );
  DLH_X1 \REGISTERS_reg[26][9]  ( .G(N2483), .D(N4104), .Q(\REGISTERS[26][9] )
         );
  DLH_X1 \REGISTERS_reg[26][8]  ( .G(N2483), .D(N4102), .Q(\REGISTERS[26][8] )
         );
  DLH_X1 \REGISTERS_reg[26][7]  ( .G(N2483), .D(N4100), .Q(\REGISTERS[26][7] )
         );
  DLH_X1 \REGISTERS_reg[26][6]  ( .G(N2483), .D(N4098), .Q(\REGISTERS[26][6] )
         );
  DLH_X1 \REGISTERS_reg[26][5]  ( .G(N2483), .D(N4096), .Q(\REGISTERS[26][5] )
         );
  DLH_X1 \REGISTERS_reg[26][4]  ( .G(N2483), .D(N4094), .Q(\REGISTERS[26][4] )
         );
  DLH_X1 \REGISTERS_reg[26][3]  ( .G(N2483), .D(N4092), .Q(\REGISTERS[26][3] )
         );
  DLH_X1 \REGISTERS_reg[26][2]  ( .G(N2483), .D(N4090), .Q(\REGISTERS[26][2] )
         );
  DLH_X1 \REGISTERS_reg[26][1]  ( .G(N2483), .D(N4088), .Q(\REGISTERS[26][1] )
         );
  DLH_X1 \REGISTERS_reg[26][0]  ( .G(N2483), .D(N4086), .Q(\REGISTERS[26][0] )
         );
  DLH_X1 \REGISTERS_reg[27][31]  ( .G(N2419), .D(N4148), .Q(
        \REGISTERS[27][31] ) );
  DLH_X1 \REGISTERS_reg[27][30]  ( .G(N2419), .D(N4146), .Q(
        \REGISTERS[27][30] ) );
  DLH_X1 \REGISTERS_reg[27][29]  ( .G(N2419), .D(N4144), .Q(
        \REGISTERS[27][29] ) );
  DLH_X1 \REGISTERS_reg[27][28]  ( .G(N2419), .D(N4142), .Q(
        \REGISTERS[27][28] ) );
  DLH_X1 \REGISTERS_reg[27][27]  ( .G(N2419), .D(N4140), .Q(
        \REGISTERS[27][27] ) );
  DLH_X1 \REGISTERS_reg[27][26]  ( .G(N2419), .D(N4138), .Q(
        \REGISTERS[27][26] ) );
  DLH_X1 \REGISTERS_reg[27][25]  ( .G(N2419), .D(N4136), .Q(
        \REGISTERS[27][25] ) );
  DLH_X1 \REGISTERS_reg[27][24]  ( .G(N2419), .D(N4134), .Q(
        \REGISTERS[27][24] ) );
  DLH_X1 \REGISTERS_reg[27][23]  ( .G(N2419), .D(N4132), .Q(
        \REGISTERS[27][23] ) );
  DLH_X1 \REGISTERS_reg[27][22]  ( .G(N2419), .D(N4130), .Q(
        \REGISTERS[27][22] ) );
  DLH_X1 \REGISTERS_reg[27][21]  ( .G(N2419), .D(N4128), .Q(
        \REGISTERS[27][21] ) );
  DLH_X1 \REGISTERS_reg[27][20]  ( .G(N2419), .D(N4126), .Q(
        \REGISTERS[27][20] ) );
  DLH_X1 \REGISTERS_reg[27][19]  ( .G(N2419), .D(N4124), .Q(
        \REGISTERS[27][19] ) );
  DLH_X1 \REGISTERS_reg[27][18]  ( .G(N2419), .D(N4122), .Q(
        \REGISTERS[27][18] ) );
  DLH_X1 \REGISTERS_reg[27][17]  ( .G(N2419), .D(N4120), .Q(
        \REGISTERS[27][17] ) );
  DLH_X1 \REGISTERS_reg[27][16]  ( .G(N2419), .D(N4118), .Q(
        \REGISTERS[27][16] ) );
  DLH_X1 \REGISTERS_reg[27][15]  ( .G(N2419), .D(N4116), .Q(
        \REGISTERS[27][15] ) );
  DLH_X1 \REGISTERS_reg[27][14]  ( .G(N2419), .D(N4114), .Q(
        \REGISTERS[27][14] ) );
  DLH_X1 \REGISTERS_reg[27][13]  ( .G(N2419), .D(N4112), .Q(
        \REGISTERS[27][13] ) );
  DLH_X1 \REGISTERS_reg[27][12]  ( .G(N2419), .D(N4110), .Q(
        \REGISTERS[27][12] ) );
  DLH_X1 \REGISTERS_reg[27][11]  ( .G(N2419), .D(N4108), .Q(
        \REGISTERS[27][11] ) );
  DLH_X1 \REGISTERS_reg[27][10]  ( .G(N2419), .D(N4106), .Q(
        \REGISTERS[27][10] ) );
  DLH_X1 \REGISTERS_reg[27][9]  ( .G(N2419), .D(N4104), .Q(\REGISTERS[27][9] )
         );
  DLH_X1 \REGISTERS_reg[27][8]  ( .G(N2419), .D(N4102), .Q(\REGISTERS[27][8] )
         );
  DLH_X1 \REGISTERS_reg[27][7]  ( .G(N2419), .D(N4100), .Q(\REGISTERS[27][7] )
         );
  DLH_X1 \REGISTERS_reg[27][6]  ( .G(N2419), .D(N4098), .Q(\REGISTERS[27][6] )
         );
  DLH_X1 \REGISTERS_reg[27][5]  ( .G(N2419), .D(N4096), .Q(\REGISTERS[27][5] )
         );
  DLH_X1 \REGISTERS_reg[27][4]  ( .G(N2419), .D(N4094), .Q(\REGISTERS[27][4] )
         );
  DLH_X1 \REGISTERS_reg[27][3]  ( .G(N2419), .D(N4092), .Q(\REGISTERS[27][3] )
         );
  DLH_X1 \REGISTERS_reg[27][2]  ( .G(N2419), .D(N4090), .Q(\REGISTERS[27][2] )
         );
  DLH_X1 \REGISTERS_reg[27][1]  ( .G(N2419), .D(N4088), .Q(\REGISTERS[27][1] )
         );
  DLH_X1 \REGISTERS_reg[27][0]  ( .G(N2419), .D(N4086), .Q(\REGISTERS[27][0] )
         );
  DLH_X1 \REGISTERS_reg[28][31]  ( .G(N2355), .D(N4148), .Q(
        \REGISTERS[28][31] ) );
  DLH_X1 \REGISTERS_reg[28][30]  ( .G(N2355), .D(N4146), .Q(
        \REGISTERS[28][30] ) );
  DLH_X1 \REGISTERS_reg[28][29]  ( .G(N2355), .D(N4144), .Q(
        \REGISTERS[28][29] ) );
  DLH_X1 \REGISTERS_reg[28][28]  ( .G(N2355), .D(N4142), .Q(
        \REGISTERS[28][28] ) );
  DLH_X1 \REGISTERS_reg[28][27]  ( .G(N2355), .D(N4140), .Q(
        \REGISTERS[28][27] ) );
  DLH_X1 \REGISTERS_reg[28][26]  ( .G(N2355), .D(N4138), .Q(
        \REGISTERS[28][26] ) );
  DLH_X1 \REGISTERS_reg[28][25]  ( .G(N2355), .D(N4136), .Q(
        \REGISTERS[28][25] ) );
  DLH_X1 \REGISTERS_reg[28][24]  ( .G(N2355), .D(N4134), .Q(
        \REGISTERS[28][24] ) );
  DLH_X1 \REGISTERS_reg[28][23]  ( .G(N2355), .D(N4132), .Q(
        \REGISTERS[28][23] ) );
  DLH_X1 \REGISTERS_reg[28][22]  ( .G(N2355), .D(N4130), .Q(
        \REGISTERS[28][22] ) );
  DLH_X1 \REGISTERS_reg[28][21]  ( .G(N2355), .D(N4128), .Q(
        \REGISTERS[28][21] ) );
  DLH_X1 \REGISTERS_reg[28][20]  ( .G(N2355), .D(N4126), .Q(
        \REGISTERS[28][20] ) );
  DLH_X1 \REGISTERS_reg[28][19]  ( .G(N2355), .D(N4124), .Q(
        \REGISTERS[28][19] ) );
  DLH_X1 \REGISTERS_reg[28][18]  ( .G(N2355), .D(N4122), .Q(
        \REGISTERS[28][18] ) );
  DLH_X1 \REGISTERS_reg[28][17]  ( .G(N2355), .D(N4120), .Q(
        \REGISTERS[28][17] ) );
  DLH_X1 \REGISTERS_reg[28][16]  ( .G(N2355), .D(N4118), .Q(
        \REGISTERS[28][16] ) );
  DLH_X1 \REGISTERS_reg[28][15]  ( .G(N2355), .D(N4116), .Q(
        \REGISTERS[28][15] ) );
  DLH_X1 \REGISTERS_reg[28][14]  ( .G(N2355), .D(N4114), .Q(
        \REGISTERS[28][14] ) );
  DLH_X1 \REGISTERS_reg[28][13]  ( .G(N2355), .D(N4112), .Q(
        \REGISTERS[28][13] ) );
  DLH_X1 \REGISTERS_reg[28][12]  ( .G(N2355), .D(N4110), .Q(
        \REGISTERS[28][12] ) );
  DLH_X1 \REGISTERS_reg[28][11]  ( .G(N2355), .D(N4108), .Q(
        \REGISTERS[28][11] ) );
  DLH_X1 \REGISTERS_reg[28][10]  ( .G(N2355), .D(N4106), .Q(
        \REGISTERS[28][10] ) );
  DLH_X1 \REGISTERS_reg[28][9]  ( .G(N2355), .D(N4104), .Q(\REGISTERS[28][9] )
         );
  DLH_X1 \REGISTERS_reg[28][8]  ( .G(N2355), .D(N4102), .Q(\REGISTERS[28][8] )
         );
  DLH_X1 \REGISTERS_reg[28][7]  ( .G(N2355), .D(N4100), .Q(\REGISTERS[28][7] )
         );
  DLH_X1 \REGISTERS_reg[28][6]  ( .G(N2355), .D(N4098), .Q(\REGISTERS[28][6] )
         );
  DLH_X1 \REGISTERS_reg[28][5]  ( .G(N2355), .D(N4096), .Q(\REGISTERS[28][5] )
         );
  DLH_X1 \REGISTERS_reg[28][4]  ( .G(N2355), .D(N4094), .Q(\REGISTERS[28][4] )
         );
  DLH_X1 \REGISTERS_reg[28][3]  ( .G(N2355), .D(N4092), .Q(\REGISTERS[28][3] )
         );
  DLH_X1 \REGISTERS_reg[28][2]  ( .G(N2355), .D(N4090), .Q(\REGISTERS[28][2] )
         );
  DLH_X1 \REGISTERS_reg[28][1]  ( .G(N2355), .D(N4088), .Q(\REGISTERS[28][1] )
         );
  DLH_X1 \REGISTERS_reg[28][0]  ( .G(N2355), .D(N4086), .Q(\REGISTERS[28][0] )
         );
  DLH_X1 \REGISTERS_reg[29][31]  ( .G(N2291), .D(N4148), .Q(
        \REGISTERS[29][31] ) );
  DLH_X1 \REGISTERS_reg[29][30]  ( .G(N2291), .D(N4146), .Q(
        \REGISTERS[29][30] ) );
  DLH_X1 \REGISTERS_reg[29][29]  ( .G(N2291), .D(N4144), .Q(
        \REGISTERS[29][29] ) );
  DLH_X1 \REGISTERS_reg[29][28]  ( .G(N2291), .D(N4142), .Q(
        \REGISTERS[29][28] ) );
  DLH_X1 \REGISTERS_reg[29][27]  ( .G(N2291), .D(N4140), .Q(
        \REGISTERS[29][27] ) );
  DLH_X1 \REGISTERS_reg[29][26]  ( .G(N2291), .D(N4138), .Q(
        \REGISTERS[29][26] ) );
  DLH_X1 \REGISTERS_reg[29][25]  ( .G(N2291), .D(N4136), .Q(
        \REGISTERS[29][25] ) );
  DLH_X1 \REGISTERS_reg[29][24]  ( .G(N2291), .D(N4134), .Q(
        \REGISTERS[29][24] ) );
  DLH_X1 \REGISTERS_reg[29][23]  ( .G(N2291), .D(N4132), .Q(
        \REGISTERS[29][23] ) );
  DLH_X1 \REGISTERS_reg[29][22]  ( .G(N2291), .D(N4130), .Q(
        \REGISTERS[29][22] ) );
  DLH_X1 \REGISTERS_reg[29][21]  ( .G(N2291), .D(N4128), .Q(
        \REGISTERS[29][21] ) );
  DLH_X1 \REGISTERS_reg[29][20]  ( .G(N2291), .D(N4126), .Q(
        \REGISTERS[29][20] ) );
  DLH_X1 \REGISTERS_reg[29][19]  ( .G(N2291), .D(N4124), .Q(
        \REGISTERS[29][19] ) );
  DLH_X1 \REGISTERS_reg[29][18]  ( .G(N2291), .D(N4122), .Q(
        \REGISTERS[29][18] ) );
  DLH_X1 \REGISTERS_reg[29][17]  ( .G(N2291), .D(N4120), .Q(
        \REGISTERS[29][17] ) );
  DLH_X1 \REGISTERS_reg[29][16]  ( .G(N2291), .D(N4118), .Q(
        \REGISTERS[29][16] ) );
  DLH_X1 \REGISTERS_reg[29][15]  ( .G(N2291), .D(N4116), .Q(
        \REGISTERS[29][15] ) );
  DLH_X1 \REGISTERS_reg[29][14]  ( .G(N2291), .D(N4114), .Q(
        \REGISTERS[29][14] ) );
  DLH_X1 \REGISTERS_reg[29][13]  ( .G(N2291), .D(N4112), .Q(
        \REGISTERS[29][13] ) );
  DLH_X1 \REGISTERS_reg[29][12]  ( .G(N2291), .D(N4110), .Q(
        \REGISTERS[29][12] ) );
  DLH_X1 \REGISTERS_reg[29][11]  ( .G(N2291), .D(N4108), .Q(
        \REGISTERS[29][11] ) );
  DLH_X1 \REGISTERS_reg[29][10]  ( .G(N2291), .D(N4106), .Q(
        \REGISTERS[29][10] ) );
  DLH_X1 \REGISTERS_reg[29][9]  ( .G(N2291), .D(N4104), .Q(\REGISTERS[29][9] )
         );
  DLH_X1 \REGISTERS_reg[29][8]  ( .G(N2291), .D(N4102), .Q(\REGISTERS[29][8] )
         );
  DLH_X1 \REGISTERS_reg[29][7]  ( .G(N2291), .D(N4100), .Q(\REGISTERS[29][7] )
         );
  DLH_X1 \REGISTERS_reg[29][6]  ( .G(N2291), .D(N4098), .Q(\REGISTERS[29][6] )
         );
  DLH_X1 \REGISTERS_reg[29][5]  ( .G(N2291), .D(N4096), .Q(\REGISTERS[29][5] )
         );
  DLH_X1 \REGISTERS_reg[29][4]  ( .G(N2291), .D(N4094), .Q(\REGISTERS[29][4] )
         );
  DLH_X1 \REGISTERS_reg[29][3]  ( .G(N2291), .D(N4092), .Q(\REGISTERS[29][3] )
         );
  DLH_X1 \REGISTERS_reg[29][2]  ( .G(N2291), .D(N4090), .Q(\REGISTERS[29][2] )
         );
  DLH_X1 \REGISTERS_reg[29][1]  ( .G(N2291), .D(N4088), .Q(\REGISTERS[29][1] )
         );
  DLH_X1 \REGISTERS_reg[29][0]  ( .G(N2291), .D(N4086), .Q(\REGISTERS[29][0] )
         );
  DLH_X1 \REGISTERS_reg[30][31]  ( .G(N2227), .D(N4148), .Q(
        \REGISTERS[30][31] ) );
  DLH_X1 \REGISTERS_reg[30][30]  ( .G(N2227), .D(N4146), .Q(
        \REGISTERS[30][30] ) );
  DLH_X1 \REGISTERS_reg[30][29]  ( .G(N2227), .D(N4144), .Q(
        \REGISTERS[30][29] ) );
  DLH_X1 \REGISTERS_reg[30][28]  ( .G(N2227), .D(N4142), .Q(
        \REGISTERS[30][28] ) );
  DLH_X1 \REGISTERS_reg[30][27]  ( .G(N2227), .D(N4140), .Q(
        \REGISTERS[30][27] ) );
  DLH_X1 \REGISTERS_reg[30][26]  ( .G(N2227), .D(N4138), .Q(
        \REGISTERS[30][26] ) );
  DLH_X1 \REGISTERS_reg[30][25]  ( .G(N2227), .D(N4136), .Q(
        \REGISTERS[30][25] ) );
  DLH_X1 \REGISTERS_reg[30][24]  ( .G(N2227), .D(N4134), .Q(
        \REGISTERS[30][24] ) );
  DLH_X1 \REGISTERS_reg[30][23]  ( .G(N2227), .D(N4132), .Q(
        \REGISTERS[30][23] ) );
  DLH_X1 \REGISTERS_reg[30][22]  ( .G(N2227), .D(N4130), .Q(
        \REGISTERS[30][22] ) );
  DLH_X1 \REGISTERS_reg[30][21]  ( .G(N2227), .D(N4128), .Q(
        \REGISTERS[30][21] ) );
  DLH_X1 \REGISTERS_reg[30][20]  ( .G(N2227), .D(N4126), .Q(
        \REGISTERS[30][20] ) );
  DLH_X1 \REGISTERS_reg[30][19]  ( .G(N2227), .D(N4124), .Q(
        \REGISTERS[30][19] ) );
  DLH_X1 \REGISTERS_reg[30][18]  ( .G(N2227), .D(N4122), .Q(
        \REGISTERS[30][18] ) );
  DLH_X1 \REGISTERS_reg[30][17]  ( .G(N2227), .D(N4120), .Q(
        \REGISTERS[30][17] ) );
  DLH_X1 \REGISTERS_reg[30][16]  ( .G(N2227), .D(N4118), .Q(
        \REGISTERS[30][16] ) );
  DLH_X1 \REGISTERS_reg[30][15]  ( .G(N2227), .D(N4116), .Q(
        \REGISTERS[30][15] ) );
  DLH_X1 \REGISTERS_reg[30][14]  ( .G(N2227), .D(N4114), .Q(
        \REGISTERS[30][14] ) );
  DLH_X1 \REGISTERS_reg[30][13]  ( .G(N2227), .D(N4112), .Q(
        \REGISTERS[30][13] ) );
  DLH_X1 \REGISTERS_reg[30][12]  ( .G(N2227), .D(N4110), .Q(
        \REGISTERS[30][12] ) );
  DLH_X1 \REGISTERS_reg[30][11]  ( .G(N2227), .D(N4108), .Q(
        \REGISTERS[30][11] ) );
  DLH_X1 \REGISTERS_reg[30][10]  ( .G(N2227), .D(N4106), .Q(
        \REGISTERS[30][10] ) );
  DLH_X1 \REGISTERS_reg[30][9]  ( .G(N2227), .D(N4104), .Q(\REGISTERS[30][9] )
         );
  DLH_X1 \REGISTERS_reg[30][8]  ( .G(N2227), .D(N4102), .Q(\REGISTERS[30][8] )
         );
  DLH_X1 \REGISTERS_reg[30][7]  ( .G(N2227), .D(N4100), .Q(\REGISTERS[30][7] )
         );
  DLH_X1 \REGISTERS_reg[30][6]  ( .G(N2227), .D(N4098), .Q(\REGISTERS[30][6] )
         );
  DLH_X1 \REGISTERS_reg[30][5]  ( .G(N2227), .D(N4096), .Q(\REGISTERS[30][5] )
         );
  DLH_X1 \REGISTERS_reg[30][4]  ( .G(N2227), .D(N4094), .Q(\REGISTERS[30][4] )
         );
  DLH_X1 \REGISTERS_reg[30][3]  ( .G(N2227), .D(N4092), .Q(\REGISTERS[30][3] )
         );
  DLH_X1 \REGISTERS_reg[30][2]  ( .G(N2227), .D(N4090), .Q(\REGISTERS[30][2] )
         );
  DLH_X1 \REGISTERS_reg[30][1]  ( .G(N2227), .D(N4088), .Q(\REGISTERS[30][1] )
         );
  DLH_X1 \REGISTERS_reg[30][0]  ( .G(N2227), .D(N4086), .Q(\REGISTERS[30][0] )
         );
  DLH_X1 \REGISTERS_reg[31][31]  ( .G(N2163), .D(N4148), .Q(
        \REGISTERS[31][31] ) );
  DLH_X1 \REGISTERS_reg[31][30]  ( .G(N2163), .D(N4146), .Q(
        \REGISTERS[31][30] ) );
  DLH_X1 \REGISTERS_reg[31][29]  ( .G(N2163), .D(N4144), .Q(
        \REGISTERS[31][29] ) );
  DLH_X1 \REGISTERS_reg[31][28]  ( .G(N2163), .D(N4142), .Q(
        \REGISTERS[31][28] ) );
  DLH_X1 \REGISTERS_reg[31][27]  ( .G(N2163), .D(N4140), .Q(
        \REGISTERS[31][27] ) );
  DLH_X1 \REGISTERS_reg[31][26]  ( .G(N2163), .D(N4138), .Q(
        \REGISTERS[31][26] ) );
  DLH_X1 \REGISTERS_reg[31][25]  ( .G(N2163), .D(N4136), .Q(
        \REGISTERS[31][25] ) );
  DLH_X1 \REGISTERS_reg[31][24]  ( .G(N2163), .D(N4134), .Q(
        \REGISTERS[31][24] ) );
  DLH_X1 \REGISTERS_reg[31][23]  ( .G(N2163), .D(N4132), .Q(
        \REGISTERS[31][23] ) );
  DLH_X1 \REGISTERS_reg[31][22]  ( .G(N2163), .D(N4130), .Q(
        \REGISTERS[31][22] ) );
  DLH_X1 \REGISTERS_reg[31][21]  ( .G(N2163), .D(N4128), .Q(
        \REGISTERS[31][21] ) );
  DLH_X1 \REGISTERS_reg[31][20]  ( .G(N2163), .D(N4126), .Q(
        \REGISTERS[31][20] ) );
  DLH_X1 \REGISTERS_reg[31][19]  ( .G(N2163), .D(N4124), .Q(
        \REGISTERS[31][19] ) );
  DLH_X1 \REGISTERS_reg[31][18]  ( .G(N2163), .D(N4122), .Q(
        \REGISTERS[31][18] ) );
  DLH_X1 \REGISTERS_reg[31][17]  ( .G(N2163), .D(N4120), .Q(
        \REGISTERS[31][17] ) );
  DLH_X1 \REGISTERS_reg[31][16]  ( .G(N2163), .D(N4118), .Q(
        \REGISTERS[31][16] ) );
  DLH_X1 \REGISTERS_reg[31][15]  ( .G(N2163), .D(N4116), .Q(
        \REGISTERS[31][15] ) );
  DLH_X1 \REGISTERS_reg[31][14]  ( .G(N2163), .D(N4114), .Q(
        \REGISTERS[31][14] ) );
  DLH_X1 \REGISTERS_reg[31][13]  ( .G(N2163), .D(N4112), .Q(
        \REGISTERS[31][13] ) );
  DLH_X1 \REGISTERS_reg[31][12]  ( .G(N2163), .D(N4110), .Q(
        \REGISTERS[31][12] ) );
  DLH_X1 \REGISTERS_reg[31][11]  ( .G(N2163), .D(N4108), .Q(
        \REGISTERS[31][11] ) );
  DLH_X1 \REGISTERS_reg[31][10]  ( .G(N2163), .D(N4106), .Q(
        \REGISTERS[31][10] ) );
  DLH_X1 \REGISTERS_reg[31][9]  ( .G(N2163), .D(N4104), .Q(\REGISTERS[31][9] )
         );
  DLH_X1 \REGISTERS_reg[31][8]  ( .G(N2163), .D(N4102), .Q(\REGISTERS[31][8] )
         );
  DLH_X1 \REGISTERS_reg[31][7]  ( .G(N2163), .D(N4100), .Q(\REGISTERS[31][7] )
         );
  DLH_X1 \REGISTERS_reg[31][6]  ( .G(N2163), .D(N4098), .Q(\REGISTERS[31][6] )
         );
  DLH_X1 \REGISTERS_reg[31][5]  ( .G(N2163), .D(N4096), .Q(\REGISTERS[31][5] )
         );
  DLH_X1 \REGISTERS_reg[31][4]  ( .G(N2163), .D(N4094), .Q(\REGISTERS[31][4] )
         );
  DLH_X1 \REGISTERS_reg[31][3]  ( .G(N2163), .D(N4092), .Q(\REGISTERS[31][3] )
         );
  DLH_X1 \REGISTERS_reg[31][2]  ( .G(N2163), .D(N4090), .Q(\REGISTERS[31][2] )
         );
  DLH_X1 \REGISTERS_reg[31][1]  ( .G(N2163), .D(N4088), .Q(\REGISTERS[31][1] )
         );
  DLH_X1 \REGISTERS_reg[31][0]  ( .G(N2163), .D(N4086), .Q(\REGISTERS[31][0] )
         );
  DLH_X1 \OUT1_reg[31]  ( .G(N4278), .D(N4215), .Q(OUT1[31]) );
  DLH_X1 \OUT1_reg[30]  ( .G(N4278), .D(N4216), .Q(OUT1[30]) );
  DLH_X1 \OUT1_reg[29]  ( .G(N4278), .D(N4217), .Q(OUT1[29]) );
  DLH_X1 \OUT1_reg[28]  ( .G(N4278), .D(N4218), .Q(OUT1[28]) );
  DLH_X1 \OUT1_reg[27]  ( .G(N4278), .D(N4219), .Q(OUT1[27]) );
  DLH_X1 \OUT1_reg[26]  ( .G(N4278), .D(N4220), .Q(OUT1[26]) );
  DLH_X1 \OUT1_reg[25]  ( .G(N4278), .D(N4221), .Q(OUT1[25]) );
  DLH_X1 \OUT1_reg[24]  ( .G(N4278), .D(N4222), .Q(OUT1[24]) );
  DLH_X1 \OUT1_reg[23]  ( .G(N4278), .D(N4223), .Q(OUT1[23]) );
  DLH_X1 \OUT1_reg[22]  ( .G(N4278), .D(N4224), .Q(OUT1[22]) );
  DLH_X1 \OUT1_reg[21]  ( .G(N4278), .D(N4225), .Q(OUT1[21]) );
  DLH_X1 \OUT1_reg[20]  ( .G(N4278), .D(N4226), .Q(OUT1[20]) );
  DLH_X1 \OUT1_reg[19]  ( .G(N4278), .D(N4227), .Q(OUT1[19]) );
  DLH_X1 \OUT1_reg[18]  ( .G(N4278), .D(N4228), .Q(OUT1[18]) );
  DLH_X1 \OUT1_reg[17]  ( .G(N4278), .D(N4229), .Q(OUT1[17]) );
  DLH_X1 \OUT1_reg[16]  ( .G(N4278), .D(N4230), .Q(OUT1[16]) );
  DLH_X1 \OUT1_reg[15]  ( .G(N4278), .D(N4231), .Q(OUT1[15]) );
  DLH_X1 \OUT1_reg[14]  ( .G(N4278), .D(N4232), .Q(OUT1[14]) );
  DLH_X1 \OUT1_reg[13]  ( .G(N4278), .D(N4233), .Q(OUT1[13]) );
  DLH_X1 \OUT1_reg[12]  ( .G(N4278), .D(N4234), .Q(OUT1[12]) );
  DLH_X1 \OUT1_reg[11]  ( .G(N4278), .D(N4235), .Q(OUT1[11]) );
  DLH_X1 \OUT1_reg[10]  ( .G(N4278), .D(N4236), .Q(OUT1[10]) );
  DLH_X1 \OUT1_reg[9]  ( .G(N4278), .D(N4237), .Q(OUT1[9]) );
  DLH_X1 \OUT1_reg[8]  ( .G(N4278), .D(N4238), .Q(OUT1[8]) );
  DLH_X1 \OUT1_reg[7]  ( .G(N4278), .D(N4239), .Q(OUT1[7]) );
  DLH_X1 \OUT1_reg[6]  ( .G(N4278), .D(N4240), .Q(OUT1[6]) );
  DLH_X1 \OUT1_reg[5]  ( .G(N4278), .D(N4241), .Q(OUT1[5]) );
  DLH_X1 \OUT1_reg[4]  ( .G(N4278), .D(N4242), .Q(OUT1[4]) );
  DLH_X1 \OUT1_reg[3]  ( .G(N4278), .D(N4243), .Q(OUT1[3]) );
  DLH_X1 \OUT1_reg[2]  ( .G(N4278), .D(N4244), .Q(OUT1[2]) );
  DLH_X1 \OUT1_reg[1]  ( .G(N4278), .D(N4245), .Q(OUT1[1]) );
  DLH_X1 \OUT1_reg[0]  ( .G(N4278), .D(N4246), .Q(OUT1[0]) );
  DLH_X1 \OUT2_reg[31]  ( .G(N4407), .D(N4344), .Q(OUT2[31]) );
  DLH_X1 \OUT2_reg[30]  ( .G(N4407), .D(N4345), .Q(OUT2[30]) );
  DLH_X1 \OUT2_reg[29]  ( .G(N4407), .D(N4346), .Q(OUT2[29]) );
  DLH_X1 \OUT2_reg[28]  ( .G(N4407), .D(N4347), .Q(OUT2[28]) );
  DLH_X1 \OUT2_reg[27]  ( .G(N4407), .D(N4348), .Q(OUT2[27]) );
  DLH_X1 \OUT2_reg[26]  ( .G(N4407), .D(N4349), .Q(OUT2[26]) );
  DLH_X1 \OUT2_reg[25]  ( .G(N4407), .D(N4350), .Q(OUT2[25]) );
  DLH_X1 \OUT2_reg[24]  ( .G(N4407), .D(N4351), .Q(OUT2[24]) );
  DLH_X1 \OUT2_reg[23]  ( .G(N4407), .D(N4352), .Q(OUT2[23]) );
  DLH_X1 \OUT2_reg[22]  ( .G(N4407), .D(N4353), .Q(OUT2[22]) );
  DLH_X1 \OUT2_reg[21]  ( .G(N4407), .D(N4354), .Q(OUT2[21]) );
  DLH_X1 \OUT2_reg[20]  ( .G(N4407), .D(N4355), .Q(OUT2[20]) );
  DLH_X1 \OUT2_reg[19]  ( .G(N4407), .D(N4356), .Q(OUT2[19]) );
  DLH_X1 \OUT2_reg[18]  ( .G(N4407), .D(N4357), .Q(OUT2[18]) );
  DLH_X1 \OUT2_reg[17]  ( .G(N4407), .D(N4358), .Q(OUT2[17]) );
  DLH_X1 \OUT2_reg[16]  ( .G(N4407), .D(N4359), .Q(OUT2[16]) );
  DLH_X1 \OUT2_reg[15]  ( .G(N4407), .D(N4360), .Q(OUT2[15]) );
  DLH_X1 \OUT2_reg[14]  ( .G(N4407), .D(N4361), .Q(OUT2[14]) );
  DLH_X1 \OUT2_reg[13]  ( .G(N4407), .D(N4362), .Q(OUT2[13]) );
  DLH_X1 \OUT2_reg[12]  ( .G(N4407), .D(N4363), .Q(OUT2[12]) );
  DLH_X1 \OUT2_reg[11]  ( .G(N4407), .D(N4364), .Q(OUT2[11]) );
  DLH_X1 \OUT2_reg[10]  ( .G(N4407), .D(N4365), .Q(OUT2[10]) );
  DLH_X1 \OUT2_reg[9]  ( .G(N4407), .D(N4366), .Q(OUT2[9]) );
  DLH_X1 \OUT2_reg[8]  ( .G(N4407), .D(N4367), .Q(OUT2[8]) );
  DLH_X1 \OUT2_reg[7]  ( .G(N4407), .D(N4368), .Q(OUT2[7]) );
  DLH_X1 \OUT2_reg[6]  ( .G(N4407), .D(N4369), .Q(OUT2[6]) );
  DLH_X1 \OUT2_reg[5]  ( .G(N4407), .D(N4370), .Q(OUT2[5]) );
  DLH_X1 \OUT2_reg[4]  ( .G(N4407), .D(N4371), .Q(OUT2[4]) );
  DLH_X1 \OUT2_reg[3]  ( .G(N4407), .D(N4372), .Q(OUT2[3]) );
  DLH_X1 \OUT2_reg[2]  ( .G(N4407), .D(N4373), .Q(OUT2[2]) );
  DLH_X1 \OUT2_reg[1]  ( .G(N4407), .D(N4374), .Q(OUT2[1]) );
  DLH_X1 \OUT2_reg[0]  ( .G(N4407), .D(N4375), .Q(OUT2[0]) );
  AND2_X1 U35 ( .A1(RD2), .A2(ENABLE), .ZN(N4407) );
  NAND2_X1 U36 ( .A1(n2), .A2(n3), .ZN(N4375) );
  NOR4_X1 U37 ( .A1(n4), .A2(n5), .A3(n6), .A4(n7), .ZN(n3) );
  OAI221_X1 U38 ( .B1(n8), .B2(n9), .C1(n10), .C2(n11), .A(n12), .ZN(n7) );
  AOI22_X1 U39 ( .A1(\REGISTERS[19][0] ), .A2(n13), .B1(\REGISTERS[18][0] ), 
        .B2(n14), .ZN(n12) );
  OAI221_X1 U40 ( .B1(n15), .B2(n16), .C1(n17), .C2(n18), .A(n19), .ZN(n6) );
  AOI22_X1 U41 ( .A1(\REGISTERS[23][0] ), .A2(n20), .B1(\REGISTERS[22][0] ), 
        .B2(n21), .ZN(n19) );
  OAI221_X1 U42 ( .B1(n22), .B2(n23), .C1(n24), .C2(n25), .A(n26), .ZN(n5) );
  AOI22_X1 U43 ( .A1(\REGISTERS[27][0] ), .A2(n27), .B1(\REGISTERS[26][0] ), 
        .B2(n28), .ZN(n26) );
  OAI221_X1 U44 ( .B1(n29), .B2(n30), .C1(n31), .C2(n32), .A(n33), .ZN(n4) );
  AOI22_X1 U45 ( .A1(\REGISTERS[29][0] ), .A2(n34), .B1(\REGISTERS[28][0] ), 
        .B2(n35), .ZN(n33) );
  NOR4_X1 U46 ( .A1(n36), .A2(n37), .A3(n38), .A4(n39), .ZN(n2) );
  AOI22_X1 U48 ( .A1(\REGISTERS[3][0] ), .A2(n45), .B1(\REGISTERS[2][0] ), 
        .B2(n46), .ZN(n44) );
  OAI221_X1 U49 ( .B1(n47), .B2(n48), .C1(n49), .C2(n50), .A(n51), .ZN(n38) );
  AOI22_X1 U50 ( .A1(\REGISTERS[7][0] ), .A2(n52), .B1(\REGISTERS[6][0] ), 
        .B2(n53), .ZN(n51) );
  OAI221_X1 U51 ( .B1(n54), .B2(n55), .C1(n56), .C2(n57), .A(n58), .ZN(n37) );
  AOI22_X1 U52 ( .A1(\REGISTERS[11][0] ), .A2(n59), .B1(\REGISTERS[10][0] ), 
        .B2(n60), .ZN(n58) );
  OAI221_X1 U53 ( .B1(n61), .B2(n62), .C1(n63), .C2(n64), .A(n65), .ZN(n36) );
  AOI22_X1 U54 ( .A1(\REGISTERS[15][0] ), .A2(n66), .B1(\REGISTERS[14][0] ), 
        .B2(n67), .ZN(n65) );
  NAND2_X1 U55 ( .A1(n68), .A2(n69), .ZN(N4374) );
  NOR4_X1 U56 ( .A1(n70), .A2(n71), .A3(n72), .A4(n73), .ZN(n69) );
  OAI221_X1 U57 ( .B1(n8), .B2(n74), .C1(n10), .C2(n75), .A(n76), .ZN(n73) );
  AOI22_X1 U58 ( .A1(\REGISTERS[19][1] ), .A2(n13), .B1(\REGISTERS[18][1] ), 
        .B2(n14), .ZN(n76) );
  OAI221_X1 U59 ( .B1(n15), .B2(n77), .C1(n17), .C2(n78), .A(n79), .ZN(n72) );
  AOI22_X1 U60 ( .A1(\REGISTERS[23][1] ), .A2(n20), .B1(\REGISTERS[22][1] ), 
        .B2(n21), .ZN(n79) );
  OAI221_X1 U61 ( .B1(n22), .B2(n80), .C1(n24), .C2(n81), .A(n82), .ZN(n71) );
  AOI22_X1 U62 ( .A1(\REGISTERS[27][1] ), .A2(n27), .B1(\REGISTERS[26][1] ), 
        .B2(n28), .ZN(n82) );
  OAI221_X1 U63 ( .B1(n29), .B2(n83), .C1(n31), .C2(n84), .A(n85), .ZN(n70) );
  AOI22_X1 U64 ( .A1(\REGISTERS[29][1] ), .A2(n34), .B1(\REGISTERS[28][1] ), 
        .B2(n35), .ZN(n85) );
  NOR4_X1 U65 ( .A1(n86), .A2(n87), .A3(n88), .A4(n89), .ZN(n68) );
  AOI22_X1 U67 ( .A1(\REGISTERS[3][1] ), .A2(n45), .B1(\REGISTERS[2][1] ), 
        .B2(n46), .ZN(n92) );
  OAI221_X1 U68 ( .B1(n47), .B2(n93), .C1(n49), .C2(n94), .A(n95), .ZN(n88) );
  AOI22_X1 U69 ( .A1(\REGISTERS[7][1] ), .A2(n52), .B1(\REGISTERS[6][1] ), 
        .B2(n53), .ZN(n95) );
  OAI221_X1 U70 ( .B1(n54), .B2(n96), .C1(n56), .C2(n97), .A(n98), .ZN(n87) );
  AOI22_X1 U71 ( .A1(\REGISTERS[11][1] ), .A2(n59), .B1(\REGISTERS[10][1] ), 
        .B2(n60), .ZN(n98) );
  OAI221_X1 U72 ( .B1(n61), .B2(n99), .C1(n63), .C2(n100), .A(n101), .ZN(n86)
         );
  AOI22_X1 U73 ( .A1(\REGISTERS[15][1] ), .A2(n66), .B1(\REGISTERS[14][1] ), 
        .B2(n67), .ZN(n101) );
  NAND2_X1 U74 ( .A1(n102), .A2(n103), .ZN(N4373) );
  NOR4_X1 U75 ( .A1(n104), .A2(n105), .A3(n106), .A4(n107), .ZN(n103) );
  OAI221_X1 U76 ( .B1(n8), .B2(n108), .C1(n10), .C2(n109), .A(n110), .ZN(n107)
         );
  AOI22_X1 U77 ( .A1(\REGISTERS[19][2] ), .A2(n13), .B1(\REGISTERS[18][2] ), 
        .B2(n14), .ZN(n110) );
  OAI221_X1 U78 ( .B1(n15), .B2(n111), .C1(n17), .C2(n112), .A(n113), .ZN(n106) );
  AOI22_X1 U79 ( .A1(\REGISTERS[23][2] ), .A2(n20), .B1(\REGISTERS[22][2] ), 
        .B2(n21), .ZN(n113) );
  OAI221_X1 U80 ( .B1(n22), .B2(n114), .C1(n24), .C2(n115), .A(n116), .ZN(n105) );
  AOI22_X1 U81 ( .A1(\REGISTERS[27][2] ), .A2(n27), .B1(\REGISTERS[26][2] ), 
        .B2(n28), .ZN(n116) );
  OAI221_X1 U82 ( .B1(n29), .B2(n117), .C1(n31), .C2(n118), .A(n119), .ZN(n104) );
  AOI22_X1 U83 ( .A1(\REGISTERS[29][2] ), .A2(n34), .B1(\REGISTERS[28][2] ), 
        .B2(n35), .ZN(n119) );
  NOR4_X1 U84 ( .A1(n120), .A2(n121), .A3(n122), .A4(n123), .ZN(n102) );
  AOI22_X1 U86 ( .A1(\REGISTERS[3][2] ), .A2(n45), .B1(\REGISTERS[2][2] ), 
        .B2(n46), .ZN(n126) );
  OAI221_X1 U87 ( .B1(n47), .B2(n127), .C1(n49), .C2(n128), .A(n129), .ZN(n122) );
  AOI22_X1 U88 ( .A1(\REGISTERS[7][2] ), .A2(n52), .B1(\REGISTERS[6][2] ), 
        .B2(n53), .ZN(n129) );
  OAI221_X1 U89 ( .B1(n54), .B2(n130), .C1(n56), .C2(n131), .A(n132), .ZN(n121) );
  AOI22_X1 U90 ( .A1(\REGISTERS[11][2] ), .A2(n59), .B1(\REGISTERS[10][2] ), 
        .B2(n60), .ZN(n132) );
  OAI221_X1 U91 ( .B1(n61), .B2(n133), .C1(n63), .C2(n134), .A(n135), .ZN(n120) );
  AOI22_X1 U92 ( .A1(\REGISTERS[15][2] ), .A2(n66), .B1(\REGISTERS[14][2] ), 
        .B2(n67), .ZN(n135) );
  NAND2_X1 U93 ( .A1(n136), .A2(n137), .ZN(N4372) );
  NOR4_X1 U94 ( .A1(n138), .A2(n139), .A3(n140), .A4(n141), .ZN(n137) );
  OAI221_X1 U95 ( .B1(n8), .B2(n142), .C1(n10), .C2(n143), .A(n144), .ZN(n141)
         );
  AOI22_X1 U96 ( .A1(\REGISTERS[19][3] ), .A2(n13), .B1(\REGISTERS[18][3] ), 
        .B2(n14), .ZN(n144) );
  OAI221_X1 U97 ( .B1(n15), .B2(n145), .C1(n17), .C2(n146), .A(n147), .ZN(n140) );
  AOI22_X1 U98 ( .A1(\REGISTERS[23][3] ), .A2(n20), .B1(\REGISTERS[22][3] ), 
        .B2(n21), .ZN(n147) );
  OAI221_X1 U99 ( .B1(n22), .B2(n148), .C1(n24), .C2(n149), .A(n150), .ZN(n139) );
  AOI22_X1 U100 ( .A1(\REGISTERS[27][3] ), .A2(n27), .B1(\REGISTERS[26][3] ), 
        .B2(n28), .ZN(n150) );
  OAI221_X1 U101 ( .B1(n29), .B2(n151), .C1(n31), .C2(n152), .A(n153), .ZN(
        n138) );
  AOI22_X1 U102 ( .A1(\REGISTERS[29][3] ), .A2(n34), .B1(\REGISTERS[28][3] ), 
        .B2(n35), .ZN(n153) );
  NOR4_X1 U103 ( .A1(n154), .A2(n155), .A3(n156), .A4(n157), .ZN(n136) );
  AOI22_X1 U105 ( .A1(\REGISTERS[3][3] ), .A2(n45), .B1(\REGISTERS[2][3] ), 
        .B2(n46), .ZN(n160) );
  OAI221_X1 U106 ( .B1(n47), .B2(n161), .C1(n49), .C2(n162), .A(n163), .ZN(
        n156) );
  AOI22_X1 U107 ( .A1(\REGISTERS[7][3] ), .A2(n52), .B1(\REGISTERS[6][3] ), 
        .B2(n53), .ZN(n163) );
  OAI221_X1 U108 ( .B1(n54), .B2(n164), .C1(n56), .C2(n165), .A(n166), .ZN(
        n155) );
  AOI22_X1 U109 ( .A1(\REGISTERS[11][3] ), .A2(n59), .B1(\REGISTERS[10][3] ), 
        .B2(n60), .ZN(n166) );
  OAI221_X1 U110 ( .B1(n61), .B2(n167), .C1(n63), .C2(n168), .A(n169), .ZN(
        n154) );
  AOI22_X1 U111 ( .A1(\REGISTERS[15][3] ), .A2(n66), .B1(\REGISTERS[14][3] ), 
        .B2(n67), .ZN(n169) );
  NAND2_X1 U112 ( .A1(n170), .A2(n171), .ZN(N4371) );
  NOR4_X1 U113 ( .A1(n172), .A2(n173), .A3(n174), .A4(n175), .ZN(n171) );
  OAI221_X1 U114 ( .B1(n8), .B2(n176), .C1(n10), .C2(n177), .A(n178), .ZN(n175) );
  AOI22_X1 U115 ( .A1(\REGISTERS[19][4] ), .A2(n13), .B1(\REGISTERS[18][4] ), 
        .B2(n14), .ZN(n178) );
  OAI221_X1 U116 ( .B1(n15), .B2(n179), .C1(n17), .C2(n180), .A(n181), .ZN(
        n174) );
  AOI22_X1 U117 ( .A1(\REGISTERS[23][4] ), .A2(n20), .B1(\REGISTERS[22][4] ), 
        .B2(n21), .ZN(n181) );
  OAI221_X1 U118 ( .B1(n22), .B2(n182), .C1(n24), .C2(n183), .A(n184), .ZN(
        n173) );
  AOI22_X1 U119 ( .A1(\REGISTERS[27][4] ), .A2(n27), .B1(\REGISTERS[26][4] ), 
        .B2(n28), .ZN(n184) );
  OAI221_X1 U120 ( .B1(n29), .B2(n185), .C1(n31), .C2(n186), .A(n187), .ZN(
        n172) );
  AOI22_X1 U121 ( .A1(\REGISTERS[29][4] ), .A2(n34), .B1(\REGISTERS[28][4] ), 
        .B2(n35), .ZN(n187) );
  NOR4_X1 U122 ( .A1(n188), .A2(n189), .A3(n190), .A4(n191), .ZN(n170) );
  AOI22_X1 U124 ( .A1(\REGISTERS[3][4] ), .A2(n45), .B1(\REGISTERS[2][4] ), 
        .B2(n46), .ZN(n194) );
  OAI221_X1 U125 ( .B1(n47), .B2(n195), .C1(n49), .C2(n196), .A(n197), .ZN(
        n190) );
  AOI22_X1 U126 ( .A1(\REGISTERS[7][4] ), .A2(n52), .B1(\REGISTERS[6][4] ), 
        .B2(n53), .ZN(n197) );
  OAI221_X1 U127 ( .B1(n54), .B2(n198), .C1(n56), .C2(n199), .A(n200), .ZN(
        n189) );
  AOI22_X1 U128 ( .A1(\REGISTERS[11][4] ), .A2(n59), .B1(\REGISTERS[10][4] ), 
        .B2(n60), .ZN(n200) );
  OAI221_X1 U129 ( .B1(n61), .B2(n201), .C1(n63), .C2(n202), .A(n203), .ZN(
        n188) );
  AOI22_X1 U130 ( .A1(\REGISTERS[15][4] ), .A2(n66), .B1(\REGISTERS[14][4] ), 
        .B2(n67), .ZN(n203) );
  NAND2_X1 U131 ( .A1(n204), .A2(n205), .ZN(N4370) );
  NOR4_X1 U132 ( .A1(n206), .A2(n207), .A3(n208), .A4(n209), .ZN(n205) );
  OAI221_X1 U133 ( .B1(n8), .B2(n210), .C1(n10), .C2(n211), .A(n212), .ZN(n209) );
  AOI22_X1 U134 ( .A1(\REGISTERS[19][5] ), .A2(n13), .B1(\REGISTERS[18][5] ), 
        .B2(n14), .ZN(n212) );
  OAI221_X1 U135 ( .B1(n15), .B2(n213), .C1(n17), .C2(n214), .A(n215), .ZN(
        n208) );
  AOI22_X1 U136 ( .A1(\REGISTERS[23][5] ), .A2(n20), .B1(\REGISTERS[22][5] ), 
        .B2(n21), .ZN(n215) );
  OAI221_X1 U137 ( .B1(n22), .B2(n216), .C1(n24), .C2(n217), .A(n218), .ZN(
        n207) );
  AOI22_X1 U138 ( .A1(\REGISTERS[27][5] ), .A2(n27), .B1(\REGISTERS[26][5] ), 
        .B2(n28), .ZN(n218) );
  OAI221_X1 U139 ( .B1(n29), .B2(n219), .C1(n31), .C2(n220), .A(n221), .ZN(
        n206) );
  AOI22_X1 U140 ( .A1(\REGISTERS[29][5] ), .A2(n34), .B1(\REGISTERS[28][5] ), 
        .B2(n35), .ZN(n221) );
  NOR4_X1 U141 ( .A1(n222), .A2(n223), .A3(n224), .A4(n225), .ZN(n204) );
  AOI22_X1 U143 ( .A1(\REGISTERS[3][5] ), .A2(n45), .B1(\REGISTERS[2][5] ), 
        .B2(n46), .ZN(n228) );
  OAI221_X1 U144 ( .B1(n47), .B2(n229), .C1(n49), .C2(n230), .A(n231), .ZN(
        n224) );
  AOI22_X1 U145 ( .A1(\REGISTERS[7][5] ), .A2(n52), .B1(\REGISTERS[6][5] ), 
        .B2(n53), .ZN(n231) );
  OAI221_X1 U146 ( .B1(n54), .B2(n232), .C1(n56), .C2(n233), .A(n234), .ZN(
        n223) );
  AOI22_X1 U147 ( .A1(\REGISTERS[11][5] ), .A2(n59), .B1(\REGISTERS[10][5] ), 
        .B2(n60), .ZN(n234) );
  OAI221_X1 U148 ( .B1(n61), .B2(n235), .C1(n63), .C2(n236), .A(n237), .ZN(
        n222) );
  AOI22_X1 U149 ( .A1(\REGISTERS[15][5] ), .A2(n66), .B1(\REGISTERS[14][5] ), 
        .B2(n67), .ZN(n237) );
  NAND2_X1 U150 ( .A1(n238), .A2(n239), .ZN(N4369) );
  NOR4_X1 U151 ( .A1(n240), .A2(n241), .A3(n242), .A4(n243), .ZN(n239) );
  OAI221_X1 U152 ( .B1(n8), .B2(n244), .C1(n10), .C2(n245), .A(n246), .ZN(n243) );
  AOI22_X1 U153 ( .A1(\REGISTERS[19][6] ), .A2(n13), .B1(\REGISTERS[18][6] ), 
        .B2(n14), .ZN(n246) );
  OAI221_X1 U154 ( .B1(n15), .B2(n247), .C1(n17), .C2(n248), .A(n249), .ZN(
        n242) );
  AOI22_X1 U155 ( .A1(\REGISTERS[23][6] ), .A2(n20), .B1(\REGISTERS[22][6] ), 
        .B2(n21), .ZN(n249) );
  OAI221_X1 U156 ( .B1(n22), .B2(n250), .C1(n24), .C2(n251), .A(n252), .ZN(
        n241) );
  AOI22_X1 U157 ( .A1(\REGISTERS[27][6] ), .A2(n27), .B1(\REGISTERS[26][6] ), 
        .B2(n28), .ZN(n252) );
  OAI221_X1 U158 ( .B1(n29), .B2(n253), .C1(n31), .C2(n254), .A(n255), .ZN(
        n240) );
  AOI22_X1 U159 ( .A1(\REGISTERS[29][6] ), .A2(n34), .B1(\REGISTERS[28][6] ), 
        .B2(n35), .ZN(n255) );
  NOR4_X1 U160 ( .A1(n256), .A2(n257), .A3(n258), .A4(n259), .ZN(n238) );
  AOI22_X1 U162 ( .A1(\REGISTERS[3][6] ), .A2(n45), .B1(\REGISTERS[2][6] ), 
        .B2(n46), .ZN(n262) );
  OAI221_X1 U163 ( .B1(n47), .B2(n263), .C1(n49), .C2(n264), .A(n265), .ZN(
        n258) );
  AOI22_X1 U164 ( .A1(\REGISTERS[7][6] ), .A2(n52), .B1(\REGISTERS[6][6] ), 
        .B2(n53), .ZN(n265) );
  OAI221_X1 U165 ( .B1(n54), .B2(n266), .C1(n56), .C2(n267), .A(n268), .ZN(
        n257) );
  AOI22_X1 U166 ( .A1(\REGISTERS[11][6] ), .A2(n59), .B1(\REGISTERS[10][6] ), 
        .B2(n60), .ZN(n268) );
  OAI221_X1 U167 ( .B1(n61), .B2(n269), .C1(n63), .C2(n270), .A(n271), .ZN(
        n256) );
  AOI22_X1 U168 ( .A1(\REGISTERS[15][6] ), .A2(n66), .B1(\REGISTERS[14][6] ), 
        .B2(n67), .ZN(n271) );
  NAND2_X1 U169 ( .A1(n272), .A2(n273), .ZN(N4368) );
  NOR4_X1 U170 ( .A1(n274), .A2(n275), .A3(n276), .A4(n277), .ZN(n273) );
  OAI221_X1 U171 ( .B1(n8), .B2(n278), .C1(n10), .C2(n279), .A(n280), .ZN(n277) );
  AOI22_X1 U172 ( .A1(\REGISTERS[19][7] ), .A2(n13), .B1(\REGISTERS[18][7] ), 
        .B2(n14), .ZN(n280) );
  OAI221_X1 U173 ( .B1(n15), .B2(n281), .C1(n17), .C2(n282), .A(n283), .ZN(
        n276) );
  AOI22_X1 U174 ( .A1(\REGISTERS[23][7] ), .A2(n20), .B1(\REGISTERS[22][7] ), 
        .B2(n21), .ZN(n283) );
  OAI221_X1 U175 ( .B1(n22), .B2(n284), .C1(n24), .C2(n285), .A(n286), .ZN(
        n275) );
  AOI22_X1 U176 ( .A1(\REGISTERS[27][7] ), .A2(n27), .B1(\REGISTERS[26][7] ), 
        .B2(n28), .ZN(n286) );
  OAI221_X1 U177 ( .B1(n29), .B2(n287), .C1(n31), .C2(n288), .A(n289), .ZN(
        n274) );
  AOI22_X1 U178 ( .A1(\REGISTERS[29][7] ), .A2(n34), .B1(\REGISTERS[28][7] ), 
        .B2(n35), .ZN(n289) );
  NOR4_X1 U179 ( .A1(n290), .A2(n291), .A3(n292), .A4(n293), .ZN(n272) );
  AOI22_X1 U181 ( .A1(\REGISTERS[3][7] ), .A2(n45), .B1(\REGISTERS[2][7] ), 
        .B2(n46), .ZN(n296) );
  OAI221_X1 U182 ( .B1(n47), .B2(n297), .C1(n49), .C2(n298), .A(n299), .ZN(
        n292) );
  AOI22_X1 U183 ( .A1(\REGISTERS[7][7] ), .A2(n52), .B1(\REGISTERS[6][7] ), 
        .B2(n53), .ZN(n299) );
  OAI221_X1 U184 ( .B1(n54), .B2(n300), .C1(n56), .C2(n301), .A(n302), .ZN(
        n291) );
  AOI22_X1 U185 ( .A1(\REGISTERS[11][7] ), .A2(n59), .B1(\REGISTERS[10][7] ), 
        .B2(n60), .ZN(n302) );
  OAI221_X1 U186 ( .B1(n61), .B2(n303), .C1(n63), .C2(n304), .A(n305), .ZN(
        n290) );
  AOI22_X1 U187 ( .A1(\REGISTERS[15][7] ), .A2(n66), .B1(\REGISTERS[14][7] ), 
        .B2(n67), .ZN(n305) );
  NAND2_X1 U188 ( .A1(n306), .A2(n307), .ZN(N4367) );
  NOR4_X1 U189 ( .A1(n308), .A2(n309), .A3(n310), .A4(n311), .ZN(n307) );
  OAI221_X1 U190 ( .B1(n8), .B2(n312), .C1(n10), .C2(n313), .A(n314), .ZN(n311) );
  AOI22_X1 U191 ( .A1(\REGISTERS[19][8] ), .A2(n13), .B1(\REGISTERS[18][8] ), 
        .B2(n14), .ZN(n314) );
  OAI221_X1 U192 ( .B1(n15), .B2(n315), .C1(n17), .C2(n316), .A(n317), .ZN(
        n310) );
  AOI22_X1 U193 ( .A1(\REGISTERS[23][8] ), .A2(n20), .B1(\REGISTERS[22][8] ), 
        .B2(n21), .ZN(n317) );
  OAI221_X1 U194 ( .B1(n22), .B2(n318), .C1(n24), .C2(n319), .A(n320), .ZN(
        n309) );
  AOI22_X1 U195 ( .A1(\REGISTERS[27][8] ), .A2(n27), .B1(\REGISTERS[26][8] ), 
        .B2(n28), .ZN(n320) );
  OAI221_X1 U196 ( .B1(n29), .B2(n321), .C1(n31), .C2(n322), .A(n323), .ZN(
        n308) );
  AOI22_X1 U197 ( .A1(\REGISTERS[29][8] ), .A2(n34), .B1(\REGISTERS[28][8] ), 
        .B2(n35), .ZN(n323) );
  NOR4_X1 U198 ( .A1(n324), .A2(n325), .A3(n326), .A4(n327), .ZN(n306) );
  AOI22_X1 U200 ( .A1(\REGISTERS[3][8] ), .A2(n45), .B1(\REGISTERS[2][8] ), 
        .B2(n46), .ZN(n330) );
  OAI221_X1 U201 ( .B1(n47), .B2(n331), .C1(n49), .C2(n332), .A(n333), .ZN(
        n326) );
  AOI22_X1 U202 ( .A1(\REGISTERS[7][8] ), .A2(n52), .B1(\REGISTERS[6][8] ), 
        .B2(n53), .ZN(n333) );
  OAI221_X1 U203 ( .B1(n54), .B2(n334), .C1(n56), .C2(n335), .A(n336), .ZN(
        n325) );
  AOI22_X1 U204 ( .A1(\REGISTERS[11][8] ), .A2(n59), .B1(\REGISTERS[10][8] ), 
        .B2(n60), .ZN(n336) );
  OAI221_X1 U205 ( .B1(n61), .B2(n337), .C1(n63), .C2(n338), .A(n339), .ZN(
        n324) );
  AOI22_X1 U206 ( .A1(\REGISTERS[15][8] ), .A2(n66), .B1(\REGISTERS[14][8] ), 
        .B2(n67), .ZN(n339) );
  NAND2_X1 U207 ( .A1(n340), .A2(n341), .ZN(N4366) );
  NOR4_X1 U208 ( .A1(n342), .A2(n343), .A3(n344), .A4(n345), .ZN(n341) );
  OAI221_X1 U209 ( .B1(n8), .B2(n346), .C1(n10), .C2(n347), .A(n348), .ZN(n345) );
  AOI22_X1 U210 ( .A1(\REGISTERS[19][9] ), .A2(n13), .B1(\REGISTERS[18][9] ), 
        .B2(n14), .ZN(n348) );
  OAI221_X1 U211 ( .B1(n15), .B2(n349), .C1(n17), .C2(n350), .A(n351), .ZN(
        n344) );
  AOI22_X1 U212 ( .A1(\REGISTERS[23][9] ), .A2(n20), .B1(\REGISTERS[22][9] ), 
        .B2(n21), .ZN(n351) );
  OAI221_X1 U213 ( .B1(n22), .B2(n352), .C1(n24), .C2(n353), .A(n354), .ZN(
        n343) );
  AOI22_X1 U214 ( .A1(\REGISTERS[27][9] ), .A2(n27), .B1(\REGISTERS[26][9] ), 
        .B2(n28), .ZN(n354) );
  OAI221_X1 U215 ( .B1(n29), .B2(n355), .C1(n31), .C2(n356), .A(n357), .ZN(
        n342) );
  AOI22_X1 U216 ( .A1(\REGISTERS[29][9] ), .A2(n34), .B1(\REGISTERS[28][9] ), 
        .B2(n35), .ZN(n357) );
  NOR4_X1 U217 ( .A1(n358), .A2(n359), .A3(n360), .A4(n361), .ZN(n340) );
  AOI22_X1 U219 ( .A1(\REGISTERS[3][9] ), .A2(n45), .B1(\REGISTERS[2][9] ), 
        .B2(n46), .ZN(n364) );
  OAI221_X1 U220 ( .B1(n47), .B2(n365), .C1(n49), .C2(n366), .A(n367), .ZN(
        n360) );
  AOI22_X1 U221 ( .A1(\REGISTERS[7][9] ), .A2(n52), .B1(\REGISTERS[6][9] ), 
        .B2(n53), .ZN(n367) );
  OAI221_X1 U222 ( .B1(n54), .B2(n368), .C1(n56), .C2(n369), .A(n370), .ZN(
        n359) );
  AOI22_X1 U223 ( .A1(\REGISTERS[11][9] ), .A2(n59), .B1(\REGISTERS[10][9] ), 
        .B2(n60), .ZN(n370) );
  OAI221_X1 U224 ( .B1(n61), .B2(n371), .C1(n63), .C2(n372), .A(n373), .ZN(
        n358) );
  AOI22_X1 U225 ( .A1(\REGISTERS[15][9] ), .A2(n66), .B1(\REGISTERS[14][9] ), 
        .B2(n67), .ZN(n373) );
  NAND2_X1 U226 ( .A1(n374), .A2(n375), .ZN(N4365) );
  NOR4_X1 U227 ( .A1(n376), .A2(n377), .A3(n378), .A4(n379), .ZN(n375) );
  OAI221_X1 U228 ( .B1(n8), .B2(n380), .C1(n10), .C2(n381), .A(n382), .ZN(n379) );
  AOI22_X1 U229 ( .A1(\REGISTERS[19][10] ), .A2(n13), .B1(\REGISTERS[18][10] ), 
        .B2(n14), .ZN(n382) );
  OAI221_X1 U230 ( .B1(n15), .B2(n383), .C1(n17), .C2(n384), .A(n385), .ZN(
        n378) );
  AOI22_X1 U231 ( .A1(\REGISTERS[23][10] ), .A2(n20), .B1(\REGISTERS[22][10] ), 
        .B2(n21), .ZN(n385) );
  OAI221_X1 U232 ( .B1(n22), .B2(n386), .C1(n24), .C2(n387), .A(n388), .ZN(
        n377) );
  AOI22_X1 U233 ( .A1(\REGISTERS[27][10] ), .A2(n27), .B1(\REGISTERS[26][10] ), 
        .B2(n28), .ZN(n388) );
  OAI221_X1 U234 ( .B1(n29), .B2(n389), .C1(n31), .C2(n390), .A(n391), .ZN(
        n376) );
  AOI22_X1 U235 ( .A1(\REGISTERS[29][10] ), .A2(n34), .B1(\REGISTERS[28][10] ), 
        .B2(n35), .ZN(n391) );
  NOR4_X1 U236 ( .A1(n392), .A2(n393), .A3(n394), .A4(n395), .ZN(n374) );
  AOI22_X1 U238 ( .A1(\REGISTERS[3][10] ), .A2(n45), .B1(\REGISTERS[2][10] ), 
        .B2(n46), .ZN(n398) );
  OAI221_X1 U239 ( .B1(n47), .B2(n399), .C1(n49), .C2(n400), .A(n401), .ZN(
        n394) );
  AOI22_X1 U240 ( .A1(\REGISTERS[7][10] ), .A2(n52), .B1(\REGISTERS[6][10] ), 
        .B2(n53), .ZN(n401) );
  OAI221_X1 U241 ( .B1(n54), .B2(n402), .C1(n56), .C2(n403), .A(n404), .ZN(
        n393) );
  AOI22_X1 U242 ( .A1(\REGISTERS[11][10] ), .A2(n59), .B1(\REGISTERS[10][10] ), 
        .B2(n60), .ZN(n404) );
  OAI221_X1 U243 ( .B1(n61), .B2(n405), .C1(n63), .C2(n406), .A(n407), .ZN(
        n392) );
  AOI22_X1 U244 ( .A1(\REGISTERS[15][10] ), .A2(n66), .B1(\REGISTERS[14][10] ), 
        .B2(n67), .ZN(n407) );
  NAND2_X1 U245 ( .A1(n408), .A2(n409), .ZN(N4364) );
  NOR4_X1 U246 ( .A1(n410), .A2(n411), .A3(n412), .A4(n413), .ZN(n409) );
  OAI221_X1 U247 ( .B1(n8), .B2(n414), .C1(n10), .C2(n415), .A(n416), .ZN(n413) );
  AOI22_X1 U248 ( .A1(\REGISTERS[19][11] ), .A2(n13), .B1(\REGISTERS[18][11] ), 
        .B2(n14), .ZN(n416) );
  OAI221_X1 U249 ( .B1(n15), .B2(n417), .C1(n17), .C2(n418), .A(n419), .ZN(
        n412) );
  AOI22_X1 U250 ( .A1(\REGISTERS[23][11] ), .A2(n20), .B1(\REGISTERS[22][11] ), 
        .B2(n21), .ZN(n419) );
  OAI221_X1 U251 ( .B1(n22), .B2(n420), .C1(n24), .C2(n421), .A(n422), .ZN(
        n411) );
  AOI22_X1 U252 ( .A1(\REGISTERS[27][11] ), .A2(n27), .B1(\REGISTERS[26][11] ), 
        .B2(n28), .ZN(n422) );
  OAI221_X1 U253 ( .B1(n29), .B2(n423), .C1(n31), .C2(n424), .A(n425), .ZN(
        n410) );
  AOI22_X1 U254 ( .A1(\REGISTERS[29][11] ), .A2(n34), .B1(\REGISTERS[28][11] ), 
        .B2(n35), .ZN(n425) );
  NOR4_X1 U255 ( .A1(n426), .A2(n427), .A3(n428), .A4(n429), .ZN(n408) );
  AOI22_X1 U257 ( .A1(\REGISTERS[3][11] ), .A2(n45), .B1(\REGISTERS[2][11] ), 
        .B2(n46), .ZN(n432) );
  OAI221_X1 U258 ( .B1(n47), .B2(n433), .C1(n49), .C2(n434), .A(n435), .ZN(
        n428) );
  AOI22_X1 U259 ( .A1(\REGISTERS[7][11] ), .A2(n52), .B1(\REGISTERS[6][11] ), 
        .B2(n53), .ZN(n435) );
  OAI221_X1 U260 ( .B1(n54), .B2(n436), .C1(n56), .C2(n437), .A(n438), .ZN(
        n427) );
  AOI22_X1 U261 ( .A1(\REGISTERS[11][11] ), .A2(n59), .B1(\REGISTERS[10][11] ), 
        .B2(n60), .ZN(n438) );
  OAI221_X1 U262 ( .B1(n61), .B2(n439), .C1(n63), .C2(n440), .A(n441), .ZN(
        n426) );
  AOI22_X1 U263 ( .A1(\REGISTERS[15][11] ), .A2(n66), .B1(\REGISTERS[14][11] ), 
        .B2(n67), .ZN(n441) );
  NAND2_X1 U264 ( .A1(n442), .A2(n443), .ZN(N4363) );
  NOR4_X1 U265 ( .A1(n444), .A2(n445), .A3(n446), .A4(n447), .ZN(n443) );
  OAI221_X1 U266 ( .B1(n8), .B2(n448), .C1(n10), .C2(n449), .A(n450), .ZN(n447) );
  AOI22_X1 U267 ( .A1(\REGISTERS[19][12] ), .A2(n13), .B1(\REGISTERS[18][12] ), 
        .B2(n14), .ZN(n450) );
  OAI221_X1 U268 ( .B1(n15), .B2(n451), .C1(n17), .C2(n452), .A(n453), .ZN(
        n446) );
  AOI22_X1 U269 ( .A1(\REGISTERS[23][12] ), .A2(n20), .B1(\REGISTERS[22][12] ), 
        .B2(n21), .ZN(n453) );
  OAI221_X1 U270 ( .B1(n22), .B2(n454), .C1(n24), .C2(n455), .A(n456), .ZN(
        n445) );
  AOI22_X1 U271 ( .A1(\REGISTERS[27][12] ), .A2(n27), .B1(\REGISTERS[26][12] ), 
        .B2(n28), .ZN(n456) );
  OAI221_X1 U272 ( .B1(n29), .B2(n457), .C1(n31), .C2(n458), .A(n459), .ZN(
        n444) );
  AOI22_X1 U273 ( .A1(\REGISTERS[29][12] ), .A2(n34), .B1(\REGISTERS[28][12] ), 
        .B2(n35), .ZN(n459) );
  NOR4_X1 U274 ( .A1(n460), .A2(n461), .A3(n462), .A4(n463), .ZN(n442) );
  AOI22_X1 U276 ( .A1(\REGISTERS[3][12] ), .A2(n45), .B1(\REGISTERS[2][12] ), 
        .B2(n46), .ZN(n466) );
  OAI221_X1 U277 ( .B1(n47), .B2(n467), .C1(n49), .C2(n468), .A(n469), .ZN(
        n462) );
  AOI22_X1 U278 ( .A1(\REGISTERS[7][12] ), .A2(n52), .B1(\REGISTERS[6][12] ), 
        .B2(n53), .ZN(n469) );
  OAI221_X1 U279 ( .B1(n54), .B2(n470), .C1(n56), .C2(n471), .A(n472), .ZN(
        n461) );
  AOI22_X1 U280 ( .A1(\REGISTERS[11][12] ), .A2(n59), .B1(\REGISTERS[10][12] ), 
        .B2(n60), .ZN(n472) );
  OAI221_X1 U281 ( .B1(n61), .B2(n473), .C1(n63), .C2(n474), .A(n475), .ZN(
        n460) );
  AOI22_X1 U282 ( .A1(\REGISTERS[15][12] ), .A2(n66), .B1(\REGISTERS[14][12] ), 
        .B2(n67), .ZN(n475) );
  NAND2_X1 U283 ( .A1(n476), .A2(n477), .ZN(N4362) );
  NOR4_X1 U284 ( .A1(n478), .A2(n479), .A3(n480), .A4(n481), .ZN(n477) );
  OAI221_X1 U285 ( .B1(n8), .B2(n482), .C1(n10), .C2(n483), .A(n484), .ZN(n481) );
  AOI22_X1 U286 ( .A1(\REGISTERS[19][13] ), .A2(n13), .B1(\REGISTERS[18][13] ), 
        .B2(n14), .ZN(n484) );
  OAI221_X1 U287 ( .B1(n15), .B2(n485), .C1(n17), .C2(n486), .A(n487), .ZN(
        n480) );
  AOI22_X1 U288 ( .A1(\REGISTERS[23][13] ), .A2(n20), .B1(\REGISTERS[22][13] ), 
        .B2(n21), .ZN(n487) );
  OAI221_X1 U289 ( .B1(n22), .B2(n488), .C1(n24), .C2(n489), .A(n490), .ZN(
        n479) );
  AOI22_X1 U290 ( .A1(\REGISTERS[27][13] ), .A2(n27), .B1(\REGISTERS[26][13] ), 
        .B2(n28), .ZN(n490) );
  OAI221_X1 U291 ( .B1(n29), .B2(n491), .C1(n31), .C2(n492), .A(n493), .ZN(
        n478) );
  AOI22_X1 U292 ( .A1(\REGISTERS[29][13] ), .A2(n34), .B1(\REGISTERS[28][13] ), 
        .B2(n35), .ZN(n493) );
  NOR4_X1 U293 ( .A1(n494), .A2(n495), .A3(n496), .A4(n497), .ZN(n476) );
  AOI22_X1 U295 ( .A1(\REGISTERS[3][13] ), .A2(n45), .B1(\REGISTERS[2][13] ), 
        .B2(n46), .ZN(n500) );
  OAI221_X1 U296 ( .B1(n47), .B2(n501), .C1(n49), .C2(n502), .A(n503), .ZN(
        n496) );
  AOI22_X1 U297 ( .A1(\REGISTERS[7][13] ), .A2(n52), .B1(\REGISTERS[6][13] ), 
        .B2(n53), .ZN(n503) );
  OAI221_X1 U298 ( .B1(n54), .B2(n504), .C1(n56), .C2(n505), .A(n506), .ZN(
        n495) );
  AOI22_X1 U299 ( .A1(\REGISTERS[11][13] ), .A2(n59), .B1(\REGISTERS[10][13] ), 
        .B2(n60), .ZN(n506) );
  OAI221_X1 U300 ( .B1(n61), .B2(n507), .C1(n63), .C2(n508), .A(n509), .ZN(
        n494) );
  AOI22_X1 U301 ( .A1(\REGISTERS[15][13] ), .A2(n66), .B1(\REGISTERS[14][13] ), 
        .B2(n67), .ZN(n509) );
  NAND2_X1 U302 ( .A1(n510), .A2(n511), .ZN(N4361) );
  NOR4_X1 U303 ( .A1(n512), .A2(n513), .A3(n514), .A4(n515), .ZN(n511) );
  OAI221_X1 U304 ( .B1(n8), .B2(n516), .C1(n10), .C2(n517), .A(n518), .ZN(n515) );
  AOI22_X1 U305 ( .A1(\REGISTERS[19][14] ), .A2(n13), .B1(\REGISTERS[18][14] ), 
        .B2(n14), .ZN(n518) );
  OAI221_X1 U306 ( .B1(n15), .B2(n519), .C1(n17), .C2(n520), .A(n521), .ZN(
        n514) );
  AOI22_X1 U307 ( .A1(\REGISTERS[23][14] ), .A2(n20), .B1(\REGISTERS[22][14] ), 
        .B2(n21), .ZN(n521) );
  OAI221_X1 U308 ( .B1(n22), .B2(n522), .C1(n24), .C2(n523), .A(n524), .ZN(
        n513) );
  AOI22_X1 U309 ( .A1(\REGISTERS[27][14] ), .A2(n27), .B1(\REGISTERS[26][14] ), 
        .B2(n28), .ZN(n524) );
  OAI221_X1 U310 ( .B1(n29), .B2(n525), .C1(n31), .C2(n526), .A(n527), .ZN(
        n512) );
  AOI22_X1 U311 ( .A1(\REGISTERS[29][14] ), .A2(n34), .B1(\REGISTERS[28][14] ), 
        .B2(n35), .ZN(n527) );
  NOR4_X1 U312 ( .A1(n528), .A2(n529), .A3(n530), .A4(n531), .ZN(n510) );
  AOI22_X1 U314 ( .A1(\REGISTERS[3][14] ), .A2(n45), .B1(\REGISTERS[2][14] ), 
        .B2(n46), .ZN(n534) );
  OAI221_X1 U315 ( .B1(n47), .B2(n535), .C1(n49), .C2(n536), .A(n537), .ZN(
        n530) );
  AOI22_X1 U316 ( .A1(\REGISTERS[7][14] ), .A2(n52), .B1(\REGISTERS[6][14] ), 
        .B2(n53), .ZN(n537) );
  OAI221_X1 U317 ( .B1(n54), .B2(n538), .C1(n56), .C2(n539), .A(n540), .ZN(
        n529) );
  AOI22_X1 U318 ( .A1(\REGISTERS[11][14] ), .A2(n59), .B1(\REGISTERS[10][14] ), 
        .B2(n60), .ZN(n540) );
  OAI221_X1 U319 ( .B1(n61), .B2(n541), .C1(n63), .C2(n542), .A(n543), .ZN(
        n528) );
  AOI22_X1 U320 ( .A1(\REGISTERS[15][14] ), .A2(n66), .B1(\REGISTERS[14][14] ), 
        .B2(n67), .ZN(n543) );
  NAND2_X1 U321 ( .A1(n544), .A2(n545), .ZN(N4360) );
  NOR4_X1 U322 ( .A1(n546), .A2(n547), .A3(n548), .A4(n549), .ZN(n545) );
  OAI221_X1 U323 ( .B1(n8), .B2(n550), .C1(n10), .C2(n551), .A(n552), .ZN(n549) );
  AOI22_X1 U324 ( .A1(\REGISTERS[19][15] ), .A2(n13), .B1(\REGISTERS[18][15] ), 
        .B2(n14), .ZN(n552) );
  OAI221_X1 U325 ( .B1(n15), .B2(n553), .C1(n17), .C2(n554), .A(n555), .ZN(
        n548) );
  AOI22_X1 U326 ( .A1(\REGISTERS[23][15] ), .A2(n20), .B1(\REGISTERS[22][15] ), 
        .B2(n21), .ZN(n555) );
  OAI221_X1 U327 ( .B1(n22), .B2(n556), .C1(n24), .C2(n557), .A(n558), .ZN(
        n547) );
  AOI22_X1 U328 ( .A1(\REGISTERS[27][15] ), .A2(n27), .B1(\REGISTERS[26][15] ), 
        .B2(n28), .ZN(n558) );
  OAI221_X1 U329 ( .B1(n29), .B2(n559), .C1(n31), .C2(n560), .A(n561), .ZN(
        n546) );
  AOI22_X1 U330 ( .A1(\REGISTERS[29][15] ), .A2(n34), .B1(\REGISTERS[28][15] ), 
        .B2(n35), .ZN(n561) );
  NOR4_X1 U331 ( .A1(n562), .A2(n563), .A3(n564), .A4(n565), .ZN(n544) );
  AOI22_X1 U333 ( .A1(\REGISTERS[3][15] ), .A2(n45), .B1(\REGISTERS[2][15] ), 
        .B2(n46), .ZN(n568) );
  OAI221_X1 U334 ( .B1(n47), .B2(n569), .C1(n49), .C2(n570), .A(n571), .ZN(
        n564) );
  AOI22_X1 U335 ( .A1(\REGISTERS[7][15] ), .A2(n52), .B1(\REGISTERS[6][15] ), 
        .B2(n53), .ZN(n571) );
  OAI221_X1 U336 ( .B1(n54), .B2(n572), .C1(n56), .C2(n573), .A(n574), .ZN(
        n563) );
  AOI22_X1 U337 ( .A1(\REGISTERS[11][15] ), .A2(n59), .B1(\REGISTERS[10][15] ), 
        .B2(n60), .ZN(n574) );
  OAI221_X1 U338 ( .B1(n61), .B2(n575), .C1(n63), .C2(n576), .A(n577), .ZN(
        n562) );
  AOI22_X1 U339 ( .A1(\REGISTERS[15][15] ), .A2(n66), .B1(\REGISTERS[14][15] ), 
        .B2(n67), .ZN(n577) );
  NAND2_X1 U340 ( .A1(n578), .A2(n579), .ZN(N4359) );
  NOR4_X1 U341 ( .A1(n580), .A2(n581), .A3(n582), .A4(n583), .ZN(n579) );
  OAI221_X1 U342 ( .B1(n8), .B2(n584), .C1(n10), .C2(n585), .A(n586), .ZN(n583) );
  AOI22_X1 U343 ( .A1(\REGISTERS[19][16] ), .A2(n13), .B1(\REGISTERS[18][16] ), 
        .B2(n14), .ZN(n586) );
  OAI221_X1 U344 ( .B1(n15), .B2(n587), .C1(n17), .C2(n588), .A(n589), .ZN(
        n582) );
  AOI22_X1 U345 ( .A1(\REGISTERS[23][16] ), .A2(n20), .B1(\REGISTERS[22][16] ), 
        .B2(n21), .ZN(n589) );
  OAI221_X1 U346 ( .B1(n22), .B2(n590), .C1(n24), .C2(n591), .A(n592), .ZN(
        n581) );
  AOI22_X1 U347 ( .A1(\REGISTERS[27][16] ), .A2(n27), .B1(\REGISTERS[26][16] ), 
        .B2(n28), .ZN(n592) );
  OAI221_X1 U348 ( .B1(n29), .B2(n593), .C1(n31), .C2(n594), .A(n595), .ZN(
        n580) );
  AOI22_X1 U349 ( .A1(\REGISTERS[29][16] ), .A2(n34), .B1(\REGISTERS[28][16] ), 
        .B2(n35), .ZN(n595) );
  NOR4_X1 U350 ( .A1(n596), .A2(n597), .A3(n598), .A4(n599), .ZN(n578) );
  AOI22_X1 U352 ( .A1(\REGISTERS[3][16] ), .A2(n45), .B1(\REGISTERS[2][16] ), 
        .B2(n46), .ZN(n602) );
  OAI221_X1 U353 ( .B1(n47), .B2(n603), .C1(n49), .C2(n604), .A(n605), .ZN(
        n598) );
  AOI22_X1 U354 ( .A1(\REGISTERS[7][16] ), .A2(n52), .B1(\REGISTERS[6][16] ), 
        .B2(n53), .ZN(n605) );
  OAI221_X1 U355 ( .B1(n54), .B2(n606), .C1(n56), .C2(n607), .A(n608), .ZN(
        n597) );
  AOI22_X1 U356 ( .A1(\REGISTERS[11][16] ), .A2(n59), .B1(\REGISTERS[10][16] ), 
        .B2(n60), .ZN(n608) );
  OAI221_X1 U357 ( .B1(n61), .B2(n609), .C1(n63), .C2(n610), .A(n611), .ZN(
        n596) );
  AOI22_X1 U358 ( .A1(\REGISTERS[15][16] ), .A2(n66), .B1(\REGISTERS[14][16] ), 
        .B2(n67), .ZN(n611) );
  NAND2_X1 U359 ( .A1(n612), .A2(n613), .ZN(N4358) );
  NOR4_X1 U360 ( .A1(n614), .A2(n615), .A3(n616), .A4(n617), .ZN(n613) );
  OAI221_X1 U361 ( .B1(n8), .B2(n618), .C1(n10), .C2(n619), .A(n620), .ZN(n617) );
  AOI22_X1 U362 ( .A1(\REGISTERS[19][17] ), .A2(n13), .B1(\REGISTERS[18][17] ), 
        .B2(n14), .ZN(n620) );
  OAI221_X1 U363 ( .B1(n15), .B2(n621), .C1(n17), .C2(n622), .A(n623), .ZN(
        n616) );
  AOI22_X1 U364 ( .A1(\REGISTERS[23][17] ), .A2(n20), .B1(\REGISTERS[22][17] ), 
        .B2(n21), .ZN(n623) );
  OAI221_X1 U365 ( .B1(n22), .B2(n624), .C1(n24), .C2(n625), .A(n626), .ZN(
        n615) );
  AOI22_X1 U366 ( .A1(\REGISTERS[27][17] ), .A2(n27), .B1(\REGISTERS[26][17] ), 
        .B2(n28), .ZN(n626) );
  OAI221_X1 U367 ( .B1(n29), .B2(n627), .C1(n31), .C2(n628), .A(n629), .ZN(
        n614) );
  AOI22_X1 U368 ( .A1(\REGISTERS[29][17] ), .A2(n34), .B1(\REGISTERS[28][17] ), 
        .B2(n35), .ZN(n629) );
  NOR4_X1 U369 ( .A1(n630), .A2(n631), .A3(n632), .A4(n633), .ZN(n612) );
  AOI22_X1 U371 ( .A1(\REGISTERS[3][17] ), .A2(n45), .B1(\REGISTERS[2][17] ), 
        .B2(n46), .ZN(n636) );
  OAI221_X1 U372 ( .B1(n47), .B2(n637), .C1(n49), .C2(n638), .A(n639), .ZN(
        n632) );
  AOI22_X1 U373 ( .A1(\REGISTERS[7][17] ), .A2(n52), .B1(\REGISTERS[6][17] ), 
        .B2(n53), .ZN(n639) );
  OAI221_X1 U374 ( .B1(n54), .B2(n640), .C1(n56), .C2(n641), .A(n642), .ZN(
        n631) );
  AOI22_X1 U375 ( .A1(\REGISTERS[11][17] ), .A2(n59), .B1(\REGISTERS[10][17] ), 
        .B2(n60), .ZN(n642) );
  OAI221_X1 U376 ( .B1(n61), .B2(n643), .C1(n63), .C2(n644), .A(n645), .ZN(
        n630) );
  AOI22_X1 U377 ( .A1(\REGISTERS[15][17] ), .A2(n66), .B1(\REGISTERS[14][17] ), 
        .B2(n67), .ZN(n645) );
  NAND2_X1 U378 ( .A1(n646), .A2(n647), .ZN(N4357) );
  NOR4_X1 U379 ( .A1(n648), .A2(n649), .A3(n650), .A4(n651), .ZN(n647) );
  OAI221_X1 U380 ( .B1(n8), .B2(n652), .C1(n10), .C2(n653), .A(n654), .ZN(n651) );
  AOI22_X1 U381 ( .A1(\REGISTERS[19][18] ), .A2(n13), .B1(\REGISTERS[18][18] ), 
        .B2(n14), .ZN(n654) );
  OAI221_X1 U382 ( .B1(n15), .B2(n655), .C1(n17), .C2(n656), .A(n657), .ZN(
        n650) );
  AOI22_X1 U383 ( .A1(\REGISTERS[23][18] ), .A2(n20), .B1(\REGISTERS[22][18] ), 
        .B2(n21), .ZN(n657) );
  OAI221_X1 U384 ( .B1(n22), .B2(n658), .C1(n24), .C2(n659), .A(n660), .ZN(
        n649) );
  AOI22_X1 U385 ( .A1(\REGISTERS[27][18] ), .A2(n27), .B1(\REGISTERS[26][18] ), 
        .B2(n28), .ZN(n660) );
  OAI221_X1 U386 ( .B1(n29), .B2(n661), .C1(n31), .C2(n662), .A(n663), .ZN(
        n648) );
  AOI22_X1 U387 ( .A1(\REGISTERS[29][18] ), .A2(n34), .B1(\REGISTERS[28][18] ), 
        .B2(n35), .ZN(n663) );
  NOR4_X1 U388 ( .A1(n664), .A2(n665), .A3(n666), .A4(n667), .ZN(n646) );
  AOI22_X1 U390 ( .A1(\REGISTERS[3][18] ), .A2(n45), .B1(\REGISTERS[2][18] ), 
        .B2(n46), .ZN(n670) );
  OAI221_X1 U391 ( .B1(n47), .B2(n671), .C1(n49), .C2(n672), .A(n673), .ZN(
        n666) );
  AOI22_X1 U392 ( .A1(\REGISTERS[7][18] ), .A2(n52), .B1(\REGISTERS[6][18] ), 
        .B2(n53), .ZN(n673) );
  OAI221_X1 U393 ( .B1(n54), .B2(n674), .C1(n56), .C2(n675), .A(n676), .ZN(
        n665) );
  AOI22_X1 U394 ( .A1(\REGISTERS[11][18] ), .A2(n59), .B1(\REGISTERS[10][18] ), 
        .B2(n60), .ZN(n676) );
  OAI221_X1 U395 ( .B1(n61), .B2(n677), .C1(n63), .C2(n678), .A(n679), .ZN(
        n664) );
  AOI22_X1 U396 ( .A1(\REGISTERS[15][18] ), .A2(n66), .B1(\REGISTERS[14][18] ), 
        .B2(n67), .ZN(n679) );
  NAND2_X1 U397 ( .A1(n680), .A2(n681), .ZN(N4356) );
  NOR4_X1 U398 ( .A1(n682), .A2(n683), .A3(n684), .A4(n685), .ZN(n681) );
  OAI221_X1 U399 ( .B1(n8), .B2(n686), .C1(n10), .C2(n687), .A(n688), .ZN(n685) );
  AOI22_X1 U400 ( .A1(\REGISTERS[19][19] ), .A2(n13), .B1(\REGISTERS[18][19] ), 
        .B2(n14), .ZN(n688) );
  OAI221_X1 U401 ( .B1(n15), .B2(n689), .C1(n17), .C2(n690), .A(n691), .ZN(
        n684) );
  AOI22_X1 U402 ( .A1(\REGISTERS[23][19] ), .A2(n20), .B1(\REGISTERS[22][19] ), 
        .B2(n21), .ZN(n691) );
  OAI221_X1 U403 ( .B1(n22), .B2(n692), .C1(n24), .C2(n693), .A(n694), .ZN(
        n683) );
  AOI22_X1 U404 ( .A1(\REGISTERS[27][19] ), .A2(n27), .B1(\REGISTERS[26][19] ), 
        .B2(n28), .ZN(n694) );
  OAI221_X1 U405 ( .B1(n29), .B2(n695), .C1(n31), .C2(n696), .A(n697), .ZN(
        n682) );
  AOI22_X1 U406 ( .A1(\REGISTERS[29][19] ), .A2(n34), .B1(\REGISTERS[28][19] ), 
        .B2(n35), .ZN(n697) );
  NOR4_X1 U407 ( .A1(n698), .A2(n699), .A3(n700), .A4(n701), .ZN(n680) );
  AOI22_X1 U409 ( .A1(\REGISTERS[3][19] ), .A2(n45), .B1(\REGISTERS[2][19] ), 
        .B2(n46), .ZN(n704) );
  OAI221_X1 U410 ( .B1(n47), .B2(n705), .C1(n49), .C2(n706), .A(n707), .ZN(
        n700) );
  AOI22_X1 U411 ( .A1(\REGISTERS[7][19] ), .A2(n52), .B1(\REGISTERS[6][19] ), 
        .B2(n53), .ZN(n707) );
  OAI221_X1 U412 ( .B1(n54), .B2(n708), .C1(n56), .C2(n709), .A(n710), .ZN(
        n699) );
  AOI22_X1 U413 ( .A1(\REGISTERS[11][19] ), .A2(n59), .B1(\REGISTERS[10][19] ), 
        .B2(n60), .ZN(n710) );
  OAI221_X1 U414 ( .B1(n61), .B2(n711), .C1(n63), .C2(n712), .A(n713), .ZN(
        n698) );
  AOI22_X1 U415 ( .A1(\REGISTERS[15][19] ), .A2(n66), .B1(\REGISTERS[14][19] ), 
        .B2(n67), .ZN(n713) );
  NAND2_X1 U416 ( .A1(n714), .A2(n715), .ZN(N4355) );
  NOR4_X1 U417 ( .A1(n716), .A2(n717), .A3(n718), .A4(n719), .ZN(n715) );
  OAI221_X1 U418 ( .B1(n8), .B2(n720), .C1(n10), .C2(n721), .A(n722), .ZN(n719) );
  AOI22_X1 U419 ( .A1(\REGISTERS[19][20] ), .A2(n13), .B1(\REGISTERS[18][20] ), 
        .B2(n14), .ZN(n722) );
  OAI221_X1 U420 ( .B1(n15), .B2(n723), .C1(n17), .C2(n724), .A(n725), .ZN(
        n718) );
  AOI22_X1 U421 ( .A1(\REGISTERS[23][20] ), .A2(n20), .B1(\REGISTERS[22][20] ), 
        .B2(n21), .ZN(n725) );
  OAI221_X1 U422 ( .B1(n22), .B2(n726), .C1(n24), .C2(n727), .A(n728), .ZN(
        n717) );
  AOI22_X1 U423 ( .A1(\REGISTERS[27][20] ), .A2(n27), .B1(\REGISTERS[26][20] ), 
        .B2(n28), .ZN(n728) );
  OAI221_X1 U424 ( .B1(n29), .B2(n729), .C1(n31), .C2(n730), .A(n731), .ZN(
        n716) );
  AOI22_X1 U425 ( .A1(\REGISTERS[29][20] ), .A2(n34), .B1(\REGISTERS[28][20] ), 
        .B2(n35), .ZN(n731) );
  NOR4_X1 U426 ( .A1(n732), .A2(n733), .A3(n734), .A4(n735), .ZN(n714) );
  AOI22_X1 U428 ( .A1(\REGISTERS[3][20] ), .A2(n45), .B1(\REGISTERS[2][20] ), 
        .B2(n46), .ZN(n738) );
  OAI221_X1 U429 ( .B1(n47), .B2(n739), .C1(n49), .C2(n740), .A(n741), .ZN(
        n734) );
  AOI22_X1 U430 ( .A1(\REGISTERS[7][20] ), .A2(n52), .B1(\REGISTERS[6][20] ), 
        .B2(n53), .ZN(n741) );
  OAI221_X1 U431 ( .B1(n54), .B2(n742), .C1(n56), .C2(n743), .A(n744), .ZN(
        n733) );
  AOI22_X1 U432 ( .A1(\REGISTERS[11][20] ), .A2(n59), .B1(\REGISTERS[10][20] ), 
        .B2(n60), .ZN(n744) );
  OAI221_X1 U433 ( .B1(n61), .B2(n745), .C1(n63), .C2(n746), .A(n747), .ZN(
        n732) );
  AOI22_X1 U434 ( .A1(\REGISTERS[15][20] ), .A2(n66), .B1(\REGISTERS[14][20] ), 
        .B2(n67), .ZN(n747) );
  NAND2_X1 U435 ( .A1(n748), .A2(n749), .ZN(N4354) );
  NOR4_X1 U436 ( .A1(n750), .A2(n751), .A3(n752), .A4(n753), .ZN(n749) );
  OAI221_X1 U437 ( .B1(n8), .B2(n754), .C1(n10), .C2(n755), .A(n756), .ZN(n753) );
  AOI22_X1 U438 ( .A1(\REGISTERS[19][21] ), .A2(n13), .B1(\REGISTERS[18][21] ), 
        .B2(n14), .ZN(n756) );
  OAI221_X1 U439 ( .B1(n15), .B2(n757), .C1(n17), .C2(n758), .A(n759), .ZN(
        n752) );
  AOI22_X1 U440 ( .A1(\REGISTERS[23][21] ), .A2(n20), .B1(\REGISTERS[22][21] ), 
        .B2(n21), .ZN(n759) );
  OAI221_X1 U441 ( .B1(n22), .B2(n760), .C1(n24), .C2(n761), .A(n762), .ZN(
        n751) );
  AOI22_X1 U442 ( .A1(\REGISTERS[27][21] ), .A2(n27), .B1(\REGISTERS[26][21] ), 
        .B2(n28), .ZN(n762) );
  OAI221_X1 U443 ( .B1(n29), .B2(n763), .C1(n31), .C2(n764), .A(n765), .ZN(
        n750) );
  AOI22_X1 U444 ( .A1(\REGISTERS[29][21] ), .A2(n34), .B1(\REGISTERS[28][21] ), 
        .B2(n35), .ZN(n765) );
  NOR4_X1 U445 ( .A1(n766), .A2(n767), .A3(n768), .A4(n769), .ZN(n748) );
  AOI22_X1 U447 ( .A1(\REGISTERS[3][21] ), .A2(n45), .B1(\REGISTERS[2][21] ), 
        .B2(n46), .ZN(n772) );
  OAI221_X1 U448 ( .B1(n47), .B2(n773), .C1(n49), .C2(n774), .A(n775), .ZN(
        n768) );
  AOI22_X1 U449 ( .A1(\REGISTERS[7][21] ), .A2(n52), .B1(\REGISTERS[6][21] ), 
        .B2(n53), .ZN(n775) );
  OAI221_X1 U450 ( .B1(n54), .B2(n776), .C1(n56), .C2(n777), .A(n778), .ZN(
        n767) );
  AOI22_X1 U451 ( .A1(\REGISTERS[11][21] ), .A2(n59), .B1(\REGISTERS[10][21] ), 
        .B2(n60), .ZN(n778) );
  OAI221_X1 U452 ( .B1(n61), .B2(n779), .C1(n63), .C2(n780), .A(n781), .ZN(
        n766) );
  AOI22_X1 U453 ( .A1(\REGISTERS[15][21] ), .A2(n66), .B1(\REGISTERS[14][21] ), 
        .B2(n67), .ZN(n781) );
  NAND2_X1 U454 ( .A1(n782), .A2(n783), .ZN(N4353) );
  NOR4_X1 U455 ( .A1(n784), .A2(n785), .A3(n786), .A4(n787), .ZN(n783) );
  OAI221_X1 U456 ( .B1(n8), .B2(n788), .C1(n10), .C2(n789), .A(n790), .ZN(n787) );
  AOI22_X1 U457 ( .A1(\REGISTERS[19][22] ), .A2(n13), .B1(\REGISTERS[18][22] ), 
        .B2(n14), .ZN(n790) );
  OAI221_X1 U458 ( .B1(n15), .B2(n791), .C1(n17), .C2(n792), .A(n793), .ZN(
        n786) );
  AOI22_X1 U459 ( .A1(\REGISTERS[23][22] ), .A2(n20), .B1(\REGISTERS[22][22] ), 
        .B2(n21), .ZN(n793) );
  OAI221_X1 U460 ( .B1(n22), .B2(n794), .C1(n24), .C2(n795), .A(n796), .ZN(
        n785) );
  AOI22_X1 U461 ( .A1(\REGISTERS[27][22] ), .A2(n27), .B1(\REGISTERS[26][22] ), 
        .B2(n28), .ZN(n796) );
  OAI221_X1 U462 ( .B1(n29), .B2(n797), .C1(n31), .C2(n798), .A(n799), .ZN(
        n784) );
  AOI22_X1 U463 ( .A1(\REGISTERS[29][22] ), .A2(n34), .B1(\REGISTERS[28][22] ), 
        .B2(n35), .ZN(n799) );
  NOR4_X1 U464 ( .A1(n800), .A2(n801), .A3(n802), .A4(n803), .ZN(n782) );
  AOI22_X1 U466 ( .A1(\REGISTERS[3][22] ), .A2(n45), .B1(\REGISTERS[2][22] ), 
        .B2(n46), .ZN(n806) );
  OAI221_X1 U467 ( .B1(n47), .B2(n807), .C1(n49), .C2(n808), .A(n809), .ZN(
        n802) );
  AOI22_X1 U468 ( .A1(\REGISTERS[7][22] ), .A2(n52), .B1(\REGISTERS[6][22] ), 
        .B2(n53), .ZN(n809) );
  OAI221_X1 U469 ( .B1(n54), .B2(n810), .C1(n56), .C2(n811), .A(n812), .ZN(
        n801) );
  AOI22_X1 U470 ( .A1(\REGISTERS[11][22] ), .A2(n59), .B1(\REGISTERS[10][22] ), 
        .B2(n60), .ZN(n812) );
  OAI221_X1 U471 ( .B1(n61), .B2(n813), .C1(n63), .C2(n814), .A(n815), .ZN(
        n800) );
  AOI22_X1 U472 ( .A1(\REGISTERS[15][22] ), .A2(n66), .B1(\REGISTERS[14][22] ), 
        .B2(n67), .ZN(n815) );
  NAND2_X1 U473 ( .A1(n816), .A2(n817), .ZN(N4352) );
  NOR4_X1 U474 ( .A1(n818), .A2(n819), .A3(n820), .A4(n821), .ZN(n817) );
  OAI221_X1 U475 ( .B1(n8), .B2(n822), .C1(n10), .C2(n823), .A(n824), .ZN(n821) );
  AOI22_X1 U476 ( .A1(\REGISTERS[19][23] ), .A2(n13), .B1(\REGISTERS[18][23] ), 
        .B2(n14), .ZN(n824) );
  OAI221_X1 U477 ( .B1(n15), .B2(n825), .C1(n17), .C2(n826), .A(n827), .ZN(
        n820) );
  AOI22_X1 U478 ( .A1(\REGISTERS[23][23] ), .A2(n20), .B1(\REGISTERS[22][23] ), 
        .B2(n21), .ZN(n827) );
  OAI221_X1 U479 ( .B1(n22), .B2(n828), .C1(n24), .C2(n829), .A(n830), .ZN(
        n819) );
  AOI22_X1 U480 ( .A1(\REGISTERS[27][23] ), .A2(n27), .B1(\REGISTERS[26][23] ), 
        .B2(n28), .ZN(n830) );
  OAI221_X1 U481 ( .B1(n29), .B2(n831), .C1(n31), .C2(n832), .A(n833), .ZN(
        n818) );
  AOI22_X1 U482 ( .A1(\REGISTERS[29][23] ), .A2(n34), .B1(\REGISTERS[28][23] ), 
        .B2(n35), .ZN(n833) );
  NOR4_X1 U483 ( .A1(n834), .A2(n835), .A3(n836), .A4(n837), .ZN(n816) );
  AOI22_X1 U485 ( .A1(\REGISTERS[3][23] ), .A2(n45), .B1(\REGISTERS[2][23] ), 
        .B2(n46), .ZN(n840) );
  OAI221_X1 U486 ( .B1(n47), .B2(n841), .C1(n49), .C2(n842), .A(n843), .ZN(
        n836) );
  AOI22_X1 U487 ( .A1(\REGISTERS[7][23] ), .A2(n52), .B1(\REGISTERS[6][23] ), 
        .B2(n53), .ZN(n843) );
  OAI221_X1 U488 ( .B1(n54), .B2(n844), .C1(n56), .C2(n845), .A(n846), .ZN(
        n835) );
  AOI22_X1 U489 ( .A1(\REGISTERS[11][23] ), .A2(n59), .B1(\REGISTERS[10][23] ), 
        .B2(n60), .ZN(n846) );
  OAI221_X1 U490 ( .B1(n61), .B2(n847), .C1(n63), .C2(n848), .A(n849), .ZN(
        n834) );
  AOI22_X1 U491 ( .A1(\REGISTERS[15][23] ), .A2(n66), .B1(\REGISTERS[14][23] ), 
        .B2(n67), .ZN(n849) );
  NAND2_X1 U492 ( .A1(n850), .A2(n851), .ZN(N4351) );
  NOR4_X1 U493 ( .A1(n852), .A2(n853), .A3(n854), .A4(n855), .ZN(n851) );
  OAI221_X1 U494 ( .B1(n8), .B2(n856), .C1(n10), .C2(n857), .A(n858), .ZN(n855) );
  AOI22_X1 U495 ( .A1(\REGISTERS[19][24] ), .A2(n13), .B1(\REGISTERS[18][24] ), 
        .B2(n14), .ZN(n858) );
  OAI221_X1 U496 ( .B1(n15), .B2(n859), .C1(n17), .C2(n860), .A(n861), .ZN(
        n854) );
  AOI22_X1 U497 ( .A1(\REGISTERS[23][24] ), .A2(n20), .B1(\REGISTERS[22][24] ), 
        .B2(n21), .ZN(n861) );
  OAI221_X1 U498 ( .B1(n22), .B2(n862), .C1(n24), .C2(n863), .A(n864), .ZN(
        n853) );
  AOI22_X1 U499 ( .A1(\REGISTERS[27][24] ), .A2(n27), .B1(\REGISTERS[26][24] ), 
        .B2(n28), .ZN(n864) );
  OAI221_X1 U500 ( .B1(n29), .B2(n865), .C1(n31), .C2(n866), .A(n867), .ZN(
        n852) );
  AOI22_X1 U501 ( .A1(\REGISTERS[29][24] ), .A2(n34), .B1(\REGISTERS[28][24] ), 
        .B2(n35), .ZN(n867) );
  NOR4_X1 U502 ( .A1(n868), .A2(n869), .A3(n870), .A4(n871), .ZN(n850) );
  AOI22_X1 U504 ( .A1(\REGISTERS[3][24] ), .A2(n45), .B1(\REGISTERS[2][24] ), 
        .B2(n46), .ZN(n874) );
  OAI221_X1 U505 ( .B1(n47), .B2(n875), .C1(n49), .C2(n876), .A(n877), .ZN(
        n870) );
  AOI22_X1 U506 ( .A1(\REGISTERS[7][24] ), .A2(n52), .B1(\REGISTERS[6][24] ), 
        .B2(n53), .ZN(n877) );
  OAI221_X1 U507 ( .B1(n54), .B2(n878), .C1(n56), .C2(n879), .A(n880), .ZN(
        n869) );
  AOI22_X1 U508 ( .A1(\REGISTERS[11][24] ), .A2(n59), .B1(\REGISTERS[10][24] ), 
        .B2(n60), .ZN(n880) );
  OAI221_X1 U509 ( .B1(n61), .B2(n881), .C1(n63), .C2(n882), .A(n883), .ZN(
        n868) );
  AOI22_X1 U510 ( .A1(\REGISTERS[15][24] ), .A2(n66), .B1(\REGISTERS[14][24] ), 
        .B2(n67), .ZN(n883) );
  NAND2_X1 U511 ( .A1(n884), .A2(n885), .ZN(N4350) );
  NOR4_X1 U512 ( .A1(n886), .A2(n887), .A3(n888), .A4(n889), .ZN(n885) );
  OAI221_X1 U513 ( .B1(n8), .B2(n890), .C1(n10), .C2(n891), .A(n892), .ZN(n889) );
  AOI22_X1 U514 ( .A1(\REGISTERS[19][25] ), .A2(n13), .B1(\REGISTERS[18][25] ), 
        .B2(n14), .ZN(n892) );
  OAI221_X1 U515 ( .B1(n15), .B2(n893), .C1(n17), .C2(n894), .A(n895), .ZN(
        n888) );
  AOI22_X1 U516 ( .A1(\REGISTERS[23][25] ), .A2(n20), .B1(\REGISTERS[22][25] ), 
        .B2(n21), .ZN(n895) );
  OAI221_X1 U517 ( .B1(n22), .B2(n896), .C1(n24), .C2(n897), .A(n898), .ZN(
        n887) );
  AOI22_X1 U518 ( .A1(\REGISTERS[27][25] ), .A2(n27), .B1(\REGISTERS[26][25] ), 
        .B2(n28), .ZN(n898) );
  OAI221_X1 U519 ( .B1(n29), .B2(n899), .C1(n31), .C2(n900), .A(n901), .ZN(
        n886) );
  AOI22_X1 U520 ( .A1(\REGISTERS[29][25] ), .A2(n34), .B1(\REGISTERS[28][25] ), 
        .B2(n35), .ZN(n901) );
  NOR4_X1 U521 ( .A1(n902), .A2(n903), .A3(n904), .A4(n905), .ZN(n884) );
  AOI22_X1 U523 ( .A1(\REGISTERS[3][25] ), .A2(n45), .B1(\REGISTERS[2][25] ), 
        .B2(n46), .ZN(n908) );
  OAI221_X1 U524 ( .B1(n47), .B2(n909), .C1(n49), .C2(n910), .A(n911), .ZN(
        n904) );
  AOI22_X1 U525 ( .A1(\REGISTERS[7][25] ), .A2(n52), .B1(\REGISTERS[6][25] ), 
        .B2(n53), .ZN(n911) );
  OAI221_X1 U526 ( .B1(n54), .B2(n912), .C1(n56), .C2(n913), .A(n914), .ZN(
        n903) );
  AOI22_X1 U527 ( .A1(\REGISTERS[11][25] ), .A2(n59), .B1(\REGISTERS[10][25] ), 
        .B2(n60), .ZN(n914) );
  OAI221_X1 U528 ( .B1(n61), .B2(n915), .C1(n63), .C2(n916), .A(n917), .ZN(
        n902) );
  AOI22_X1 U529 ( .A1(\REGISTERS[15][25] ), .A2(n66), .B1(\REGISTERS[14][25] ), 
        .B2(n67), .ZN(n917) );
  NAND2_X1 U530 ( .A1(n918), .A2(n919), .ZN(N4349) );
  NOR4_X1 U531 ( .A1(n920), .A2(n921), .A3(n922), .A4(n923), .ZN(n919) );
  OAI221_X1 U532 ( .B1(n8), .B2(n924), .C1(n10), .C2(n925), .A(n926), .ZN(n923) );
  AOI22_X1 U533 ( .A1(\REGISTERS[19][26] ), .A2(n13), .B1(\REGISTERS[18][26] ), 
        .B2(n14), .ZN(n926) );
  OAI221_X1 U534 ( .B1(n15), .B2(n927), .C1(n17), .C2(n928), .A(n929), .ZN(
        n922) );
  AOI22_X1 U535 ( .A1(\REGISTERS[23][26] ), .A2(n20), .B1(\REGISTERS[22][26] ), 
        .B2(n21), .ZN(n929) );
  OAI221_X1 U536 ( .B1(n22), .B2(n930), .C1(n24), .C2(n931), .A(n932), .ZN(
        n921) );
  AOI22_X1 U537 ( .A1(\REGISTERS[27][26] ), .A2(n27), .B1(\REGISTERS[26][26] ), 
        .B2(n28), .ZN(n932) );
  OAI221_X1 U538 ( .B1(n29), .B2(n933), .C1(n31), .C2(n934), .A(n935), .ZN(
        n920) );
  AOI22_X1 U539 ( .A1(\REGISTERS[29][26] ), .A2(n34), .B1(\REGISTERS[28][26] ), 
        .B2(n35), .ZN(n935) );
  NOR4_X1 U540 ( .A1(n936), .A2(n937), .A3(n938), .A4(n939), .ZN(n918) );
  AOI22_X1 U542 ( .A1(\REGISTERS[3][26] ), .A2(n45), .B1(\REGISTERS[2][26] ), 
        .B2(n46), .ZN(n942) );
  OAI221_X1 U543 ( .B1(n47), .B2(n943), .C1(n49), .C2(n944), .A(n945), .ZN(
        n938) );
  AOI22_X1 U544 ( .A1(\REGISTERS[7][26] ), .A2(n52), .B1(\REGISTERS[6][26] ), 
        .B2(n53), .ZN(n945) );
  OAI221_X1 U545 ( .B1(n54), .B2(n946), .C1(n56), .C2(n947), .A(n948), .ZN(
        n937) );
  AOI22_X1 U546 ( .A1(\REGISTERS[11][26] ), .A2(n59), .B1(\REGISTERS[10][26] ), 
        .B2(n60), .ZN(n948) );
  OAI221_X1 U547 ( .B1(n61), .B2(n949), .C1(n63), .C2(n950), .A(n951), .ZN(
        n936) );
  AOI22_X1 U548 ( .A1(\REGISTERS[15][26] ), .A2(n66), .B1(\REGISTERS[14][26] ), 
        .B2(n67), .ZN(n951) );
  NAND2_X1 U549 ( .A1(n952), .A2(n953), .ZN(N4348) );
  NOR4_X1 U550 ( .A1(n954), .A2(n955), .A3(n956), .A4(n957), .ZN(n953) );
  OAI221_X1 U551 ( .B1(n8), .B2(n958), .C1(n10), .C2(n959), .A(n960), .ZN(n957) );
  AOI22_X1 U552 ( .A1(\REGISTERS[19][27] ), .A2(n13), .B1(\REGISTERS[18][27] ), 
        .B2(n14), .ZN(n960) );
  OAI221_X1 U553 ( .B1(n15), .B2(n961), .C1(n17), .C2(n962), .A(n963), .ZN(
        n956) );
  AOI22_X1 U554 ( .A1(\REGISTERS[23][27] ), .A2(n20), .B1(\REGISTERS[22][27] ), 
        .B2(n21), .ZN(n963) );
  OAI221_X1 U555 ( .B1(n22), .B2(n964), .C1(n24), .C2(n965), .A(n966), .ZN(
        n955) );
  AOI22_X1 U556 ( .A1(\REGISTERS[27][27] ), .A2(n27), .B1(\REGISTERS[26][27] ), 
        .B2(n28), .ZN(n966) );
  OAI221_X1 U557 ( .B1(n29), .B2(n967), .C1(n31), .C2(n968), .A(n969), .ZN(
        n954) );
  AOI22_X1 U558 ( .A1(\REGISTERS[29][27] ), .A2(n34), .B1(\REGISTERS[28][27] ), 
        .B2(n35), .ZN(n969) );
  NOR4_X1 U559 ( .A1(n970), .A2(n971), .A3(n972), .A4(n973), .ZN(n952) );
  AOI22_X1 U561 ( .A1(\REGISTERS[3][27] ), .A2(n45), .B1(\REGISTERS[2][27] ), 
        .B2(n46), .ZN(n976) );
  OAI221_X1 U562 ( .B1(n47), .B2(n977), .C1(n49), .C2(n978), .A(n979), .ZN(
        n972) );
  AOI22_X1 U563 ( .A1(\REGISTERS[7][27] ), .A2(n52), .B1(\REGISTERS[6][27] ), 
        .B2(n53), .ZN(n979) );
  OAI221_X1 U564 ( .B1(n54), .B2(n980), .C1(n56), .C2(n981), .A(n982), .ZN(
        n971) );
  AOI22_X1 U565 ( .A1(\REGISTERS[11][27] ), .A2(n59), .B1(\REGISTERS[10][27] ), 
        .B2(n60), .ZN(n982) );
  OAI221_X1 U566 ( .B1(n61), .B2(n983), .C1(n63), .C2(n984), .A(n985), .ZN(
        n970) );
  AOI22_X1 U567 ( .A1(\REGISTERS[15][27] ), .A2(n66), .B1(\REGISTERS[14][27] ), 
        .B2(n67), .ZN(n985) );
  NAND2_X1 U568 ( .A1(n986), .A2(n987), .ZN(N4347) );
  NOR4_X1 U569 ( .A1(n988), .A2(n989), .A3(n990), .A4(n991), .ZN(n987) );
  OAI221_X1 U570 ( .B1(n8), .B2(n992), .C1(n10), .C2(n993), .A(n994), .ZN(n991) );
  AOI22_X1 U571 ( .A1(\REGISTERS[19][28] ), .A2(n13), .B1(\REGISTERS[18][28] ), 
        .B2(n14), .ZN(n994) );
  OAI221_X1 U572 ( .B1(n15), .B2(n995), .C1(n17), .C2(n996), .A(n997), .ZN(
        n990) );
  AOI22_X1 U573 ( .A1(\REGISTERS[23][28] ), .A2(n20), .B1(\REGISTERS[22][28] ), 
        .B2(n21), .ZN(n997) );
  OAI221_X1 U574 ( .B1(n22), .B2(n998), .C1(n24), .C2(n999), .A(n1000), .ZN(
        n989) );
  AOI22_X1 U575 ( .A1(\REGISTERS[27][28] ), .A2(n27), .B1(\REGISTERS[26][28] ), 
        .B2(n28), .ZN(n1000) );
  OAI221_X1 U576 ( .B1(n29), .B2(n1001), .C1(n31), .C2(n1002), .A(n1003), .ZN(
        n988) );
  AOI22_X1 U577 ( .A1(\REGISTERS[29][28] ), .A2(n34), .B1(\REGISTERS[28][28] ), 
        .B2(n35), .ZN(n1003) );
  NOR4_X1 U578 ( .A1(n1004), .A2(n1005), .A3(n1006), .A4(n1007), .ZN(n986) );
  AOI22_X1 U580 ( .A1(\REGISTERS[3][28] ), .A2(n45), .B1(\REGISTERS[2][28] ), 
        .B2(n46), .ZN(n1010) );
  OAI221_X1 U581 ( .B1(n47), .B2(n1011), .C1(n49), .C2(n1012), .A(n1013), .ZN(
        n1006) );
  AOI22_X1 U582 ( .A1(\REGISTERS[7][28] ), .A2(n52), .B1(\REGISTERS[6][28] ), 
        .B2(n53), .ZN(n1013) );
  OAI221_X1 U583 ( .B1(n54), .B2(n1014), .C1(n56), .C2(n1015), .A(n1016), .ZN(
        n1005) );
  AOI22_X1 U584 ( .A1(\REGISTERS[11][28] ), .A2(n59), .B1(\REGISTERS[10][28] ), 
        .B2(n60), .ZN(n1016) );
  OAI221_X1 U585 ( .B1(n61), .B2(n1017), .C1(n63), .C2(n1018), .A(n1019), .ZN(
        n1004) );
  AOI22_X1 U586 ( .A1(\REGISTERS[15][28] ), .A2(n66), .B1(\REGISTERS[14][28] ), 
        .B2(n67), .ZN(n1019) );
  NAND2_X1 U587 ( .A1(n1020), .A2(n1021), .ZN(N4346) );
  NOR4_X1 U588 ( .A1(n1022), .A2(n1023), .A3(n1024), .A4(n1025), .ZN(n1021) );
  OAI221_X1 U589 ( .B1(n8), .B2(n1026), .C1(n10), .C2(n1027), .A(n1028), .ZN(
        n1025) );
  AOI22_X1 U590 ( .A1(\REGISTERS[19][29] ), .A2(n13), .B1(\REGISTERS[18][29] ), 
        .B2(n14), .ZN(n1028) );
  OAI221_X1 U591 ( .B1(n15), .B2(n1029), .C1(n17), .C2(n1030), .A(n1031), .ZN(
        n1024) );
  AOI22_X1 U592 ( .A1(\REGISTERS[23][29] ), .A2(n20), .B1(\REGISTERS[22][29] ), 
        .B2(n21), .ZN(n1031) );
  OAI221_X1 U593 ( .B1(n22), .B2(n1032), .C1(n24), .C2(n1033), .A(n1034), .ZN(
        n1023) );
  AOI22_X1 U594 ( .A1(\REGISTERS[27][29] ), .A2(n27), .B1(\REGISTERS[26][29] ), 
        .B2(n28), .ZN(n1034) );
  OAI221_X1 U595 ( .B1(n29), .B2(n1035), .C1(n31), .C2(n1036), .A(n1037), .ZN(
        n1022) );
  AOI22_X1 U596 ( .A1(\REGISTERS[29][29] ), .A2(n34), .B1(\REGISTERS[28][29] ), 
        .B2(n35), .ZN(n1037) );
  NOR4_X1 U597 ( .A1(n1038), .A2(n1039), .A3(n1040), .A4(n1041), .ZN(n1020) );
  AOI22_X1 U599 ( .A1(\REGISTERS[3][29] ), .A2(n45), .B1(\REGISTERS[2][29] ), 
        .B2(n46), .ZN(n1044) );
  OAI221_X1 U600 ( .B1(n47), .B2(n1045), .C1(n49), .C2(n1046), .A(n1047), .ZN(
        n1040) );
  AOI22_X1 U601 ( .A1(\REGISTERS[7][29] ), .A2(n52), .B1(\REGISTERS[6][29] ), 
        .B2(n53), .ZN(n1047) );
  OAI221_X1 U602 ( .B1(n54), .B2(n1048), .C1(n56), .C2(n1049), .A(n1050), .ZN(
        n1039) );
  AOI22_X1 U603 ( .A1(\REGISTERS[11][29] ), .A2(n59), .B1(\REGISTERS[10][29] ), 
        .B2(n60), .ZN(n1050) );
  OAI221_X1 U604 ( .B1(n61), .B2(n1051), .C1(n63), .C2(n1052), .A(n1053), .ZN(
        n1038) );
  AOI22_X1 U605 ( .A1(\REGISTERS[15][29] ), .A2(n66), .B1(\REGISTERS[14][29] ), 
        .B2(n67), .ZN(n1053) );
  NAND2_X1 U606 ( .A1(n1054), .A2(n1055), .ZN(N4345) );
  NOR4_X1 U607 ( .A1(n1056), .A2(n1057), .A3(n1058), .A4(n1059), .ZN(n1055) );
  OAI221_X1 U608 ( .B1(n8), .B2(n1060), .C1(n10), .C2(n1061), .A(n1062), .ZN(
        n1059) );
  AOI22_X1 U609 ( .A1(\REGISTERS[19][30] ), .A2(n13), .B1(\REGISTERS[18][30] ), 
        .B2(n14), .ZN(n1062) );
  OAI221_X1 U610 ( .B1(n15), .B2(n1063), .C1(n17), .C2(n1064), .A(n1065), .ZN(
        n1058) );
  AOI22_X1 U611 ( .A1(\REGISTERS[23][30] ), .A2(n20), .B1(\REGISTERS[22][30] ), 
        .B2(n21), .ZN(n1065) );
  OAI221_X1 U612 ( .B1(n22), .B2(n1066), .C1(n24), .C2(n1067), .A(n1068), .ZN(
        n1057) );
  AOI22_X1 U613 ( .A1(\REGISTERS[27][30] ), .A2(n27), .B1(\REGISTERS[26][30] ), 
        .B2(n28), .ZN(n1068) );
  OAI221_X1 U614 ( .B1(n29), .B2(n1069), .C1(n31), .C2(n1070), .A(n1071), .ZN(
        n1056) );
  AOI22_X1 U615 ( .A1(\REGISTERS[29][30] ), .A2(n34), .B1(\REGISTERS[28][30] ), 
        .B2(n35), .ZN(n1071) );
  NOR4_X1 U616 ( .A1(n1072), .A2(n1073), .A3(n1074), .A4(n1075), .ZN(n1054) );
  AOI22_X1 U618 ( .A1(\REGISTERS[3][30] ), .A2(n45), .B1(\REGISTERS[2][30] ), 
        .B2(n46), .ZN(n1078) );
  OAI221_X1 U619 ( .B1(n47), .B2(n1079), .C1(n49), .C2(n1080), .A(n1081), .ZN(
        n1074) );
  AOI22_X1 U620 ( .A1(\REGISTERS[7][30] ), .A2(n52), .B1(\REGISTERS[6][30] ), 
        .B2(n53), .ZN(n1081) );
  OAI221_X1 U621 ( .B1(n54), .B2(n1082), .C1(n56), .C2(n1083), .A(n1084), .ZN(
        n1073) );
  AOI22_X1 U622 ( .A1(\REGISTERS[11][30] ), .A2(n59), .B1(\REGISTERS[10][30] ), 
        .B2(n60), .ZN(n1084) );
  OAI221_X1 U623 ( .B1(n61), .B2(n1085), .C1(n63), .C2(n1086), .A(n1087), .ZN(
        n1072) );
  AOI22_X1 U624 ( .A1(\REGISTERS[15][30] ), .A2(n66), .B1(\REGISTERS[14][30] ), 
        .B2(n67), .ZN(n1087) );
  NAND2_X1 U625 ( .A1(n1088), .A2(n1089), .ZN(N4344) );
  NOR4_X1 U626 ( .A1(n1090), .A2(n1091), .A3(n1092), .A4(n1093), .ZN(n1089) );
  OAI221_X1 U627 ( .B1(n8), .B2(n1094), .C1(n10), .C2(n1095), .A(n1096), .ZN(
        n1093) );
  AOI22_X1 U628 ( .A1(\REGISTERS[19][31] ), .A2(n13), .B1(\REGISTERS[18][31] ), 
        .B2(n14), .ZN(n1096) );
  OAI221_X1 U633 ( .B1(n15), .B2(n1101), .C1(n17), .C2(n1102), .A(n1103), .ZN(
        n1092) );
  AOI22_X1 U634 ( .A1(\REGISTERS[23][31] ), .A2(n20), .B1(\REGISTERS[22][31] ), 
        .B2(n21), .ZN(n1103) );
  AND2_X1 U638 ( .A1(n1106), .A2(n1107), .ZN(n1097) );
  AND2_X1 U640 ( .A1(n1106), .A2(ADD_RD2[0]), .ZN(n1099) );
  AND2_X1 U641 ( .A1(ADD_RD2[4]), .A2(n1108), .ZN(n1106) );
  OAI221_X1 U642 ( .B1(n22), .B2(n1109), .C1(n24), .C2(n1110), .A(n1111), .ZN(
        n1091) );
  AOI22_X1 U643 ( .A1(\REGISTERS[27][31] ), .A2(n27), .B1(\REGISTERS[26][31] ), 
        .B2(n28), .ZN(n1111) );
  OAI221_X1 U648 ( .B1(n29), .B2(n1114), .C1(n31), .C2(n1115), .A(n1116), .ZN(
        n1090) );
  AOI22_X1 U649 ( .A1(\REGISTERS[29][31] ), .A2(n34), .B1(\REGISTERS[28][31] ), 
        .B2(n35), .ZN(n1116) );
  AND2_X1 U653 ( .A1(n1117), .A2(n1107), .ZN(n1112) );
  AND2_X1 U655 ( .A1(ADD_RD2[0]), .A2(n1117), .ZN(n1113) );
  AND2_X1 U656 ( .A1(ADD_RD2[4]), .A2(ADD_RD2[3]), .ZN(n1117) );
  NOR4_X1 U657 ( .A1(n1118), .A2(n1119), .A3(n1120), .A4(n1121), .ZN(n1088) );
  AOI22_X1 U659 ( .A1(\REGISTERS[3][31] ), .A2(n45), .B1(\REGISTERS[2][31] ), 
        .B2(n46), .ZN(n1124) );
  OAI221_X1 U664 ( .B1(n47), .B2(n1127), .C1(n49), .C2(n1128), .A(n1129), .ZN(
        n1120) );
  AOI22_X1 U665 ( .A1(\REGISTERS[7][31] ), .A2(n52), .B1(\REGISTERS[6][31] ), 
        .B2(n53), .ZN(n1129) );
  AND2_X1 U669 ( .A1(n1130), .A2(n1107), .ZN(n1125) );
  AND2_X1 U671 ( .A1(n1130), .A2(ADD_RD2[0]), .ZN(n1126) );
  NOR2_X1 U672 ( .A1(ADD_RD2[3]), .A2(ADD_RD2[4]), .ZN(n1130) );
  OAI221_X1 U673 ( .B1(n54), .B2(n1131), .C1(n56), .C2(n1132), .A(n1133), .ZN(
        n1119) );
  AOI22_X1 U674 ( .A1(\REGISTERS[11][31] ), .A2(n59), .B1(\REGISTERS[10][31] ), 
        .B2(n60), .ZN(n1133) );
  NOR2_X1 U677 ( .A1(n1136), .A2(ADD_RD2[2]), .ZN(n1098) );
  NOR2_X1 U680 ( .A1(ADD_RD2[1]), .A2(ADD_RD2[2]), .ZN(n1100) );
  OAI221_X1 U681 ( .B1(n61), .B2(n1137), .C1(n63), .C2(n1138), .A(n1139), .ZN(
        n1118) );
  AOI22_X1 U682 ( .A1(\REGISTERS[15][31] ), .A2(n66), .B1(\REGISTERS[14][31] ), 
        .B2(n67), .ZN(n1139) );
  NOR2_X1 U685 ( .A1(n1140), .A2(n1136), .ZN(n1104) );
  INV_X1 U686 ( .A(ADD_RD2[1]), .ZN(n1136) );
  AND2_X1 U688 ( .A1(n1141), .A2(n1107), .ZN(n1134) );
  INV_X1 U689 ( .A(ADD_RD2[0]), .ZN(n1107) );
  INV_X1 U692 ( .A(ADD_RD2[2]), .ZN(n1140) );
  AND2_X1 U693 ( .A1(n1141), .A2(ADD_RD2[0]), .ZN(n1135) );
  NOR2_X1 U694 ( .A1(n1108), .A2(ADD_RD2[4]), .ZN(n1141) );
  INV_X1 U695 ( .A(ADD_RD2[3]), .ZN(n1108) );
  AND2_X1 U696 ( .A1(RD1), .A2(ENABLE), .ZN(N4278) );
  NAND2_X1 U697 ( .A1(n1142), .A2(n1143), .ZN(N4246) );
  NOR4_X1 U698 ( .A1(n1144), .A2(n1145), .A3(n1146), .A4(n1147), .ZN(n1143) );
  OAI221_X1 U699 ( .B1(n9), .B2(n1148), .C1(n11), .C2(n1149), .A(n1150), .ZN(
        n1147) );
  AOI22_X1 U700 ( .A1(n1151), .A2(\REGISTERS[19][0] ), .B1(n1152), .B2(
        \REGISTERS[18][0] ), .ZN(n1150) );
  INV_X1 U701 ( .A(\REGISTERS[16][0] ), .ZN(n11) );
  INV_X1 U702 ( .A(\REGISTERS[17][0] ), .ZN(n9) );
  OAI221_X1 U703 ( .B1(n16), .B2(n1153), .C1(n18), .C2(n1154), .A(n1155), .ZN(
        n1146) );
  AOI22_X1 U704 ( .A1(n1156), .A2(\REGISTERS[23][0] ), .B1(n1157), .B2(
        \REGISTERS[22][0] ), .ZN(n1155) );
  INV_X1 U705 ( .A(\REGISTERS[20][0] ), .ZN(n18) );
  INV_X1 U706 ( .A(\REGISTERS[21][0] ), .ZN(n16) );
  OAI221_X1 U707 ( .B1(n23), .B2(n1158), .C1(n25), .C2(n1159), .A(n1160), .ZN(
        n1145) );
  AOI22_X1 U708 ( .A1(n1161), .A2(\REGISTERS[27][0] ), .B1(n1162), .B2(
        \REGISTERS[26][0] ), .ZN(n1160) );
  INV_X1 U709 ( .A(\REGISTERS[24][0] ), .ZN(n25) );
  INV_X1 U710 ( .A(\REGISTERS[25][0] ), .ZN(n23) );
  OAI221_X1 U711 ( .B1(n30), .B2(n1163), .C1(n32), .C2(n1164), .A(n1165), .ZN(
        n1144) );
  AOI22_X1 U712 ( .A1(n1166), .A2(\REGISTERS[29][0] ), .B1(n1167), .B2(
        \REGISTERS[28][0] ), .ZN(n1165) );
  INV_X1 U713 ( .A(\REGISTERS[30][0] ), .ZN(n32) );
  INV_X1 U714 ( .A(\REGISTERS[31][0] ), .ZN(n30) );
  NOR4_X1 U715 ( .A1(n1168), .A2(n1169), .A3(n1170), .A4(n1171), .ZN(n1142) );
  AOI22_X1 U717 ( .A1(n1175), .A2(\REGISTERS[3][0] ), .B1(n1176), .B2(
        \REGISTERS[2][0] ), .ZN(n1174) );
  INV_X1 U718 ( .A(\REGISTERS[1][0] ), .ZN(n41) );
  OAI221_X1 U719 ( .B1(n48), .B2(n1177), .C1(n50), .C2(n1178), .A(n1179), .ZN(
        n1170) );
  AOI22_X1 U720 ( .A1(n1180), .A2(\REGISTERS[7][0] ), .B1(n1181), .B2(
        \REGISTERS[6][0] ), .ZN(n1179) );
  INV_X1 U721 ( .A(\REGISTERS[4][0] ), .ZN(n50) );
  INV_X1 U722 ( .A(\REGISTERS[5][0] ), .ZN(n48) );
  OAI221_X1 U723 ( .B1(n55), .B2(n1182), .C1(n57), .C2(n1183), .A(n1184), .ZN(
        n1169) );
  AOI22_X1 U724 ( .A1(n1185), .A2(\REGISTERS[11][0] ), .B1(n1186), .B2(
        \REGISTERS[10][0] ), .ZN(n1184) );
  INV_X1 U725 ( .A(\REGISTERS[8][0] ), .ZN(n57) );
  INV_X1 U726 ( .A(\REGISTERS[9][0] ), .ZN(n55) );
  OAI221_X1 U727 ( .B1(n62), .B2(n1187), .C1(n64), .C2(n1188), .A(n1189), .ZN(
        n1168) );
  AOI22_X1 U728 ( .A1(n1190), .A2(\REGISTERS[15][0] ), .B1(n1191), .B2(
        \REGISTERS[14][0] ), .ZN(n1189) );
  INV_X1 U729 ( .A(\REGISTERS[12][0] ), .ZN(n64) );
  INV_X1 U730 ( .A(\REGISTERS[13][0] ), .ZN(n62) );
  NAND2_X1 U731 ( .A1(n1192), .A2(n1193), .ZN(N4245) );
  NOR4_X1 U732 ( .A1(n1194), .A2(n1195), .A3(n1196), .A4(n1197), .ZN(n1193) );
  OAI221_X1 U733 ( .B1(n74), .B2(n1148), .C1(n75), .C2(n1149), .A(n1198), .ZN(
        n1197) );
  AOI22_X1 U734 ( .A1(n1151), .A2(\REGISTERS[19][1] ), .B1(n1152), .B2(
        \REGISTERS[18][1] ), .ZN(n1198) );
  INV_X1 U735 ( .A(\REGISTERS[16][1] ), .ZN(n75) );
  INV_X1 U736 ( .A(\REGISTERS[17][1] ), .ZN(n74) );
  OAI221_X1 U737 ( .B1(n77), .B2(n1153), .C1(n78), .C2(n1154), .A(n1199), .ZN(
        n1196) );
  AOI22_X1 U738 ( .A1(n1156), .A2(\REGISTERS[23][1] ), .B1(n1157), .B2(
        \REGISTERS[22][1] ), .ZN(n1199) );
  INV_X1 U739 ( .A(\REGISTERS[20][1] ), .ZN(n78) );
  INV_X1 U740 ( .A(\REGISTERS[21][1] ), .ZN(n77) );
  OAI221_X1 U741 ( .B1(n80), .B2(n1158), .C1(n81), .C2(n1159), .A(n1200), .ZN(
        n1195) );
  AOI22_X1 U742 ( .A1(n1161), .A2(\REGISTERS[27][1] ), .B1(n1162), .B2(
        \REGISTERS[26][1] ), .ZN(n1200) );
  INV_X1 U743 ( .A(\REGISTERS[24][1] ), .ZN(n81) );
  INV_X1 U744 ( .A(\REGISTERS[25][1] ), .ZN(n80) );
  OAI221_X1 U745 ( .B1(n83), .B2(n1163), .C1(n84), .C2(n1164), .A(n1201), .ZN(
        n1194) );
  AOI22_X1 U746 ( .A1(n1166), .A2(\REGISTERS[29][1] ), .B1(n1167), .B2(
        \REGISTERS[28][1] ), .ZN(n1201) );
  INV_X1 U747 ( .A(\REGISTERS[30][1] ), .ZN(n84) );
  INV_X1 U748 ( .A(\REGISTERS[31][1] ), .ZN(n83) );
  NOR4_X1 U749 ( .A1(n1202), .A2(n1203), .A3(n1204), .A4(n1205), .ZN(n1192) );
  AOI22_X1 U751 ( .A1(n1175), .A2(\REGISTERS[3][1] ), .B1(n1176), .B2(
        \REGISTERS[2][1] ), .ZN(n1206) );
  INV_X1 U752 ( .A(\REGISTERS[1][1] ), .ZN(n90) );
  OAI221_X1 U753 ( .B1(n93), .B2(n1177), .C1(n94), .C2(n1178), .A(n1207), .ZN(
        n1204) );
  AOI22_X1 U754 ( .A1(n1180), .A2(\REGISTERS[7][1] ), .B1(n1181), .B2(
        \REGISTERS[6][1] ), .ZN(n1207) );
  INV_X1 U755 ( .A(\REGISTERS[4][1] ), .ZN(n94) );
  INV_X1 U756 ( .A(\REGISTERS[5][1] ), .ZN(n93) );
  OAI221_X1 U757 ( .B1(n96), .B2(n1182), .C1(n97), .C2(n1183), .A(n1208), .ZN(
        n1203) );
  AOI22_X1 U758 ( .A1(n1185), .A2(\REGISTERS[11][1] ), .B1(n1186), .B2(
        \REGISTERS[10][1] ), .ZN(n1208) );
  INV_X1 U759 ( .A(\REGISTERS[8][1] ), .ZN(n97) );
  INV_X1 U760 ( .A(\REGISTERS[9][1] ), .ZN(n96) );
  OAI221_X1 U761 ( .B1(n99), .B2(n1187), .C1(n100), .C2(n1188), .A(n1209), 
        .ZN(n1202) );
  AOI22_X1 U762 ( .A1(n1190), .A2(\REGISTERS[15][1] ), .B1(n1191), .B2(
        \REGISTERS[14][1] ), .ZN(n1209) );
  INV_X1 U763 ( .A(\REGISTERS[12][1] ), .ZN(n100) );
  INV_X1 U764 ( .A(\REGISTERS[13][1] ), .ZN(n99) );
  NAND2_X1 U765 ( .A1(n1210), .A2(n1211), .ZN(N4244) );
  NOR4_X1 U766 ( .A1(n1212), .A2(n1213), .A3(n1214), .A4(n1215), .ZN(n1211) );
  OAI221_X1 U767 ( .B1(n108), .B2(n1148), .C1(n109), .C2(n1149), .A(n1216), 
        .ZN(n1215) );
  AOI22_X1 U768 ( .A1(n1151), .A2(\REGISTERS[19][2] ), .B1(n1152), .B2(
        \REGISTERS[18][2] ), .ZN(n1216) );
  INV_X1 U769 ( .A(\REGISTERS[16][2] ), .ZN(n109) );
  INV_X1 U770 ( .A(\REGISTERS[17][2] ), .ZN(n108) );
  OAI221_X1 U771 ( .B1(n111), .B2(n1153), .C1(n112), .C2(n1154), .A(n1217), 
        .ZN(n1214) );
  AOI22_X1 U772 ( .A1(n1156), .A2(\REGISTERS[23][2] ), .B1(n1157), .B2(
        \REGISTERS[22][2] ), .ZN(n1217) );
  INV_X1 U773 ( .A(\REGISTERS[20][2] ), .ZN(n112) );
  INV_X1 U774 ( .A(\REGISTERS[21][2] ), .ZN(n111) );
  OAI221_X1 U775 ( .B1(n114), .B2(n1158), .C1(n115), .C2(n1159), .A(n1218), 
        .ZN(n1213) );
  AOI22_X1 U776 ( .A1(n1161), .A2(\REGISTERS[27][2] ), .B1(n1162), .B2(
        \REGISTERS[26][2] ), .ZN(n1218) );
  INV_X1 U777 ( .A(\REGISTERS[24][2] ), .ZN(n115) );
  INV_X1 U778 ( .A(\REGISTERS[25][2] ), .ZN(n114) );
  OAI221_X1 U779 ( .B1(n117), .B2(n1163), .C1(n118), .C2(n1164), .A(n1219), 
        .ZN(n1212) );
  AOI22_X1 U780 ( .A1(n1166), .A2(\REGISTERS[29][2] ), .B1(n1167), .B2(
        \REGISTERS[28][2] ), .ZN(n1219) );
  INV_X1 U781 ( .A(\REGISTERS[30][2] ), .ZN(n118) );
  INV_X1 U782 ( .A(\REGISTERS[31][2] ), .ZN(n117) );
  NOR4_X1 U783 ( .A1(n1220), .A2(n1221), .A3(n1222), .A4(n1223), .ZN(n1210) );
  AOI22_X1 U785 ( .A1(n1175), .A2(\REGISTERS[3][2] ), .B1(n1176), .B2(
        \REGISTERS[2][2] ), .ZN(n1224) );
  INV_X1 U786 ( .A(\REGISTERS[1][2] ), .ZN(n124) );
  OAI221_X1 U787 ( .B1(n127), .B2(n1177), .C1(n128), .C2(n1178), .A(n1225), 
        .ZN(n1222) );
  AOI22_X1 U788 ( .A1(n1180), .A2(\REGISTERS[7][2] ), .B1(n1181), .B2(
        \REGISTERS[6][2] ), .ZN(n1225) );
  INV_X1 U789 ( .A(\REGISTERS[4][2] ), .ZN(n128) );
  INV_X1 U790 ( .A(\REGISTERS[5][2] ), .ZN(n127) );
  OAI221_X1 U791 ( .B1(n130), .B2(n1182), .C1(n131), .C2(n1183), .A(n1226), 
        .ZN(n1221) );
  AOI22_X1 U792 ( .A1(n1185), .A2(\REGISTERS[11][2] ), .B1(n1186), .B2(
        \REGISTERS[10][2] ), .ZN(n1226) );
  INV_X1 U793 ( .A(\REGISTERS[8][2] ), .ZN(n131) );
  INV_X1 U794 ( .A(\REGISTERS[9][2] ), .ZN(n130) );
  OAI221_X1 U795 ( .B1(n133), .B2(n1187), .C1(n134), .C2(n1188), .A(n1227), 
        .ZN(n1220) );
  AOI22_X1 U796 ( .A1(n1190), .A2(\REGISTERS[15][2] ), .B1(n1191), .B2(
        \REGISTERS[14][2] ), .ZN(n1227) );
  INV_X1 U797 ( .A(\REGISTERS[12][2] ), .ZN(n134) );
  INV_X1 U798 ( .A(\REGISTERS[13][2] ), .ZN(n133) );
  NAND2_X1 U799 ( .A1(n1228), .A2(n1229), .ZN(N4243) );
  NOR4_X1 U800 ( .A1(n1230), .A2(n1231), .A3(n1232), .A4(n1233), .ZN(n1229) );
  OAI221_X1 U801 ( .B1(n142), .B2(n1148), .C1(n143), .C2(n1149), .A(n1234), 
        .ZN(n1233) );
  AOI22_X1 U802 ( .A1(n1151), .A2(\REGISTERS[19][3] ), .B1(n1152), .B2(
        \REGISTERS[18][3] ), .ZN(n1234) );
  INV_X1 U803 ( .A(\REGISTERS[16][3] ), .ZN(n143) );
  INV_X1 U804 ( .A(\REGISTERS[17][3] ), .ZN(n142) );
  OAI221_X1 U805 ( .B1(n145), .B2(n1153), .C1(n146), .C2(n1154), .A(n1235), 
        .ZN(n1232) );
  AOI22_X1 U806 ( .A1(n1156), .A2(\REGISTERS[23][3] ), .B1(n1157), .B2(
        \REGISTERS[22][3] ), .ZN(n1235) );
  INV_X1 U807 ( .A(\REGISTERS[20][3] ), .ZN(n146) );
  INV_X1 U808 ( .A(\REGISTERS[21][3] ), .ZN(n145) );
  OAI221_X1 U809 ( .B1(n148), .B2(n1158), .C1(n149), .C2(n1159), .A(n1236), 
        .ZN(n1231) );
  AOI22_X1 U810 ( .A1(n1161), .A2(\REGISTERS[27][3] ), .B1(n1162), .B2(
        \REGISTERS[26][3] ), .ZN(n1236) );
  INV_X1 U811 ( .A(\REGISTERS[24][3] ), .ZN(n149) );
  INV_X1 U812 ( .A(\REGISTERS[25][3] ), .ZN(n148) );
  OAI221_X1 U813 ( .B1(n151), .B2(n1163), .C1(n152), .C2(n1164), .A(n1237), 
        .ZN(n1230) );
  AOI22_X1 U814 ( .A1(n1166), .A2(\REGISTERS[29][3] ), .B1(n1167), .B2(
        \REGISTERS[28][3] ), .ZN(n1237) );
  INV_X1 U815 ( .A(\REGISTERS[30][3] ), .ZN(n152) );
  INV_X1 U816 ( .A(\REGISTERS[31][3] ), .ZN(n151) );
  NOR4_X1 U817 ( .A1(n1238), .A2(n1239), .A3(n1240), .A4(n1241), .ZN(n1228) );
  AOI22_X1 U819 ( .A1(n1175), .A2(\REGISTERS[3][3] ), .B1(n1176), .B2(
        \REGISTERS[2][3] ), .ZN(n1242) );
  INV_X1 U820 ( .A(\REGISTERS[1][3] ), .ZN(n158) );
  OAI221_X1 U821 ( .B1(n161), .B2(n1177), .C1(n162), .C2(n1178), .A(n1243), 
        .ZN(n1240) );
  AOI22_X1 U822 ( .A1(n1180), .A2(\REGISTERS[7][3] ), .B1(n1181), .B2(
        \REGISTERS[6][3] ), .ZN(n1243) );
  INV_X1 U823 ( .A(\REGISTERS[4][3] ), .ZN(n162) );
  INV_X1 U824 ( .A(\REGISTERS[5][3] ), .ZN(n161) );
  OAI221_X1 U825 ( .B1(n164), .B2(n1182), .C1(n165), .C2(n1183), .A(n1244), 
        .ZN(n1239) );
  AOI22_X1 U826 ( .A1(n1185), .A2(\REGISTERS[11][3] ), .B1(n1186), .B2(
        \REGISTERS[10][3] ), .ZN(n1244) );
  INV_X1 U827 ( .A(\REGISTERS[8][3] ), .ZN(n165) );
  INV_X1 U828 ( .A(\REGISTERS[9][3] ), .ZN(n164) );
  OAI221_X1 U829 ( .B1(n167), .B2(n1187), .C1(n168), .C2(n1188), .A(n1245), 
        .ZN(n1238) );
  AOI22_X1 U830 ( .A1(n1190), .A2(\REGISTERS[15][3] ), .B1(n1191), .B2(
        \REGISTERS[14][3] ), .ZN(n1245) );
  INV_X1 U831 ( .A(\REGISTERS[12][3] ), .ZN(n168) );
  INV_X1 U832 ( .A(\REGISTERS[13][3] ), .ZN(n167) );
  NAND2_X1 U833 ( .A1(n1246), .A2(n1247), .ZN(N4242) );
  NOR4_X1 U834 ( .A1(n1248), .A2(n1249), .A3(n1250), .A4(n1251), .ZN(n1247) );
  OAI221_X1 U835 ( .B1(n176), .B2(n1148), .C1(n177), .C2(n1149), .A(n1252), 
        .ZN(n1251) );
  AOI22_X1 U836 ( .A1(n1151), .A2(\REGISTERS[19][4] ), .B1(n1152), .B2(
        \REGISTERS[18][4] ), .ZN(n1252) );
  INV_X1 U837 ( .A(\REGISTERS[16][4] ), .ZN(n177) );
  INV_X1 U838 ( .A(\REGISTERS[17][4] ), .ZN(n176) );
  OAI221_X1 U839 ( .B1(n179), .B2(n1153), .C1(n180), .C2(n1154), .A(n1253), 
        .ZN(n1250) );
  AOI22_X1 U840 ( .A1(n1156), .A2(\REGISTERS[23][4] ), .B1(n1157), .B2(
        \REGISTERS[22][4] ), .ZN(n1253) );
  INV_X1 U841 ( .A(\REGISTERS[20][4] ), .ZN(n180) );
  INV_X1 U842 ( .A(\REGISTERS[21][4] ), .ZN(n179) );
  OAI221_X1 U843 ( .B1(n182), .B2(n1158), .C1(n183), .C2(n1159), .A(n1254), 
        .ZN(n1249) );
  AOI22_X1 U844 ( .A1(n1161), .A2(\REGISTERS[27][4] ), .B1(n1162), .B2(
        \REGISTERS[26][4] ), .ZN(n1254) );
  INV_X1 U845 ( .A(\REGISTERS[24][4] ), .ZN(n183) );
  INV_X1 U846 ( .A(\REGISTERS[25][4] ), .ZN(n182) );
  OAI221_X1 U847 ( .B1(n185), .B2(n1163), .C1(n186), .C2(n1164), .A(n1255), 
        .ZN(n1248) );
  AOI22_X1 U848 ( .A1(n1166), .A2(\REGISTERS[29][4] ), .B1(n1167), .B2(
        \REGISTERS[28][4] ), .ZN(n1255) );
  INV_X1 U849 ( .A(\REGISTERS[30][4] ), .ZN(n186) );
  INV_X1 U850 ( .A(\REGISTERS[31][4] ), .ZN(n185) );
  NOR4_X1 U851 ( .A1(n1256), .A2(n1257), .A3(n1258), .A4(n1259), .ZN(n1246) );
  AOI22_X1 U853 ( .A1(n1175), .A2(\REGISTERS[3][4] ), .B1(n1176), .B2(
        \REGISTERS[2][4] ), .ZN(n1260) );
  INV_X1 U854 ( .A(\REGISTERS[1][4] ), .ZN(n192) );
  OAI221_X1 U855 ( .B1(n195), .B2(n1177), .C1(n196), .C2(n1178), .A(n1261), 
        .ZN(n1258) );
  AOI22_X1 U856 ( .A1(n1180), .A2(\REGISTERS[7][4] ), .B1(n1181), .B2(
        \REGISTERS[6][4] ), .ZN(n1261) );
  INV_X1 U857 ( .A(\REGISTERS[4][4] ), .ZN(n196) );
  INV_X1 U858 ( .A(\REGISTERS[5][4] ), .ZN(n195) );
  OAI221_X1 U859 ( .B1(n198), .B2(n1182), .C1(n199), .C2(n1183), .A(n1262), 
        .ZN(n1257) );
  AOI22_X1 U860 ( .A1(n1185), .A2(\REGISTERS[11][4] ), .B1(n1186), .B2(
        \REGISTERS[10][4] ), .ZN(n1262) );
  INV_X1 U861 ( .A(\REGISTERS[8][4] ), .ZN(n199) );
  INV_X1 U862 ( .A(\REGISTERS[9][4] ), .ZN(n198) );
  OAI221_X1 U863 ( .B1(n201), .B2(n1187), .C1(n202), .C2(n1188), .A(n1263), 
        .ZN(n1256) );
  AOI22_X1 U864 ( .A1(n1190), .A2(\REGISTERS[15][4] ), .B1(n1191), .B2(
        \REGISTERS[14][4] ), .ZN(n1263) );
  INV_X1 U865 ( .A(\REGISTERS[12][4] ), .ZN(n202) );
  INV_X1 U866 ( .A(\REGISTERS[13][4] ), .ZN(n201) );
  NAND2_X1 U867 ( .A1(n1264), .A2(n1265), .ZN(N4241) );
  NOR4_X1 U868 ( .A1(n1266), .A2(n1267), .A3(n1268), .A4(n1269), .ZN(n1265) );
  OAI221_X1 U869 ( .B1(n210), .B2(n1148), .C1(n211), .C2(n1149), .A(n1270), 
        .ZN(n1269) );
  AOI22_X1 U870 ( .A1(n1151), .A2(\REGISTERS[19][5] ), .B1(n1152), .B2(
        \REGISTERS[18][5] ), .ZN(n1270) );
  INV_X1 U871 ( .A(\REGISTERS[16][5] ), .ZN(n211) );
  INV_X1 U872 ( .A(\REGISTERS[17][5] ), .ZN(n210) );
  OAI221_X1 U873 ( .B1(n213), .B2(n1153), .C1(n214), .C2(n1154), .A(n1271), 
        .ZN(n1268) );
  AOI22_X1 U874 ( .A1(n1156), .A2(\REGISTERS[23][5] ), .B1(n1157), .B2(
        \REGISTERS[22][5] ), .ZN(n1271) );
  INV_X1 U875 ( .A(\REGISTERS[20][5] ), .ZN(n214) );
  INV_X1 U876 ( .A(\REGISTERS[21][5] ), .ZN(n213) );
  OAI221_X1 U877 ( .B1(n216), .B2(n1158), .C1(n217), .C2(n1159), .A(n1272), 
        .ZN(n1267) );
  AOI22_X1 U878 ( .A1(n1161), .A2(\REGISTERS[27][5] ), .B1(n1162), .B2(
        \REGISTERS[26][5] ), .ZN(n1272) );
  INV_X1 U879 ( .A(\REGISTERS[24][5] ), .ZN(n217) );
  INV_X1 U880 ( .A(\REGISTERS[25][5] ), .ZN(n216) );
  OAI221_X1 U881 ( .B1(n219), .B2(n1163), .C1(n220), .C2(n1164), .A(n1273), 
        .ZN(n1266) );
  AOI22_X1 U882 ( .A1(n1166), .A2(\REGISTERS[29][5] ), .B1(n1167), .B2(
        \REGISTERS[28][5] ), .ZN(n1273) );
  INV_X1 U883 ( .A(\REGISTERS[30][5] ), .ZN(n220) );
  INV_X1 U884 ( .A(\REGISTERS[31][5] ), .ZN(n219) );
  NOR4_X1 U885 ( .A1(n1274), .A2(n1275), .A3(n1276), .A4(n1277), .ZN(n1264) );
  AOI22_X1 U887 ( .A1(n1175), .A2(\REGISTERS[3][5] ), .B1(n1176), .B2(
        \REGISTERS[2][5] ), .ZN(n1278) );
  INV_X1 U888 ( .A(\REGISTERS[1][5] ), .ZN(n226) );
  OAI221_X1 U889 ( .B1(n229), .B2(n1177), .C1(n230), .C2(n1178), .A(n1279), 
        .ZN(n1276) );
  AOI22_X1 U890 ( .A1(n1180), .A2(\REGISTERS[7][5] ), .B1(n1181), .B2(
        \REGISTERS[6][5] ), .ZN(n1279) );
  INV_X1 U891 ( .A(\REGISTERS[4][5] ), .ZN(n230) );
  INV_X1 U892 ( .A(\REGISTERS[5][5] ), .ZN(n229) );
  OAI221_X1 U893 ( .B1(n232), .B2(n1182), .C1(n233), .C2(n1183), .A(n1280), 
        .ZN(n1275) );
  AOI22_X1 U894 ( .A1(n1185), .A2(\REGISTERS[11][5] ), .B1(n1186), .B2(
        \REGISTERS[10][5] ), .ZN(n1280) );
  INV_X1 U895 ( .A(\REGISTERS[8][5] ), .ZN(n233) );
  INV_X1 U896 ( .A(\REGISTERS[9][5] ), .ZN(n232) );
  OAI221_X1 U897 ( .B1(n235), .B2(n1187), .C1(n236), .C2(n1188), .A(n1281), 
        .ZN(n1274) );
  AOI22_X1 U898 ( .A1(n1190), .A2(\REGISTERS[15][5] ), .B1(n1191), .B2(
        \REGISTERS[14][5] ), .ZN(n1281) );
  INV_X1 U899 ( .A(\REGISTERS[12][5] ), .ZN(n236) );
  INV_X1 U900 ( .A(\REGISTERS[13][5] ), .ZN(n235) );
  NAND2_X1 U901 ( .A1(n1282), .A2(n1283), .ZN(N4240) );
  NOR4_X1 U902 ( .A1(n1284), .A2(n1285), .A3(n1286), .A4(n1287), .ZN(n1283) );
  OAI221_X1 U903 ( .B1(n244), .B2(n1148), .C1(n245), .C2(n1149), .A(n1288), 
        .ZN(n1287) );
  AOI22_X1 U904 ( .A1(n1151), .A2(\REGISTERS[19][6] ), .B1(n1152), .B2(
        \REGISTERS[18][6] ), .ZN(n1288) );
  INV_X1 U905 ( .A(\REGISTERS[16][6] ), .ZN(n245) );
  INV_X1 U906 ( .A(\REGISTERS[17][6] ), .ZN(n244) );
  OAI221_X1 U907 ( .B1(n247), .B2(n1153), .C1(n248), .C2(n1154), .A(n1289), 
        .ZN(n1286) );
  AOI22_X1 U908 ( .A1(n1156), .A2(\REGISTERS[23][6] ), .B1(n1157), .B2(
        \REGISTERS[22][6] ), .ZN(n1289) );
  INV_X1 U909 ( .A(\REGISTERS[20][6] ), .ZN(n248) );
  INV_X1 U910 ( .A(\REGISTERS[21][6] ), .ZN(n247) );
  OAI221_X1 U911 ( .B1(n250), .B2(n1158), .C1(n251), .C2(n1159), .A(n1290), 
        .ZN(n1285) );
  AOI22_X1 U912 ( .A1(n1161), .A2(\REGISTERS[27][6] ), .B1(n1162), .B2(
        \REGISTERS[26][6] ), .ZN(n1290) );
  INV_X1 U913 ( .A(\REGISTERS[24][6] ), .ZN(n251) );
  INV_X1 U914 ( .A(\REGISTERS[25][6] ), .ZN(n250) );
  OAI221_X1 U915 ( .B1(n253), .B2(n1163), .C1(n254), .C2(n1164), .A(n1291), 
        .ZN(n1284) );
  AOI22_X1 U916 ( .A1(n1166), .A2(\REGISTERS[29][6] ), .B1(n1167), .B2(
        \REGISTERS[28][6] ), .ZN(n1291) );
  INV_X1 U917 ( .A(\REGISTERS[30][6] ), .ZN(n254) );
  INV_X1 U918 ( .A(\REGISTERS[31][6] ), .ZN(n253) );
  NOR4_X1 U919 ( .A1(n1292), .A2(n1293), .A3(n1294), .A4(n1295), .ZN(n1282) );
  AOI22_X1 U921 ( .A1(n1175), .A2(\REGISTERS[3][6] ), .B1(n1176), .B2(
        \REGISTERS[2][6] ), .ZN(n1296) );
  INV_X1 U922 ( .A(\REGISTERS[1][6] ), .ZN(n260) );
  OAI221_X1 U923 ( .B1(n263), .B2(n1177), .C1(n264), .C2(n1178), .A(n1297), 
        .ZN(n1294) );
  AOI22_X1 U924 ( .A1(n1180), .A2(\REGISTERS[7][6] ), .B1(n1181), .B2(
        \REGISTERS[6][6] ), .ZN(n1297) );
  INV_X1 U925 ( .A(\REGISTERS[4][6] ), .ZN(n264) );
  INV_X1 U926 ( .A(\REGISTERS[5][6] ), .ZN(n263) );
  OAI221_X1 U927 ( .B1(n266), .B2(n1182), .C1(n267), .C2(n1183), .A(n1298), 
        .ZN(n1293) );
  AOI22_X1 U928 ( .A1(n1185), .A2(\REGISTERS[11][6] ), .B1(n1186), .B2(
        \REGISTERS[10][6] ), .ZN(n1298) );
  INV_X1 U929 ( .A(\REGISTERS[8][6] ), .ZN(n267) );
  INV_X1 U930 ( .A(\REGISTERS[9][6] ), .ZN(n266) );
  OAI221_X1 U931 ( .B1(n269), .B2(n1187), .C1(n270), .C2(n1188), .A(n1299), 
        .ZN(n1292) );
  AOI22_X1 U932 ( .A1(n1190), .A2(\REGISTERS[15][6] ), .B1(n1191), .B2(
        \REGISTERS[14][6] ), .ZN(n1299) );
  INV_X1 U933 ( .A(\REGISTERS[12][6] ), .ZN(n270) );
  INV_X1 U934 ( .A(\REGISTERS[13][6] ), .ZN(n269) );
  NAND2_X1 U935 ( .A1(n1300), .A2(n1301), .ZN(N4239) );
  NOR4_X1 U936 ( .A1(n1302), .A2(n1303), .A3(n1304), .A4(n1305), .ZN(n1301) );
  OAI221_X1 U937 ( .B1(n278), .B2(n1148), .C1(n279), .C2(n1149), .A(n1306), 
        .ZN(n1305) );
  AOI22_X1 U938 ( .A1(n1151), .A2(\REGISTERS[19][7] ), .B1(n1152), .B2(
        \REGISTERS[18][7] ), .ZN(n1306) );
  INV_X1 U939 ( .A(\REGISTERS[16][7] ), .ZN(n279) );
  INV_X1 U940 ( .A(\REGISTERS[17][7] ), .ZN(n278) );
  OAI221_X1 U941 ( .B1(n281), .B2(n1153), .C1(n282), .C2(n1154), .A(n1307), 
        .ZN(n1304) );
  AOI22_X1 U942 ( .A1(n1156), .A2(\REGISTERS[23][7] ), .B1(n1157), .B2(
        \REGISTERS[22][7] ), .ZN(n1307) );
  INV_X1 U943 ( .A(\REGISTERS[20][7] ), .ZN(n282) );
  INV_X1 U944 ( .A(\REGISTERS[21][7] ), .ZN(n281) );
  OAI221_X1 U945 ( .B1(n284), .B2(n1158), .C1(n285), .C2(n1159), .A(n1308), 
        .ZN(n1303) );
  AOI22_X1 U946 ( .A1(n1161), .A2(\REGISTERS[27][7] ), .B1(n1162), .B2(
        \REGISTERS[26][7] ), .ZN(n1308) );
  INV_X1 U947 ( .A(\REGISTERS[24][7] ), .ZN(n285) );
  INV_X1 U948 ( .A(\REGISTERS[25][7] ), .ZN(n284) );
  OAI221_X1 U949 ( .B1(n287), .B2(n1163), .C1(n288), .C2(n1164), .A(n1309), 
        .ZN(n1302) );
  AOI22_X1 U950 ( .A1(n1166), .A2(\REGISTERS[29][7] ), .B1(n1167), .B2(
        \REGISTERS[28][7] ), .ZN(n1309) );
  INV_X1 U951 ( .A(\REGISTERS[30][7] ), .ZN(n288) );
  INV_X1 U952 ( .A(\REGISTERS[31][7] ), .ZN(n287) );
  NOR4_X1 U953 ( .A1(n1310), .A2(n1311), .A3(n1312), .A4(n1313), .ZN(n1300) );
  AOI22_X1 U955 ( .A1(n1175), .A2(\REGISTERS[3][7] ), .B1(n1176), .B2(
        \REGISTERS[2][7] ), .ZN(n1314) );
  INV_X1 U956 ( .A(\REGISTERS[1][7] ), .ZN(n294) );
  OAI221_X1 U957 ( .B1(n297), .B2(n1177), .C1(n298), .C2(n1178), .A(n1315), 
        .ZN(n1312) );
  AOI22_X1 U958 ( .A1(n1180), .A2(\REGISTERS[7][7] ), .B1(n1181), .B2(
        \REGISTERS[6][7] ), .ZN(n1315) );
  INV_X1 U959 ( .A(\REGISTERS[4][7] ), .ZN(n298) );
  INV_X1 U960 ( .A(\REGISTERS[5][7] ), .ZN(n297) );
  OAI221_X1 U961 ( .B1(n300), .B2(n1182), .C1(n301), .C2(n1183), .A(n1316), 
        .ZN(n1311) );
  AOI22_X1 U962 ( .A1(n1185), .A2(\REGISTERS[11][7] ), .B1(n1186), .B2(
        \REGISTERS[10][7] ), .ZN(n1316) );
  INV_X1 U963 ( .A(\REGISTERS[8][7] ), .ZN(n301) );
  INV_X1 U964 ( .A(\REGISTERS[9][7] ), .ZN(n300) );
  OAI221_X1 U965 ( .B1(n303), .B2(n1187), .C1(n304), .C2(n1188), .A(n1317), 
        .ZN(n1310) );
  AOI22_X1 U966 ( .A1(n1190), .A2(\REGISTERS[15][7] ), .B1(n1191), .B2(
        \REGISTERS[14][7] ), .ZN(n1317) );
  INV_X1 U967 ( .A(\REGISTERS[12][7] ), .ZN(n304) );
  INV_X1 U968 ( .A(\REGISTERS[13][7] ), .ZN(n303) );
  NAND2_X1 U969 ( .A1(n1318), .A2(n1319), .ZN(N4238) );
  NOR4_X1 U970 ( .A1(n1320), .A2(n1321), .A3(n1322), .A4(n1323), .ZN(n1319) );
  OAI221_X1 U971 ( .B1(n312), .B2(n1148), .C1(n313), .C2(n1149), .A(n1324), 
        .ZN(n1323) );
  AOI22_X1 U972 ( .A1(n1151), .A2(\REGISTERS[19][8] ), .B1(n1152), .B2(
        \REGISTERS[18][8] ), .ZN(n1324) );
  INV_X1 U973 ( .A(\REGISTERS[16][8] ), .ZN(n313) );
  INV_X1 U974 ( .A(\REGISTERS[17][8] ), .ZN(n312) );
  OAI221_X1 U975 ( .B1(n315), .B2(n1153), .C1(n316), .C2(n1154), .A(n1325), 
        .ZN(n1322) );
  AOI22_X1 U976 ( .A1(n1156), .A2(\REGISTERS[23][8] ), .B1(n1157), .B2(
        \REGISTERS[22][8] ), .ZN(n1325) );
  INV_X1 U977 ( .A(\REGISTERS[20][8] ), .ZN(n316) );
  INV_X1 U978 ( .A(\REGISTERS[21][8] ), .ZN(n315) );
  OAI221_X1 U979 ( .B1(n318), .B2(n1158), .C1(n319), .C2(n1159), .A(n1326), 
        .ZN(n1321) );
  AOI22_X1 U980 ( .A1(n1161), .A2(\REGISTERS[27][8] ), .B1(n1162), .B2(
        \REGISTERS[26][8] ), .ZN(n1326) );
  INV_X1 U981 ( .A(\REGISTERS[24][8] ), .ZN(n319) );
  INV_X1 U982 ( .A(\REGISTERS[25][8] ), .ZN(n318) );
  OAI221_X1 U983 ( .B1(n321), .B2(n1163), .C1(n322), .C2(n1164), .A(n1327), 
        .ZN(n1320) );
  AOI22_X1 U984 ( .A1(n1166), .A2(\REGISTERS[29][8] ), .B1(n1167), .B2(
        \REGISTERS[28][8] ), .ZN(n1327) );
  INV_X1 U985 ( .A(\REGISTERS[30][8] ), .ZN(n322) );
  INV_X1 U986 ( .A(\REGISTERS[31][8] ), .ZN(n321) );
  NOR4_X1 U987 ( .A1(n1328), .A2(n1329), .A3(n1330), .A4(n1331), .ZN(n1318) );
  AOI22_X1 U989 ( .A1(n1175), .A2(\REGISTERS[3][8] ), .B1(n1176), .B2(
        \REGISTERS[2][8] ), .ZN(n1332) );
  INV_X1 U990 ( .A(\REGISTERS[1][8] ), .ZN(n328) );
  OAI221_X1 U991 ( .B1(n331), .B2(n1177), .C1(n332), .C2(n1178), .A(n1333), 
        .ZN(n1330) );
  AOI22_X1 U992 ( .A1(n1180), .A2(\REGISTERS[7][8] ), .B1(n1181), .B2(
        \REGISTERS[6][8] ), .ZN(n1333) );
  INV_X1 U993 ( .A(\REGISTERS[4][8] ), .ZN(n332) );
  INV_X1 U994 ( .A(\REGISTERS[5][8] ), .ZN(n331) );
  OAI221_X1 U995 ( .B1(n334), .B2(n1182), .C1(n335), .C2(n1183), .A(n1334), 
        .ZN(n1329) );
  AOI22_X1 U996 ( .A1(n1185), .A2(\REGISTERS[11][8] ), .B1(n1186), .B2(
        \REGISTERS[10][8] ), .ZN(n1334) );
  INV_X1 U997 ( .A(\REGISTERS[8][8] ), .ZN(n335) );
  INV_X1 U998 ( .A(\REGISTERS[9][8] ), .ZN(n334) );
  OAI221_X1 U999 ( .B1(n337), .B2(n1187), .C1(n338), .C2(n1188), .A(n1335), 
        .ZN(n1328) );
  AOI22_X1 U1000 ( .A1(n1190), .A2(\REGISTERS[15][8] ), .B1(n1191), .B2(
        \REGISTERS[14][8] ), .ZN(n1335) );
  INV_X1 U1001 ( .A(\REGISTERS[12][8] ), .ZN(n338) );
  INV_X1 U1002 ( .A(\REGISTERS[13][8] ), .ZN(n337) );
  NAND2_X1 U1003 ( .A1(n1336), .A2(n1337), .ZN(N4237) );
  NOR4_X1 U1004 ( .A1(n1338), .A2(n1339), .A3(n1340), .A4(n1341), .ZN(n1337)
         );
  OAI221_X1 U1005 ( .B1(n346), .B2(n1148), .C1(n347), .C2(n1149), .A(n1342), 
        .ZN(n1341) );
  AOI22_X1 U1006 ( .A1(n1151), .A2(\REGISTERS[19][9] ), .B1(n1152), .B2(
        \REGISTERS[18][9] ), .ZN(n1342) );
  INV_X1 U1007 ( .A(\REGISTERS[16][9] ), .ZN(n347) );
  INV_X1 U1008 ( .A(\REGISTERS[17][9] ), .ZN(n346) );
  OAI221_X1 U1009 ( .B1(n349), .B2(n1153), .C1(n350), .C2(n1154), .A(n1343), 
        .ZN(n1340) );
  AOI22_X1 U1010 ( .A1(n1156), .A2(\REGISTERS[23][9] ), .B1(n1157), .B2(
        \REGISTERS[22][9] ), .ZN(n1343) );
  INV_X1 U1011 ( .A(\REGISTERS[20][9] ), .ZN(n350) );
  INV_X1 U1012 ( .A(\REGISTERS[21][9] ), .ZN(n349) );
  OAI221_X1 U1013 ( .B1(n352), .B2(n1158), .C1(n353), .C2(n1159), .A(n1344), 
        .ZN(n1339) );
  AOI22_X1 U1014 ( .A1(n1161), .A2(\REGISTERS[27][9] ), .B1(n1162), .B2(
        \REGISTERS[26][9] ), .ZN(n1344) );
  INV_X1 U1015 ( .A(\REGISTERS[24][9] ), .ZN(n353) );
  INV_X1 U1016 ( .A(\REGISTERS[25][9] ), .ZN(n352) );
  OAI221_X1 U1017 ( .B1(n355), .B2(n1163), .C1(n356), .C2(n1164), .A(n1345), 
        .ZN(n1338) );
  AOI22_X1 U1018 ( .A1(n1166), .A2(\REGISTERS[29][9] ), .B1(n1167), .B2(
        \REGISTERS[28][9] ), .ZN(n1345) );
  INV_X1 U1019 ( .A(\REGISTERS[30][9] ), .ZN(n356) );
  INV_X1 U1020 ( .A(\REGISTERS[31][9] ), .ZN(n355) );
  NOR4_X1 U1021 ( .A1(n1346), .A2(n1347), .A3(n1348), .A4(n1349), .ZN(n1336)
         );
  AOI22_X1 U1023 ( .A1(n1175), .A2(\REGISTERS[3][9] ), .B1(n1176), .B2(
        \REGISTERS[2][9] ), .ZN(n1350) );
  INV_X1 U1024 ( .A(\REGISTERS[1][9] ), .ZN(n362) );
  OAI221_X1 U1025 ( .B1(n365), .B2(n1177), .C1(n366), .C2(n1178), .A(n1351), 
        .ZN(n1348) );
  AOI22_X1 U1026 ( .A1(n1180), .A2(\REGISTERS[7][9] ), .B1(n1181), .B2(
        \REGISTERS[6][9] ), .ZN(n1351) );
  INV_X1 U1027 ( .A(\REGISTERS[4][9] ), .ZN(n366) );
  INV_X1 U1028 ( .A(\REGISTERS[5][9] ), .ZN(n365) );
  OAI221_X1 U1029 ( .B1(n368), .B2(n1182), .C1(n369), .C2(n1183), .A(n1352), 
        .ZN(n1347) );
  AOI22_X1 U1030 ( .A1(n1185), .A2(\REGISTERS[11][9] ), .B1(n1186), .B2(
        \REGISTERS[10][9] ), .ZN(n1352) );
  INV_X1 U1031 ( .A(\REGISTERS[8][9] ), .ZN(n369) );
  INV_X1 U1032 ( .A(\REGISTERS[9][9] ), .ZN(n368) );
  OAI221_X1 U1033 ( .B1(n371), .B2(n1187), .C1(n372), .C2(n1188), .A(n1353), 
        .ZN(n1346) );
  AOI22_X1 U1034 ( .A1(n1190), .A2(\REGISTERS[15][9] ), .B1(n1191), .B2(
        \REGISTERS[14][9] ), .ZN(n1353) );
  INV_X1 U1035 ( .A(\REGISTERS[12][9] ), .ZN(n372) );
  INV_X1 U1036 ( .A(\REGISTERS[13][9] ), .ZN(n371) );
  NAND2_X1 U1037 ( .A1(n1354), .A2(n1355), .ZN(N4236) );
  NOR4_X1 U1038 ( .A1(n1356), .A2(n1357), .A3(n1358), .A4(n1359), .ZN(n1355)
         );
  OAI221_X1 U1039 ( .B1(n380), .B2(n1148), .C1(n381), .C2(n1149), .A(n1360), 
        .ZN(n1359) );
  AOI22_X1 U1040 ( .A1(n1151), .A2(\REGISTERS[19][10] ), .B1(n1152), .B2(
        \REGISTERS[18][10] ), .ZN(n1360) );
  INV_X1 U1041 ( .A(\REGISTERS[16][10] ), .ZN(n381) );
  INV_X1 U1042 ( .A(\REGISTERS[17][10] ), .ZN(n380) );
  OAI221_X1 U1043 ( .B1(n383), .B2(n1153), .C1(n384), .C2(n1154), .A(n1361), 
        .ZN(n1358) );
  AOI22_X1 U1044 ( .A1(n1156), .A2(\REGISTERS[23][10] ), .B1(n1157), .B2(
        \REGISTERS[22][10] ), .ZN(n1361) );
  INV_X1 U1045 ( .A(\REGISTERS[20][10] ), .ZN(n384) );
  INV_X1 U1046 ( .A(\REGISTERS[21][10] ), .ZN(n383) );
  OAI221_X1 U1047 ( .B1(n386), .B2(n1158), .C1(n387), .C2(n1159), .A(n1362), 
        .ZN(n1357) );
  AOI22_X1 U1048 ( .A1(n1161), .A2(\REGISTERS[27][10] ), .B1(n1162), .B2(
        \REGISTERS[26][10] ), .ZN(n1362) );
  INV_X1 U1049 ( .A(\REGISTERS[24][10] ), .ZN(n387) );
  INV_X1 U1050 ( .A(\REGISTERS[25][10] ), .ZN(n386) );
  OAI221_X1 U1051 ( .B1(n389), .B2(n1163), .C1(n390), .C2(n1164), .A(n1363), 
        .ZN(n1356) );
  AOI22_X1 U1052 ( .A1(n1166), .A2(\REGISTERS[29][10] ), .B1(n1167), .B2(
        \REGISTERS[28][10] ), .ZN(n1363) );
  INV_X1 U1053 ( .A(\REGISTERS[30][10] ), .ZN(n390) );
  INV_X1 U1054 ( .A(\REGISTERS[31][10] ), .ZN(n389) );
  NOR4_X1 U1055 ( .A1(n1364), .A2(n1365), .A3(n1366), .A4(n1367), .ZN(n1354)
         );
  AOI22_X1 U1057 ( .A1(n1175), .A2(\REGISTERS[3][10] ), .B1(n1176), .B2(
        \REGISTERS[2][10] ), .ZN(n1368) );
  INV_X1 U1058 ( .A(\REGISTERS[1][10] ), .ZN(n396) );
  OAI221_X1 U1059 ( .B1(n399), .B2(n1177), .C1(n400), .C2(n1178), .A(n1369), 
        .ZN(n1366) );
  AOI22_X1 U1060 ( .A1(n1180), .A2(\REGISTERS[7][10] ), .B1(n1181), .B2(
        \REGISTERS[6][10] ), .ZN(n1369) );
  INV_X1 U1061 ( .A(\REGISTERS[4][10] ), .ZN(n400) );
  INV_X1 U1062 ( .A(\REGISTERS[5][10] ), .ZN(n399) );
  OAI221_X1 U1063 ( .B1(n402), .B2(n1182), .C1(n403), .C2(n1183), .A(n1370), 
        .ZN(n1365) );
  AOI22_X1 U1064 ( .A1(n1185), .A2(\REGISTERS[11][10] ), .B1(n1186), .B2(
        \REGISTERS[10][10] ), .ZN(n1370) );
  INV_X1 U1065 ( .A(\REGISTERS[8][10] ), .ZN(n403) );
  INV_X1 U1066 ( .A(\REGISTERS[9][10] ), .ZN(n402) );
  OAI221_X1 U1067 ( .B1(n405), .B2(n1187), .C1(n406), .C2(n1188), .A(n1371), 
        .ZN(n1364) );
  AOI22_X1 U1068 ( .A1(n1190), .A2(\REGISTERS[15][10] ), .B1(n1191), .B2(
        \REGISTERS[14][10] ), .ZN(n1371) );
  INV_X1 U1069 ( .A(\REGISTERS[12][10] ), .ZN(n406) );
  INV_X1 U1070 ( .A(\REGISTERS[13][10] ), .ZN(n405) );
  NAND2_X1 U1071 ( .A1(n1372), .A2(n1373), .ZN(N4235) );
  NOR4_X1 U1072 ( .A1(n1374), .A2(n1375), .A3(n1376), .A4(n1377), .ZN(n1373)
         );
  OAI221_X1 U1073 ( .B1(n414), .B2(n1148), .C1(n415), .C2(n1149), .A(n1378), 
        .ZN(n1377) );
  AOI22_X1 U1074 ( .A1(n1151), .A2(\REGISTERS[19][11] ), .B1(n1152), .B2(
        \REGISTERS[18][11] ), .ZN(n1378) );
  INV_X1 U1075 ( .A(\REGISTERS[16][11] ), .ZN(n415) );
  INV_X1 U1076 ( .A(\REGISTERS[17][11] ), .ZN(n414) );
  OAI221_X1 U1077 ( .B1(n417), .B2(n1153), .C1(n418), .C2(n1154), .A(n1379), 
        .ZN(n1376) );
  AOI22_X1 U1078 ( .A1(n1156), .A2(\REGISTERS[23][11] ), .B1(n1157), .B2(
        \REGISTERS[22][11] ), .ZN(n1379) );
  INV_X1 U1079 ( .A(\REGISTERS[20][11] ), .ZN(n418) );
  INV_X1 U1080 ( .A(\REGISTERS[21][11] ), .ZN(n417) );
  OAI221_X1 U1081 ( .B1(n420), .B2(n1158), .C1(n421), .C2(n1159), .A(n1380), 
        .ZN(n1375) );
  AOI22_X1 U1082 ( .A1(n1161), .A2(\REGISTERS[27][11] ), .B1(n1162), .B2(
        \REGISTERS[26][11] ), .ZN(n1380) );
  INV_X1 U1083 ( .A(\REGISTERS[24][11] ), .ZN(n421) );
  INV_X1 U1084 ( .A(\REGISTERS[25][11] ), .ZN(n420) );
  OAI221_X1 U1085 ( .B1(n423), .B2(n1163), .C1(n424), .C2(n1164), .A(n1381), 
        .ZN(n1374) );
  AOI22_X1 U1086 ( .A1(n1166), .A2(\REGISTERS[29][11] ), .B1(n1167), .B2(
        \REGISTERS[28][11] ), .ZN(n1381) );
  INV_X1 U1087 ( .A(\REGISTERS[30][11] ), .ZN(n424) );
  INV_X1 U1088 ( .A(\REGISTERS[31][11] ), .ZN(n423) );
  NOR4_X1 U1089 ( .A1(n1382), .A2(n1383), .A3(n1384), .A4(n1385), .ZN(n1372)
         );
  AOI22_X1 U1091 ( .A1(n1175), .A2(\REGISTERS[3][11] ), .B1(n1176), .B2(
        \REGISTERS[2][11] ), .ZN(n1386) );
  INV_X1 U1092 ( .A(\REGISTERS[1][11] ), .ZN(n430) );
  OAI221_X1 U1093 ( .B1(n433), .B2(n1177), .C1(n434), .C2(n1178), .A(n1387), 
        .ZN(n1384) );
  AOI22_X1 U1094 ( .A1(n1180), .A2(\REGISTERS[7][11] ), .B1(n1181), .B2(
        \REGISTERS[6][11] ), .ZN(n1387) );
  INV_X1 U1095 ( .A(\REGISTERS[4][11] ), .ZN(n434) );
  INV_X1 U1096 ( .A(\REGISTERS[5][11] ), .ZN(n433) );
  OAI221_X1 U1097 ( .B1(n436), .B2(n1182), .C1(n437), .C2(n1183), .A(n1388), 
        .ZN(n1383) );
  AOI22_X1 U1098 ( .A1(n1185), .A2(\REGISTERS[11][11] ), .B1(n1186), .B2(
        \REGISTERS[10][11] ), .ZN(n1388) );
  INV_X1 U1099 ( .A(\REGISTERS[8][11] ), .ZN(n437) );
  INV_X1 U1100 ( .A(\REGISTERS[9][11] ), .ZN(n436) );
  OAI221_X1 U1101 ( .B1(n439), .B2(n1187), .C1(n440), .C2(n1188), .A(n1389), 
        .ZN(n1382) );
  AOI22_X1 U1102 ( .A1(n1190), .A2(\REGISTERS[15][11] ), .B1(n1191), .B2(
        \REGISTERS[14][11] ), .ZN(n1389) );
  INV_X1 U1103 ( .A(\REGISTERS[12][11] ), .ZN(n440) );
  INV_X1 U1104 ( .A(\REGISTERS[13][11] ), .ZN(n439) );
  NAND2_X1 U1105 ( .A1(n1390), .A2(n1391), .ZN(N4234) );
  NOR4_X1 U1106 ( .A1(n1392), .A2(n1393), .A3(n1394), .A4(n1395), .ZN(n1391)
         );
  OAI221_X1 U1107 ( .B1(n448), .B2(n1148), .C1(n449), .C2(n1149), .A(n1396), 
        .ZN(n1395) );
  AOI22_X1 U1108 ( .A1(n1151), .A2(\REGISTERS[19][12] ), .B1(n1152), .B2(
        \REGISTERS[18][12] ), .ZN(n1396) );
  INV_X1 U1109 ( .A(\REGISTERS[16][12] ), .ZN(n449) );
  INV_X1 U1110 ( .A(\REGISTERS[17][12] ), .ZN(n448) );
  OAI221_X1 U1111 ( .B1(n451), .B2(n1153), .C1(n452), .C2(n1154), .A(n1397), 
        .ZN(n1394) );
  AOI22_X1 U1112 ( .A1(n1156), .A2(\REGISTERS[23][12] ), .B1(n1157), .B2(
        \REGISTERS[22][12] ), .ZN(n1397) );
  INV_X1 U1113 ( .A(\REGISTERS[20][12] ), .ZN(n452) );
  INV_X1 U1114 ( .A(\REGISTERS[21][12] ), .ZN(n451) );
  OAI221_X1 U1115 ( .B1(n454), .B2(n1158), .C1(n455), .C2(n1159), .A(n1398), 
        .ZN(n1393) );
  AOI22_X1 U1116 ( .A1(n1161), .A2(\REGISTERS[27][12] ), .B1(n1162), .B2(
        \REGISTERS[26][12] ), .ZN(n1398) );
  INV_X1 U1117 ( .A(\REGISTERS[24][12] ), .ZN(n455) );
  INV_X1 U1118 ( .A(\REGISTERS[25][12] ), .ZN(n454) );
  OAI221_X1 U1119 ( .B1(n457), .B2(n1163), .C1(n458), .C2(n1164), .A(n1399), 
        .ZN(n1392) );
  AOI22_X1 U1120 ( .A1(n1166), .A2(\REGISTERS[29][12] ), .B1(n1167), .B2(
        \REGISTERS[28][12] ), .ZN(n1399) );
  INV_X1 U1121 ( .A(\REGISTERS[30][12] ), .ZN(n458) );
  INV_X1 U1122 ( .A(\REGISTERS[31][12] ), .ZN(n457) );
  NOR4_X1 U1123 ( .A1(n1400), .A2(n1401), .A3(n1402), .A4(n1403), .ZN(n1390)
         );
  AOI22_X1 U1125 ( .A1(n1175), .A2(\REGISTERS[3][12] ), .B1(n1176), .B2(
        \REGISTERS[2][12] ), .ZN(n1404) );
  INV_X1 U1126 ( .A(\REGISTERS[1][12] ), .ZN(n464) );
  OAI221_X1 U1127 ( .B1(n467), .B2(n1177), .C1(n468), .C2(n1178), .A(n1405), 
        .ZN(n1402) );
  AOI22_X1 U1128 ( .A1(n1180), .A2(\REGISTERS[7][12] ), .B1(n1181), .B2(
        \REGISTERS[6][12] ), .ZN(n1405) );
  INV_X1 U1129 ( .A(\REGISTERS[4][12] ), .ZN(n468) );
  INV_X1 U1130 ( .A(\REGISTERS[5][12] ), .ZN(n467) );
  OAI221_X1 U1131 ( .B1(n470), .B2(n1182), .C1(n471), .C2(n1183), .A(n1406), 
        .ZN(n1401) );
  AOI22_X1 U1132 ( .A1(n1185), .A2(\REGISTERS[11][12] ), .B1(n1186), .B2(
        \REGISTERS[10][12] ), .ZN(n1406) );
  INV_X1 U1133 ( .A(\REGISTERS[8][12] ), .ZN(n471) );
  INV_X1 U1134 ( .A(\REGISTERS[9][12] ), .ZN(n470) );
  OAI221_X1 U1135 ( .B1(n473), .B2(n1187), .C1(n474), .C2(n1188), .A(n1407), 
        .ZN(n1400) );
  AOI22_X1 U1136 ( .A1(n1190), .A2(\REGISTERS[15][12] ), .B1(n1191), .B2(
        \REGISTERS[14][12] ), .ZN(n1407) );
  INV_X1 U1137 ( .A(\REGISTERS[12][12] ), .ZN(n474) );
  INV_X1 U1138 ( .A(\REGISTERS[13][12] ), .ZN(n473) );
  NAND2_X1 U1139 ( .A1(n1408), .A2(n1409), .ZN(N4233) );
  NOR4_X1 U1140 ( .A1(n1410), .A2(n1411), .A3(n1412), .A4(n1413), .ZN(n1409)
         );
  OAI221_X1 U1141 ( .B1(n482), .B2(n1148), .C1(n483), .C2(n1149), .A(n1414), 
        .ZN(n1413) );
  AOI22_X1 U1142 ( .A1(n1151), .A2(\REGISTERS[19][13] ), .B1(n1152), .B2(
        \REGISTERS[18][13] ), .ZN(n1414) );
  INV_X1 U1143 ( .A(\REGISTERS[16][13] ), .ZN(n483) );
  INV_X1 U1144 ( .A(\REGISTERS[17][13] ), .ZN(n482) );
  OAI221_X1 U1145 ( .B1(n485), .B2(n1153), .C1(n486), .C2(n1154), .A(n1415), 
        .ZN(n1412) );
  AOI22_X1 U1146 ( .A1(n1156), .A2(\REGISTERS[23][13] ), .B1(n1157), .B2(
        \REGISTERS[22][13] ), .ZN(n1415) );
  INV_X1 U1147 ( .A(\REGISTERS[20][13] ), .ZN(n486) );
  INV_X1 U1148 ( .A(\REGISTERS[21][13] ), .ZN(n485) );
  OAI221_X1 U1149 ( .B1(n488), .B2(n1158), .C1(n489), .C2(n1159), .A(n1416), 
        .ZN(n1411) );
  AOI22_X1 U1150 ( .A1(n1161), .A2(\REGISTERS[27][13] ), .B1(n1162), .B2(
        \REGISTERS[26][13] ), .ZN(n1416) );
  INV_X1 U1151 ( .A(\REGISTERS[24][13] ), .ZN(n489) );
  INV_X1 U1152 ( .A(\REGISTERS[25][13] ), .ZN(n488) );
  OAI221_X1 U1153 ( .B1(n491), .B2(n1163), .C1(n492), .C2(n1164), .A(n1417), 
        .ZN(n1410) );
  AOI22_X1 U1154 ( .A1(n1166), .A2(\REGISTERS[29][13] ), .B1(n1167), .B2(
        \REGISTERS[28][13] ), .ZN(n1417) );
  INV_X1 U1155 ( .A(\REGISTERS[30][13] ), .ZN(n492) );
  INV_X1 U1156 ( .A(\REGISTERS[31][13] ), .ZN(n491) );
  NOR4_X1 U1157 ( .A1(n1418), .A2(n1419), .A3(n1420), .A4(n1421), .ZN(n1408)
         );
  AOI22_X1 U1159 ( .A1(n1175), .A2(\REGISTERS[3][13] ), .B1(n1176), .B2(
        \REGISTERS[2][13] ), .ZN(n1422) );
  INV_X1 U1160 ( .A(\REGISTERS[1][13] ), .ZN(n498) );
  OAI221_X1 U1161 ( .B1(n501), .B2(n1177), .C1(n502), .C2(n1178), .A(n1423), 
        .ZN(n1420) );
  AOI22_X1 U1162 ( .A1(n1180), .A2(\REGISTERS[7][13] ), .B1(n1181), .B2(
        \REGISTERS[6][13] ), .ZN(n1423) );
  INV_X1 U1163 ( .A(\REGISTERS[4][13] ), .ZN(n502) );
  INV_X1 U1164 ( .A(\REGISTERS[5][13] ), .ZN(n501) );
  OAI221_X1 U1165 ( .B1(n504), .B2(n1182), .C1(n505), .C2(n1183), .A(n1424), 
        .ZN(n1419) );
  AOI22_X1 U1166 ( .A1(n1185), .A2(\REGISTERS[11][13] ), .B1(n1186), .B2(
        \REGISTERS[10][13] ), .ZN(n1424) );
  INV_X1 U1167 ( .A(\REGISTERS[8][13] ), .ZN(n505) );
  INV_X1 U1168 ( .A(\REGISTERS[9][13] ), .ZN(n504) );
  OAI221_X1 U1169 ( .B1(n507), .B2(n1187), .C1(n508), .C2(n1188), .A(n1425), 
        .ZN(n1418) );
  AOI22_X1 U1170 ( .A1(n1190), .A2(\REGISTERS[15][13] ), .B1(n1191), .B2(
        \REGISTERS[14][13] ), .ZN(n1425) );
  INV_X1 U1171 ( .A(\REGISTERS[12][13] ), .ZN(n508) );
  INV_X1 U1172 ( .A(\REGISTERS[13][13] ), .ZN(n507) );
  NAND2_X1 U1173 ( .A1(n1426), .A2(n1427), .ZN(N4232) );
  NOR4_X1 U1174 ( .A1(n1428), .A2(n1429), .A3(n1430), .A4(n1431), .ZN(n1427)
         );
  OAI221_X1 U1175 ( .B1(n516), .B2(n1148), .C1(n517), .C2(n1149), .A(n1432), 
        .ZN(n1431) );
  AOI22_X1 U1176 ( .A1(n1151), .A2(\REGISTERS[19][14] ), .B1(n1152), .B2(
        \REGISTERS[18][14] ), .ZN(n1432) );
  INV_X1 U1177 ( .A(\REGISTERS[16][14] ), .ZN(n517) );
  INV_X1 U1178 ( .A(\REGISTERS[17][14] ), .ZN(n516) );
  OAI221_X1 U1179 ( .B1(n519), .B2(n1153), .C1(n520), .C2(n1154), .A(n1433), 
        .ZN(n1430) );
  AOI22_X1 U1180 ( .A1(n1156), .A2(\REGISTERS[23][14] ), .B1(n1157), .B2(
        \REGISTERS[22][14] ), .ZN(n1433) );
  INV_X1 U1181 ( .A(\REGISTERS[20][14] ), .ZN(n520) );
  INV_X1 U1182 ( .A(\REGISTERS[21][14] ), .ZN(n519) );
  OAI221_X1 U1183 ( .B1(n522), .B2(n1158), .C1(n523), .C2(n1159), .A(n1434), 
        .ZN(n1429) );
  AOI22_X1 U1184 ( .A1(n1161), .A2(\REGISTERS[27][14] ), .B1(n1162), .B2(
        \REGISTERS[26][14] ), .ZN(n1434) );
  INV_X1 U1185 ( .A(\REGISTERS[24][14] ), .ZN(n523) );
  INV_X1 U1186 ( .A(\REGISTERS[25][14] ), .ZN(n522) );
  OAI221_X1 U1187 ( .B1(n525), .B2(n1163), .C1(n526), .C2(n1164), .A(n1435), 
        .ZN(n1428) );
  AOI22_X1 U1188 ( .A1(n1166), .A2(\REGISTERS[29][14] ), .B1(n1167), .B2(
        \REGISTERS[28][14] ), .ZN(n1435) );
  INV_X1 U1189 ( .A(\REGISTERS[30][14] ), .ZN(n526) );
  INV_X1 U1190 ( .A(\REGISTERS[31][14] ), .ZN(n525) );
  NOR4_X1 U1191 ( .A1(n1436), .A2(n1437), .A3(n1438), .A4(n1439), .ZN(n1426)
         );
  AOI22_X1 U1193 ( .A1(n1175), .A2(\REGISTERS[3][14] ), .B1(n1176), .B2(
        \REGISTERS[2][14] ), .ZN(n1440) );
  INV_X1 U1194 ( .A(\REGISTERS[1][14] ), .ZN(n532) );
  OAI221_X1 U1195 ( .B1(n535), .B2(n1177), .C1(n536), .C2(n1178), .A(n1441), 
        .ZN(n1438) );
  AOI22_X1 U1196 ( .A1(n1180), .A2(\REGISTERS[7][14] ), .B1(n1181), .B2(
        \REGISTERS[6][14] ), .ZN(n1441) );
  INV_X1 U1197 ( .A(\REGISTERS[4][14] ), .ZN(n536) );
  INV_X1 U1198 ( .A(\REGISTERS[5][14] ), .ZN(n535) );
  OAI221_X1 U1199 ( .B1(n538), .B2(n1182), .C1(n539), .C2(n1183), .A(n1442), 
        .ZN(n1437) );
  AOI22_X1 U1200 ( .A1(n1185), .A2(\REGISTERS[11][14] ), .B1(n1186), .B2(
        \REGISTERS[10][14] ), .ZN(n1442) );
  INV_X1 U1201 ( .A(\REGISTERS[8][14] ), .ZN(n539) );
  INV_X1 U1202 ( .A(\REGISTERS[9][14] ), .ZN(n538) );
  OAI221_X1 U1203 ( .B1(n541), .B2(n1187), .C1(n542), .C2(n1188), .A(n1443), 
        .ZN(n1436) );
  AOI22_X1 U1204 ( .A1(n1190), .A2(\REGISTERS[15][14] ), .B1(n1191), .B2(
        \REGISTERS[14][14] ), .ZN(n1443) );
  INV_X1 U1205 ( .A(\REGISTERS[12][14] ), .ZN(n542) );
  INV_X1 U1206 ( .A(\REGISTERS[13][14] ), .ZN(n541) );
  NAND2_X1 U1207 ( .A1(n1444), .A2(n1445), .ZN(N4231) );
  NOR4_X1 U1208 ( .A1(n1446), .A2(n1447), .A3(n1448), .A4(n1449), .ZN(n1445)
         );
  OAI221_X1 U1209 ( .B1(n550), .B2(n1148), .C1(n551), .C2(n1149), .A(n1450), 
        .ZN(n1449) );
  AOI22_X1 U1210 ( .A1(n1151), .A2(\REGISTERS[19][15] ), .B1(n1152), .B2(
        \REGISTERS[18][15] ), .ZN(n1450) );
  INV_X1 U1211 ( .A(\REGISTERS[16][15] ), .ZN(n551) );
  INV_X1 U1212 ( .A(\REGISTERS[17][15] ), .ZN(n550) );
  OAI221_X1 U1213 ( .B1(n553), .B2(n1153), .C1(n554), .C2(n1154), .A(n1451), 
        .ZN(n1448) );
  AOI22_X1 U1214 ( .A1(n1156), .A2(\REGISTERS[23][15] ), .B1(n1157), .B2(
        \REGISTERS[22][15] ), .ZN(n1451) );
  INV_X1 U1215 ( .A(\REGISTERS[20][15] ), .ZN(n554) );
  INV_X1 U1216 ( .A(\REGISTERS[21][15] ), .ZN(n553) );
  OAI221_X1 U1217 ( .B1(n556), .B2(n1158), .C1(n557), .C2(n1159), .A(n1452), 
        .ZN(n1447) );
  AOI22_X1 U1218 ( .A1(n1161), .A2(\REGISTERS[27][15] ), .B1(n1162), .B2(
        \REGISTERS[26][15] ), .ZN(n1452) );
  INV_X1 U1219 ( .A(\REGISTERS[24][15] ), .ZN(n557) );
  INV_X1 U1220 ( .A(\REGISTERS[25][15] ), .ZN(n556) );
  OAI221_X1 U1221 ( .B1(n559), .B2(n1163), .C1(n560), .C2(n1164), .A(n1453), 
        .ZN(n1446) );
  AOI22_X1 U1222 ( .A1(n1166), .A2(\REGISTERS[29][15] ), .B1(n1167), .B2(
        \REGISTERS[28][15] ), .ZN(n1453) );
  INV_X1 U1223 ( .A(\REGISTERS[30][15] ), .ZN(n560) );
  INV_X1 U1224 ( .A(\REGISTERS[31][15] ), .ZN(n559) );
  NOR4_X1 U1225 ( .A1(n1454), .A2(n1455), .A3(n1456), .A4(n1457), .ZN(n1444)
         );
  AOI22_X1 U1227 ( .A1(n1175), .A2(\REGISTERS[3][15] ), .B1(n1176), .B2(
        \REGISTERS[2][15] ), .ZN(n1458) );
  INV_X1 U1228 ( .A(\REGISTERS[1][15] ), .ZN(n566) );
  OAI221_X1 U1229 ( .B1(n569), .B2(n1177), .C1(n570), .C2(n1178), .A(n1459), 
        .ZN(n1456) );
  AOI22_X1 U1230 ( .A1(n1180), .A2(\REGISTERS[7][15] ), .B1(n1181), .B2(
        \REGISTERS[6][15] ), .ZN(n1459) );
  INV_X1 U1231 ( .A(\REGISTERS[4][15] ), .ZN(n570) );
  INV_X1 U1232 ( .A(\REGISTERS[5][15] ), .ZN(n569) );
  OAI221_X1 U1233 ( .B1(n572), .B2(n1182), .C1(n573), .C2(n1183), .A(n1460), 
        .ZN(n1455) );
  AOI22_X1 U1234 ( .A1(n1185), .A2(\REGISTERS[11][15] ), .B1(n1186), .B2(
        \REGISTERS[10][15] ), .ZN(n1460) );
  INV_X1 U1235 ( .A(\REGISTERS[8][15] ), .ZN(n573) );
  INV_X1 U1236 ( .A(\REGISTERS[9][15] ), .ZN(n572) );
  OAI221_X1 U1237 ( .B1(n575), .B2(n1187), .C1(n576), .C2(n1188), .A(n1461), 
        .ZN(n1454) );
  AOI22_X1 U1238 ( .A1(n1190), .A2(\REGISTERS[15][15] ), .B1(n1191), .B2(
        \REGISTERS[14][15] ), .ZN(n1461) );
  INV_X1 U1239 ( .A(\REGISTERS[12][15] ), .ZN(n576) );
  INV_X1 U1240 ( .A(\REGISTERS[13][15] ), .ZN(n575) );
  NAND2_X1 U1241 ( .A1(n1462), .A2(n1463), .ZN(N4230) );
  NOR4_X1 U1242 ( .A1(n1464), .A2(n1465), .A3(n1466), .A4(n1467), .ZN(n1463)
         );
  OAI221_X1 U1243 ( .B1(n584), .B2(n1148), .C1(n585), .C2(n1149), .A(n1468), 
        .ZN(n1467) );
  AOI22_X1 U1244 ( .A1(n1151), .A2(\REGISTERS[19][16] ), .B1(n1152), .B2(
        \REGISTERS[18][16] ), .ZN(n1468) );
  INV_X1 U1245 ( .A(\REGISTERS[16][16] ), .ZN(n585) );
  INV_X1 U1246 ( .A(\REGISTERS[17][16] ), .ZN(n584) );
  OAI221_X1 U1247 ( .B1(n587), .B2(n1153), .C1(n588), .C2(n1154), .A(n1469), 
        .ZN(n1466) );
  AOI22_X1 U1248 ( .A1(n1156), .A2(\REGISTERS[23][16] ), .B1(n1157), .B2(
        \REGISTERS[22][16] ), .ZN(n1469) );
  INV_X1 U1249 ( .A(\REGISTERS[20][16] ), .ZN(n588) );
  INV_X1 U1250 ( .A(\REGISTERS[21][16] ), .ZN(n587) );
  OAI221_X1 U1251 ( .B1(n590), .B2(n1158), .C1(n591), .C2(n1159), .A(n1470), 
        .ZN(n1465) );
  AOI22_X1 U1252 ( .A1(n1161), .A2(\REGISTERS[27][16] ), .B1(n1162), .B2(
        \REGISTERS[26][16] ), .ZN(n1470) );
  INV_X1 U1253 ( .A(\REGISTERS[24][16] ), .ZN(n591) );
  INV_X1 U1254 ( .A(\REGISTERS[25][16] ), .ZN(n590) );
  OAI221_X1 U1255 ( .B1(n593), .B2(n1163), .C1(n594), .C2(n1164), .A(n1471), 
        .ZN(n1464) );
  AOI22_X1 U1256 ( .A1(n1166), .A2(\REGISTERS[29][16] ), .B1(n1167), .B2(
        \REGISTERS[28][16] ), .ZN(n1471) );
  INV_X1 U1257 ( .A(\REGISTERS[30][16] ), .ZN(n594) );
  INV_X1 U1258 ( .A(\REGISTERS[31][16] ), .ZN(n593) );
  NOR4_X1 U1259 ( .A1(n1472), .A2(n1473), .A3(n1474), .A4(n1475), .ZN(n1462)
         );
  AOI22_X1 U1261 ( .A1(n1175), .A2(\REGISTERS[3][16] ), .B1(n1176), .B2(
        \REGISTERS[2][16] ), .ZN(n1476) );
  INV_X1 U1262 ( .A(\REGISTERS[1][16] ), .ZN(n600) );
  OAI221_X1 U1263 ( .B1(n603), .B2(n1177), .C1(n604), .C2(n1178), .A(n1477), 
        .ZN(n1474) );
  AOI22_X1 U1264 ( .A1(n1180), .A2(\REGISTERS[7][16] ), .B1(n1181), .B2(
        \REGISTERS[6][16] ), .ZN(n1477) );
  INV_X1 U1265 ( .A(\REGISTERS[4][16] ), .ZN(n604) );
  INV_X1 U1266 ( .A(\REGISTERS[5][16] ), .ZN(n603) );
  OAI221_X1 U1267 ( .B1(n606), .B2(n1182), .C1(n607), .C2(n1183), .A(n1478), 
        .ZN(n1473) );
  AOI22_X1 U1268 ( .A1(n1185), .A2(\REGISTERS[11][16] ), .B1(n1186), .B2(
        \REGISTERS[10][16] ), .ZN(n1478) );
  INV_X1 U1269 ( .A(\REGISTERS[8][16] ), .ZN(n607) );
  INV_X1 U1270 ( .A(\REGISTERS[9][16] ), .ZN(n606) );
  OAI221_X1 U1271 ( .B1(n609), .B2(n1187), .C1(n610), .C2(n1188), .A(n1479), 
        .ZN(n1472) );
  AOI22_X1 U1272 ( .A1(n1190), .A2(\REGISTERS[15][16] ), .B1(n1191), .B2(
        \REGISTERS[14][16] ), .ZN(n1479) );
  INV_X1 U1273 ( .A(\REGISTERS[12][16] ), .ZN(n610) );
  INV_X1 U1274 ( .A(\REGISTERS[13][16] ), .ZN(n609) );
  NAND2_X1 U1275 ( .A1(n1480), .A2(n1481), .ZN(N4229) );
  NOR4_X1 U1276 ( .A1(n1482), .A2(n1483), .A3(n1484), .A4(n1485), .ZN(n1481)
         );
  OAI221_X1 U1277 ( .B1(n618), .B2(n1148), .C1(n619), .C2(n1149), .A(n1486), 
        .ZN(n1485) );
  AOI22_X1 U1278 ( .A1(n1151), .A2(\REGISTERS[19][17] ), .B1(n1152), .B2(
        \REGISTERS[18][17] ), .ZN(n1486) );
  INV_X1 U1279 ( .A(\REGISTERS[16][17] ), .ZN(n619) );
  INV_X1 U1280 ( .A(\REGISTERS[17][17] ), .ZN(n618) );
  OAI221_X1 U1281 ( .B1(n621), .B2(n1153), .C1(n622), .C2(n1154), .A(n1487), 
        .ZN(n1484) );
  AOI22_X1 U1282 ( .A1(n1156), .A2(\REGISTERS[23][17] ), .B1(n1157), .B2(
        \REGISTERS[22][17] ), .ZN(n1487) );
  INV_X1 U1283 ( .A(\REGISTERS[20][17] ), .ZN(n622) );
  INV_X1 U1284 ( .A(\REGISTERS[21][17] ), .ZN(n621) );
  OAI221_X1 U1285 ( .B1(n624), .B2(n1158), .C1(n625), .C2(n1159), .A(n1488), 
        .ZN(n1483) );
  AOI22_X1 U1286 ( .A1(n1161), .A2(\REGISTERS[27][17] ), .B1(n1162), .B2(
        \REGISTERS[26][17] ), .ZN(n1488) );
  INV_X1 U1287 ( .A(\REGISTERS[24][17] ), .ZN(n625) );
  INV_X1 U1288 ( .A(\REGISTERS[25][17] ), .ZN(n624) );
  OAI221_X1 U1289 ( .B1(n627), .B2(n1163), .C1(n628), .C2(n1164), .A(n1489), 
        .ZN(n1482) );
  AOI22_X1 U1290 ( .A1(n1166), .A2(\REGISTERS[29][17] ), .B1(n1167), .B2(
        \REGISTERS[28][17] ), .ZN(n1489) );
  INV_X1 U1291 ( .A(\REGISTERS[30][17] ), .ZN(n628) );
  INV_X1 U1292 ( .A(\REGISTERS[31][17] ), .ZN(n627) );
  NOR4_X1 U1293 ( .A1(n1490), .A2(n1491), .A3(n1492), .A4(n1493), .ZN(n1480)
         );
  AOI22_X1 U1295 ( .A1(n1175), .A2(\REGISTERS[3][17] ), .B1(n1176), .B2(
        \REGISTERS[2][17] ), .ZN(n1494) );
  INV_X1 U1296 ( .A(\REGISTERS[1][17] ), .ZN(n634) );
  OAI221_X1 U1297 ( .B1(n637), .B2(n1177), .C1(n638), .C2(n1178), .A(n1495), 
        .ZN(n1492) );
  AOI22_X1 U1298 ( .A1(n1180), .A2(\REGISTERS[7][17] ), .B1(n1181), .B2(
        \REGISTERS[6][17] ), .ZN(n1495) );
  INV_X1 U1299 ( .A(\REGISTERS[4][17] ), .ZN(n638) );
  INV_X1 U1300 ( .A(\REGISTERS[5][17] ), .ZN(n637) );
  OAI221_X1 U1301 ( .B1(n640), .B2(n1182), .C1(n641), .C2(n1183), .A(n1496), 
        .ZN(n1491) );
  AOI22_X1 U1302 ( .A1(n1185), .A2(\REGISTERS[11][17] ), .B1(n1186), .B2(
        \REGISTERS[10][17] ), .ZN(n1496) );
  INV_X1 U1303 ( .A(\REGISTERS[8][17] ), .ZN(n641) );
  INV_X1 U1304 ( .A(\REGISTERS[9][17] ), .ZN(n640) );
  OAI221_X1 U1305 ( .B1(n643), .B2(n1187), .C1(n644), .C2(n1188), .A(n1497), 
        .ZN(n1490) );
  AOI22_X1 U1306 ( .A1(n1190), .A2(\REGISTERS[15][17] ), .B1(n1191), .B2(
        \REGISTERS[14][17] ), .ZN(n1497) );
  INV_X1 U1307 ( .A(\REGISTERS[12][17] ), .ZN(n644) );
  INV_X1 U1308 ( .A(\REGISTERS[13][17] ), .ZN(n643) );
  NAND2_X1 U1309 ( .A1(n1498), .A2(n1499), .ZN(N4228) );
  NOR4_X1 U1310 ( .A1(n1500), .A2(n1501), .A3(n1502), .A4(n1503), .ZN(n1499)
         );
  OAI221_X1 U1311 ( .B1(n652), .B2(n1148), .C1(n653), .C2(n1149), .A(n1504), 
        .ZN(n1503) );
  AOI22_X1 U1312 ( .A1(n1151), .A2(\REGISTERS[19][18] ), .B1(n1152), .B2(
        \REGISTERS[18][18] ), .ZN(n1504) );
  INV_X1 U1313 ( .A(\REGISTERS[16][18] ), .ZN(n653) );
  INV_X1 U1314 ( .A(\REGISTERS[17][18] ), .ZN(n652) );
  OAI221_X1 U1315 ( .B1(n655), .B2(n1153), .C1(n656), .C2(n1154), .A(n1505), 
        .ZN(n1502) );
  AOI22_X1 U1316 ( .A1(n1156), .A2(\REGISTERS[23][18] ), .B1(n1157), .B2(
        \REGISTERS[22][18] ), .ZN(n1505) );
  INV_X1 U1317 ( .A(\REGISTERS[20][18] ), .ZN(n656) );
  INV_X1 U1318 ( .A(\REGISTERS[21][18] ), .ZN(n655) );
  OAI221_X1 U1319 ( .B1(n658), .B2(n1158), .C1(n659), .C2(n1159), .A(n1506), 
        .ZN(n1501) );
  AOI22_X1 U1320 ( .A1(n1161), .A2(\REGISTERS[27][18] ), .B1(n1162), .B2(
        \REGISTERS[26][18] ), .ZN(n1506) );
  INV_X1 U1321 ( .A(\REGISTERS[24][18] ), .ZN(n659) );
  INV_X1 U1322 ( .A(\REGISTERS[25][18] ), .ZN(n658) );
  OAI221_X1 U1323 ( .B1(n661), .B2(n1163), .C1(n662), .C2(n1164), .A(n1507), 
        .ZN(n1500) );
  AOI22_X1 U1324 ( .A1(n1166), .A2(\REGISTERS[29][18] ), .B1(n1167), .B2(
        \REGISTERS[28][18] ), .ZN(n1507) );
  INV_X1 U1325 ( .A(\REGISTERS[30][18] ), .ZN(n662) );
  INV_X1 U1326 ( .A(\REGISTERS[31][18] ), .ZN(n661) );
  NOR4_X1 U1327 ( .A1(n1508), .A2(n1509), .A3(n1510), .A4(n1511), .ZN(n1498)
         );
  AOI22_X1 U1329 ( .A1(n1175), .A2(\REGISTERS[3][18] ), .B1(n1176), .B2(
        \REGISTERS[2][18] ), .ZN(n1512) );
  INV_X1 U1330 ( .A(\REGISTERS[1][18] ), .ZN(n668) );
  OAI221_X1 U1331 ( .B1(n671), .B2(n1177), .C1(n672), .C2(n1178), .A(n1513), 
        .ZN(n1510) );
  AOI22_X1 U1332 ( .A1(n1180), .A2(\REGISTERS[7][18] ), .B1(n1181), .B2(
        \REGISTERS[6][18] ), .ZN(n1513) );
  INV_X1 U1333 ( .A(\REGISTERS[4][18] ), .ZN(n672) );
  INV_X1 U1334 ( .A(\REGISTERS[5][18] ), .ZN(n671) );
  OAI221_X1 U1335 ( .B1(n674), .B2(n1182), .C1(n675), .C2(n1183), .A(n1514), 
        .ZN(n1509) );
  AOI22_X1 U1336 ( .A1(n1185), .A2(\REGISTERS[11][18] ), .B1(n1186), .B2(
        \REGISTERS[10][18] ), .ZN(n1514) );
  INV_X1 U1337 ( .A(\REGISTERS[8][18] ), .ZN(n675) );
  INV_X1 U1338 ( .A(\REGISTERS[9][18] ), .ZN(n674) );
  OAI221_X1 U1339 ( .B1(n677), .B2(n1187), .C1(n678), .C2(n1188), .A(n1515), 
        .ZN(n1508) );
  AOI22_X1 U1340 ( .A1(n1190), .A2(\REGISTERS[15][18] ), .B1(n1191), .B2(
        \REGISTERS[14][18] ), .ZN(n1515) );
  INV_X1 U1341 ( .A(\REGISTERS[12][18] ), .ZN(n678) );
  INV_X1 U1342 ( .A(\REGISTERS[13][18] ), .ZN(n677) );
  NAND2_X1 U1343 ( .A1(n1516), .A2(n1517), .ZN(N4227) );
  NOR4_X1 U1344 ( .A1(n1518), .A2(n1519), .A3(n1520), .A4(n1521), .ZN(n1517)
         );
  OAI221_X1 U1345 ( .B1(n686), .B2(n1148), .C1(n687), .C2(n1149), .A(n1522), 
        .ZN(n1521) );
  AOI22_X1 U1346 ( .A1(n1151), .A2(\REGISTERS[19][19] ), .B1(n1152), .B2(
        \REGISTERS[18][19] ), .ZN(n1522) );
  INV_X1 U1347 ( .A(\REGISTERS[16][19] ), .ZN(n687) );
  INV_X1 U1348 ( .A(\REGISTERS[17][19] ), .ZN(n686) );
  OAI221_X1 U1349 ( .B1(n689), .B2(n1153), .C1(n690), .C2(n1154), .A(n1523), 
        .ZN(n1520) );
  AOI22_X1 U1350 ( .A1(n1156), .A2(\REGISTERS[23][19] ), .B1(n1157), .B2(
        \REGISTERS[22][19] ), .ZN(n1523) );
  INV_X1 U1351 ( .A(\REGISTERS[20][19] ), .ZN(n690) );
  INV_X1 U1352 ( .A(\REGISTERS[21][19] ), .ZN(n689) );
  OAI221_X1 U1353 ( .B1(n692), .B2(n1158), .C1(n693), .C2(n1159), .A(n1524), 
        .ZN(n1519) );
  AOI22_X1 U1354 ( .A1(n1161), .A2(\REGISTERS[27][19] ), .B1(n1162), .B2(
        \REGISTERS[26][19] ), .ZN(n1524) );
  INV_X1 U1355 ( .A(\REGISTERS[24][19] ), .ZN(n693) );
  INV_X1 U1356 ( .A(\REGISTERS[25][19] ), .ZN(n692) );
  OAI221_X1 U1357 ( .B1(n695), .B2(n1163), .C1(n696), .C2(n1164), .A(n1525), 
        .ZN(n1518) );
  AOI22_X1 U1358 ( .A1(n1166), .A2(\REGISTERS[29][19] ), .B1(n1167), .B2(
        \REGISTERS[28][19] ), .ZN(n1525) );
  INV_X1 U1359 ( .A(\REGISTERS[30][19] ), .ZN(n696) );
  INV_X1 U1360 ( .A(\REGISTERS[31][19] ), .ZN(n695) );
  NOR4_X1 U1361 ( .A1(n1526), .A2(n1527), .A3(n1528), .A4(n1529), .ZN(n1516)
         );
  AOI22_X1 U1363 ( .A1(n1175), .A2(\REGISTERS[3][19] ), .B1(n1176), .B2(
        \REGISTERS[2][19] ), .ZN(n1530) );
  INV_X1 U1364 ( .A(\REGISTERS[1][19] ), .ZN(n702) );
  OAI221_X1 U1365 ( .B1(n705), .B2(n1177), .C1(n706), .C2(n1178), .A(n1531), 
        .ZN(n1528) );
  AOI22_X1 U1366 ( .A1(n1180), .A2(\REGISTERS[7][19] ), .B1(n1181), .B2(
        \REGISTERS[6][19] ), .ZN(n1531) );
  INV_X1 U1367 ( .A(\REGISTERS[4][19] ), .ZN(n706) );
  INV_X1 U1368 ( .A(\REGISTERS[5][19] ), .ZN(n705) );
  OAI221_X1 U1369 ( .B1(n708), .B2(n1182), .C1(n709), .C2(n1183), .A(n1532), 
        .ZN(n1527) );
  AOI22_X1 U1370 ( .A1(n1185), .A2(\REGISTERS[11][19] ), .B1(n1186), .B2(
        \REGISTERS[10][19] ), .ZN(n1532) );
  INV_X1 U1371 ( .A(\REGISTERS[8][19] ), .ZN(n709) );
  INV_X1 U1372 ( .A(\REGISTERS[9][19] ), .ZN(n708) );
  OAI221_X1 U1373 ( .B1(n711), .B2(n1187), .C1(n712), .C2(n1188), .A(n1533), 
        .ZN(n1526) );
  AOI22_X1 U1374 ( .A1(n1190), .A2(\REGISTERS[15][19] ), .B1(n1191), .B2(
        \REGISTERS[14][19] ), .ZN(n1533) );
  INV_X1 U1375 ( .A(\REGISTERS[12][19] ), .ZN(n712) );
  INV_X1 U1376 ( .A(\REGISTERS[13][19] ), .ZN(n711) );
  NAND2_X1 U1377 ( .A1(n1534), .A2(n1535), .ZN(N4226) );
  NOR4_X1 U1378 ( .A1(n1536), .A2(n1537), .A3(n1538), .A4(n1539), .ZN(n1535)
         );
  OAI221_X1 U1379 ( .B1(n720), .B2(n1148), .C1(n721), .C2(n1149), .A(n1540), 
        .ZN(n1539) );
  AOI22_X1 U1380 ( .A1(n1151), .A2(\REGISTERS[19][20] ), .B1(n1152), .B2(
        \REGISTERS[18][20] ), .ZN(n1540) );
  INV_X1 U1381 ( .A(\REGISTERS[16][20] ), .ZN(n721) );
  INV_X1 U1382 ( .A(\REGISTERS[17][20] ), .ZN(n720) );
  OAI221_X1 U1383 ( .B1(n723), .B2(n1153), .C1(n724), .C2(n1154), .A(n1541), 
        .ZN(n1538) );
  AOI22_X1 U1384 ( .A1(n1156), .A2(\REGISTERS[23][20] ), .B1(n1157), .B2(
        \REGISTERS[22][20] ), .ZN(n1541) );
  INV_X1 U1385 ( .A(\REGISTERS[20][20] ), .ZN(n724) );
  INV_X1 U1386 ( .A(\REGISTERS[21][20] ), .ZN(n723) );
  OAI221_X1 U1387 ( .B1(n726), .B2(n1158), .C1(n727), .C2(n1159), .A(n1542), 
        .ZN(n1537) );
  AOI22_X1 U1388 ( .A1(n1161), .A2(\REGISTERS[27][20] ), .B1(n1162), .B2(
        \REGISTERS[26][20] ), .ZN(n1542) );
  INV_X1 U1389 ( .A(\REGISTERS[24][20] ), .ZN(n727) );
  INV_X1 U1390 ( .A(\REGISTERS[25][20] ), .ZN(n726) );
  OAI221_X1 U1391 ( .B1(n729), .B2(n1163), .C1(n730), .C2(n1164), .A(n1543), 
        .ZN(n1536) );
  AOI22_X1 U1392 ( .A1(n1166), .A2(\REGISTERS[29][20] ), .B1(n1167), .B2(
        \REGISTERS[28][20] ), .ZN(n1543) );
  INV_X1 U1393 ( .A(\REGISTERS[30][20] ), .ZN(n730) );
  INV_X1 U1394 ( .A(\REGISTERS[31][20] ), .ZN(n729) );
  NOR4_X1 U1395 ( .A1(n1544), .A2(n1545), .A3(n1546), .A4(n1547), .ZN(n1534)
         );
  AOI22_X1 U1397 ( .A1(n1175), .A2(\REGISTERS[3][20] ), .B1(n1176), .B2(
        \REGISTERS[2][20] ), .ZN(n1548) );
  INV_X1 U1398 ( .A(\REGISTERS[1][20] ), .ZN(n736) );
  OAI221_X1 U1399 ( .B1(n739), .B2(n1177), .C1(n740), .C2(n1178), .A(n1549), 
        .ZN(n1546) );
  AOI22_X1 U1400 ( .A1(n1180), .A2(\REGISTERS[7][20] ), .B1(n1181), .B2(
        \REGISTERS[6][20] ), .ZN(n1549) );
  INV_X1 U1401 ( .A(\REGISTERS[4][20] ), .ZN(n740) );
  INV_X1 U1402 ( .A(\REGISTERS[5][20] ), .ZN(n739) );
  OAI221_X1 U1403 ( .B1(n742), .B2(n1182), .C1(n743), .C2(n1183), .A(n1550), 
        .ZN(n1545) );
  AOI22_X1 U1404 ( .A1(n1185), .A2(\REGISTERS[11][20] ), .B1(n1186), .B2(
        \REGISTERS[10][20] ), .ZN(n1550) );
  INV_X1 U1405 ( .A(\REGISTERS[8][20] ), .ZN(n743) );
  INV_X1 U1406 ( .A(\REGISTERS[9][20] ), .ZN(n742) );
  OAI221_X1 U1407 ( .B1(n745), .B2(n1187), .C1(n746), .C2(n1188), .A(n1551), 
        .ZN(n1544) );
  AOI22_X1 U1408 ( .A1(n1190), .A2(\REGISTERS[15][20] ), .B1(n1191), .B2(
        \REGISTERS[14][20] ), .ZN(n1551) );
  INV_X1 U1409 ( .A(\REGISTERS[12][20] ), .ZN(n746) );
  INV_X1 U1410 ( .A(\REGISTERS[13][20] ), .ZN(n745) );
  NAND2_X1 U1411 ( .A1(n1552), .A2(n1553), .ZN(N4225) );
  NOR4_X1 U1412 ( .A1(n1554), .A2(n1555), .A3(n1556), .A4(n1557), .ZN(n1553)
         );
  OAI221_X1 U1413 ( .B1(n754), .B2(n1148), .C1(n755), .C2(n1149), .A(n1558), 
        .ZN(n1557) );
  AOI22_X1 U1414 ( .A1(n1151), .A2(\REGISTERS[19][21] ), .B1(n1152), .B2(
        \REGISTERS[18][21] ), .ZN(n1558) );
  INV_X1 U1415 ( .A(\REGISTERS[16][21] ), .ZN(n755) );
  INV_X1 U1416 ( .A(\REGISTERS[17][21] ), .ZN(n754) );
  OAI221_X1 U1417 ( .B1(n757), .B2(n1153), .C1(n758), .C2(n1154), .A(n1559), 
        .ZN(n1556) );
  AOI22_X1 U1418 ( .A1(n1156), .A2(\REGISTERS[23][21] ), .B1(n1157), .B2(
        \REGISTERS[22][21] ), .ZN(n1559) );
  INV_X1 U1419 ( .A(\REGISTERS[20][21] ), .ZN(n758) );
  INV_X1 U1420 ( .A(\REGISTERS[21][21] ), .ZN(n757) );
  OAI221_X1 U1421 ( .B1(n760), .B2(n1158), .C1(n761), .C2(n1159), .A(n1560), 
        .ZN(n1555) );
  AOI22_X1 U1422 ( .A1(n1161), .A2(\REGISTERS[27][21] ), .B1(n1162), .B2(
        \REGISTERS[26][21] ), .ZN(n1560) );
  INV_X1 U1423 ( .A(\REGISTERS[24][21] ), .ZN(n761) );
  INV_X1 U1424 ( .A(\REGISTERS[25][21] ), .ZN(n760) );
  OAI221_X1 U1425 ( .B1(n763), .B2(n1163), .C1(n764), .C2(n1164), .A(n1561), 
        .ZN(n1554) );
  AOI22_X1 U1426 ( .A1(n1166), .A2(\REGISTERS[29][21] ), .B1(n1167), .B2(
        \REGISTERS[28][21] ), .ZN(n1561) );
  INV_X1 U1427 ( .A(\REGISTERS[30][21] ), .ZN(n764) );
  INV_X1 U1428 ( .A(\REGISTERS[31][21] ), .ZN(n763) );
  NOR4_X1 U1429 ( .A1(n1562), .A2(n1563), .A3(n1564), .A4(n1565), .ZN(n1552)
         );
  AOI22_X1 U1431 ( .A1(n1175), .A2(\REGISTERS[3][21] ), .B1(n1176), .B2(
        \REGISTERS[2][21] ), .ZN(n1566) );
  INV_X1 U1432 ( .A(\REGISTERS[1][21] ), .ZN(n770) );
  OAI221_X1 U1433 ( .B1(n773), .B2(n1177), .C1(n774), .C2(n1178), .A(n1567), 
        .ZN(n1564) );
  AOI22_X1 U1434 ( .A1(n1180), .A2(\REGISTERS[7][21] ), .B1(n1181), .B2(
        \REGISTERS[6][21] ), .ZN(n1567) );
  INV_X1 U1435 ( .A(\REGISTERS[4][21] ), .ZN(n774) );
  INV_X1 U1436 ( .A(\REGISTERS[5][21] ), .ZN(n773) );
  OAI221_X1 U1437 ( .B1(n776), .B2(n1182), .C1(n777), .C2(n1183), .A(n1568), 
        .ZN(n1563) );
  AOI22_X1 U1438 ( .A1(n1185), .A2(\REGISTERS[11][21] ), .B1(n1186), .B2(
        \REGISTERS[10][21] ), .ZN(n1568) );
  INV_X1 U1439 ( .A(\REGISTERS[8][21] ), .ZN(n777) );
  INV_X1 U1440 ( .A(\REGISTERS[9][21] ), .ZN(n776) );
  OAI221_X1 U1441 ( .B1(n779), .B2(n1187), .C1(n780), .C2(n1188), .A(n1569), 
        .ZN(n1562) );
  AOI22_X1 U1442 ( .A1(n1190), .A2(\REGISTERS[15][21] ), .B1(n1191), .B2(
        \REGISTERS[14][21] ), .ZN(n1569) );
  INV_X1 U1443 ( .A(\REGISTERS[12][21] ), .ZN(n780) );
  INV_X1 U1444 ( .A(\REGISTERS[13][21] ), .ZN(n779) );
  NAND2_X1 U1445 ( .A1(n1570), .A2(n1571), .ZN(N4224) );
  NOR4_X1 U1446 ( .A1(n1572), .A2(n1573), .A3(n1574), .A4(n1575), .ZN(n1571)
         );
  OAI221_X1 U1447 ( .B1(n788), .B2(n1148), .C1(n789), .C2(n1149), .A(n1576), 
        .ZN(n1575) );
  AOI22_X1 U1448 ( .A1(n1151), .A2(\REGISTERS[19][22] ), .B1(n1152), .B2(
        \REGISTERS[18][22] ), .ZN(n1576) );
  INV_X1 U1449 ( .A(\REGISTERS[16][22] ), .ZN(n789) );
  INV_X1 U1450 ( .A(\REGISTERS[17][22] ), .ZN(n788) );
  OAI221_X1 U1451 ( .B1(n791), .B2(n1153), .C1(n792), .C2(n1154), .A(n1577), 
        .ZN(n1574) );
  AOI22_X1 U1452 ( .A1(n1156), .A2(\REGISTERS[23][22] ), .B1(n1157), .B2(
        \REGISTERS[22][22] ), .ZN(n1577) );
  INV_X1 U1453 ( .A(\REGISTERS[20][22] ), .ZN(n792) );
  INV_X1 U1454 ( .A(\REGISTERS[21][22] ), .ZN(n791) );
  OAI221_X1 U1455 ( .B1(n794), .B2(n1158), .C1(n795), .C2(n1159), .A(n1578), 
        .ZN(n1573) );
  AOI22_X1 U1456 ( .A1(n1161), .A2(\REGISTERS[27][22] ), .B1(n1162), .B2(
        \REGISTERS[26][22] ), .ZN(n1578) );
  INV_X1 U1457 ( .A(\REGISTERS[24][22] ), .ZN(n795) );
  INV_X1 U1458 ( .A(\REGISTERS[25][22] ), .ZN(n794) );
  OAI221_X1 U1459 ( .B1(n797), .B2(n1163), .C1(n798), .C2(n1164), .A(n1579), 
        .ZN(n1572) );
  AOI22_X1 U1460 ( .A1(n1166), .A2(\REGISTERS[29][22] ), .B1(n1167), .B2(
        \REGISTERS[28][22] ), .ZN(n1579) );
  INV_X1 U1461 ( .A(\REGISTERS[30][22] ), .ZN(n798) );
  INV_X1 U1462 ( .A(\REGISTERS[31][22] ), .ZN(n797) );
  NOR4_X1 U1463 ( .A1(n1580), .A2(n1581), .A3(n1582), .A4(n1583), .ZN(n1570)
         );
  AOI22_X1 U1465 ( .A1(n1175), .A2(\REGISTERS[3][22] ), .B1(n1176), .B2(
        \REGISTERS[2][22] ), .ZN(n1584) );
  INV_X1 U1466 ( .A(\REGISTERS[1][22] ), .ZN(n804) );
  OAI221_X1 U1467 ( .B1(n807), .B2(n1177), .C1(n808), .C2(n1178), .A(n1585), 
        .ZN(n1582) );
  AOI22_X1 U1468 ( .A1(n1180), .A2(\REGISTERS[7][22] ), .B1(n1181), .B2(
        \REGISTERS[6][22] ), .ZN(n1585) );
  INV_X1 U1469 ( .A(\REGISTERS[4][22] ), .ZN(n808) );
  INV_X1 U1470 ( .A(\REGISTERS[5][22] ), .ZN(n807) );
  OAI221_X1 U1471 ( .B1(n810), .B2(n1182), .C1(n811), .C2(n1183), .A(n1586), 
        .ZN(n1581) );
  AOI22_X1 U1472 ( .A1(n1185), .A2(\REGISTERS[11][22] ), .B1(n1186), .B2(
        \REGISTERS[10][22] ), .ZN(n1586) );
  INV_X1 U1473 ( .A(\REGISTERS[8][22] ), .ZN(n811) );
  INV_X1 U1474 ( .A(\REGISTERS[9][22] ), .ZN(n810) );
  OAI221_X1 U1475 ( .B1(n813), .B2(n1187), .C1(n814), .C2(n1188), .A(n1587), 
        .ZN(n1580) );
  AOI22_X1 U1476 ( .A1(n1190), .A2(\REGISTERS[15][22] ), .B1(n1191), .B2(
        \REGISTERS[14][22] ), .ZN(n1587) );
  INV_X1 U1477 ( .A(\REGISTERS[12][22] ), .ZN(n814) );
  INV_X1 U1478 ( .A(\REGISTERS[13][22] ), .ZN(n813) );
  NAND2_X1 U1479 ( .A1(n1588), .A2(n1589), .ZN(N4223) );
  NOR4_X1 U1480 ( .A1(n1590), .A2(n1591), .A3(n1592), .A4(n1593), .ZN(n1589)
         );
  OAI221_X1 U1481 ( .B1(n822), .B2(n1148), .C1(n823), .C2(n1149), .A(n1594), 
        .ZN(n1593) );
  AOI22_X1 U1482 ( .A1(n1151), .A2(\REGISTERS[19][23] ), .B1(n1152), .B2(
        \REGISTERS[18][23] ), .ZN(n1594) );
  INV_X1 U1483 ( .A(\REGISTERS[16][23] ), .ZN(n823) );
  INV_X1 U1484 ( .A(\REGISTERS[17][23] ), .ZN(n822) );
  OAI221_X1 U1485 ( .B1(n825), .B2(n1153), .C1(n826), .C2(n1154), .A(n1595), 
        .ZN(n1592) );
  AOI22_X1 U1486 ( .A1(n1156), .A2(\REGISTERS[23][23] ), .B1(n1157), .B2(
        \REGISTERS[22][23] ), .ZN(n1595) );
  INV_X1 U1487 ( .A(\REGISTERS[20][23] ), .ZN(n826) );
  INV_X1 U1488 ( .A(\REGISTERS[21][23] ), .ZN(n825) );
  OAI221_X1 U1489 ( .B1(n828), .B2(n1158), .C1(n829), .C2(n1159), .A(n1596), 
        .ZN(n1591) );
  AOI22_X1 U1490 ( .A1(n1161), .A2(\REGISTERS[27][23] ), .B1(n1162), .B2(
        \REGISTERS[26][23] ), .ZN(n1596) );
  INV_X1 U1491 ( .A(\REGISTERS[24][23] ), .ZN(n829) );
  INV_X1 U1492 ( .A(\REGISTERS[25][23] ), .ZN(n828) );
  OAI221_X1 U1493 ( .B1(n831), .B2(n1163), .C1(n832), .C2(n1164), .A(n1597), 
        .ZN(n1590) );
  AOI22_X1 U1494 ( .A1(n1166), .A2(\REGISTERS[29][23] ), .B1(n1167), .B2(
        \REGISTERS[28][23] ), .ZN(n1597) );
  INV_X1 U1495 ( .A(\REGISTERS[30][23] ), .ZN(n832) );
  INV_X1 U1496 ( .A(\REGISTERS[31][23] ), .ZN(n831) );
  NOR4_X1 U1497 ( .A1(n1598), .A2(n1599), .A3(n1600), .A4(n1601), .ZN(n1588)
         );
  AOI22_X1 U1499 ( .A1(n1175), .A2(\REGISTERS[3][23] ), .B1(n1176), .B2(
        \REGISTERS[2][23] ), .ZN(n1602) );
  INV_X1 U1500 ( .A(\REGISTERS[1][23] ), .ZN(n838) );
  OAI221_X1 U1501 ( .B1(n841), .B2(n1177), .C1(n842), .C2(n1178), .A(n1603), 
        .ZN(n1600) );
  AOI22_X1 U1502 ( .A1(n1180), .A2(\REGISTERS[7][23] ), .B1(n1181), .B2(
        \REGISTERS[6][23] ), .ZN(n1603) );
  INV_X1 U1503 ( .A(\REGISTERS[4][23] ), .ZN(n842) );
  INV_X1 U1504 ( .A(\REGISTERS[5][23] ), .ZN(n841) );
  OAI221_X1 U1505 ( .B1(n844), .B2(n1182), .C1(n845), .C2(n1183), .A(n1604), 
        .ZN(n1599) );
  AOI22_X1 U1506 ( .A1(n1185), .A2(\REGISTERS[11][23] ), .B1(n1186), .B2(
        \REGISTERS[10][23] ), .ZN(n1604) );
  INV_X1 U1507 ( .A(\REGISTERS[8][23] ), .ZN(n845) );
  INV_X1 U1508 ( .A(\REGISTERS[9][23] ), .ZN(n844) );
  OAI221_X1 U1509 ( .B1(n847), .B2(n1187), .C1(n848), .C2(n1188), .A(n1605), 
        .ZN(n1598) );
  AOI22_X1 U1510 ( .A1(n1190), .A2(\REGISTERS[15][23] ), .B1(n1191), .B2(
        \REGISTERS[14][23] ), .ZN(n1605) );
  INV_X1 U1511 ( .A(\REGISTERS[12][23] ), .ZN(n848) );
  INV_X1 U1512 ( .A(\REGISTERS[13][23] ), .ZN(n847) );
  NAND2_X1 U1513 ( .A1(n1606), .A2(n1607), .ZN(N4222) );
  NOR4_X1 U1514 ( .A1(n1608), .A2(n1609), .A3(n1610), .A4(n1611), .ZN(n1607)
         );
  OAI221_X1 U1515 ( .B1(n856), .B2(n1148), .C1(n857), .C2(n1149), .A(n1612), 
        .ZN(n1611) );
  AOI22_X1 U1516 ( .A1(n1151), .A2(\REGISTERS[19][24] ), .B1(n1152), .B2(
        \REGISTERS[18][24] ), .ZN(n1612) );
  INV_X1 U1517 ( .A(\REGISTERS[16][24] ), .ZN(n857) );
  INV_X1 U1518 ( .A(\REGISTERS[17][24] ), .ZN(n856) );
  OAI221_X1 U1519 ( .B1(n859), .B2(n1153), .C1(n860), .C2(n1154), .A(n1613), 
        .ZN(n1610) );
  AOI22_X1 U1520 ( .A1(n1156), .A2(\REGISTERS[23][24] ), .B1(n1157), .B2(
        \REGISTERS[22][24] ), .ZN(n1613) );
  INV_X1 U1521 ( .A(\REGISTERS[20][24] ), .ZN(n860) );
  INV_X1 U1522 ( .A(\REGISTERS[21][24] ), .ZN(n859) );
  OAI221_X1 U1523 ( .B1(n862), .B2(n1158), .C1(n863), .C2(n1159), .A(n1614), 
        .ZN(n1609) );
  AOI22_X1 U1524 ( .A1(n1161), .A2(\REGISTERS[27][24] ), .B1(n1162), .B2(
        \REGISTERS[26][24] ), .ZN(n1614) );
  INV_X1 U1525 ( .A(\REGISTERS[24][24] ), .ZN(n863) );
  INV_X1 U1526 ( .A(\REGISTERS[25][24] ), .ZN(n862) );
  OAI221_X1 U1527 ( .B1(n865), .B2(n1163), .C1(n866), .C2(n1164), .A(n1615), 
        .ZN(n1608) );
  AOI22_X1 U1528 ( .A1(n1166), .A2(\REGISTERS[29][24] ), .B1(n1167), .B2(
        \REGISTERS[28][24] ), .ZN(n1615) );
  INV_X1 U1529 ( .A(\REGISTERS[30][24] ), .ZN(n866) );
  INV_X1 U1530 ( .A(\REGISTERS[31][24] ), .ZN(n865) );
  NOR4_X1 U1531 ( .A1(n1616), .A2(n1617), .A3(n1618), .A4(n1619), .ZN(n1606)
         );
  AOI22_X1 U1533 ( .A1(n1175), .A2(\REGISTERS[3][24] ), .B1(n1176), .B2(
        \REGISTERS[2][24] ), .ZN(n1620) );
  INV_X1 U1534 ( .A(\REGISTERS[1][24] ), .ZN(n872) );
  OAI221_X1 U1535 ( .B1(n875), .B2(n1177), .C1(n876), .C2(n1178), .A(n1621), 
        .ZN(n1618) );
  AOI22_X1 U1536 ( .A1(n1180), .A2(\REGISTERS[7][24] ), .B1(n1181), .B2(
        \REGISTERS[6][24] ), .ZN(n1621) );
  INV_X1 U1537 ( .A(\REGISTERS[4][24] ), .ZN(n876) );
  INV_X1 U1538 ( .A(\REGISTERS[5][24] ), .ZN(n875) );
  OAI221_X1 U1539 ( .B1(n878), .B2(n1182), .C1(n879), .C2(n1183), .A(n1622), 
        .ZN(n1617) );
  AOI22_X1 U1540 ( .A1(n1185), .A2(\REGISTERS[11][24] ), .B1(n1186), .B2(
        \REGISTERS[10][24] ), .ZN(n1622) );
  INV_X1 U1541 ( .A(\REGISTERS[8][24] ), .ZN(n879) );
  INV_X1 U1542 ( .A(\REGISTERS[9][24] ), .ZN(n878) );
  OAI221_X1 U1543 ( .B1(n881), .B2(n1187), .C1(n882), .C2(n1188), .A(n1623), 
        .ZN(n1616) );
  AOI22_X1 U1544 ( .A1(n1190), .A2(\REGISTERS[15][24] ), .B1(n1191), .B2(
        \REGISTERS[14][24] ), .ZN(n1623) );
  INV_X1 U1545 ( .A(\REGISTERS[12][24] ), .ZN(n882) );
  INV_X1 U1546 ( .A(\REGISTERS[13][24] ), .ZN(n881) );
  NAND2_X1 U1547 ( .A1(n1624), .A2(n1625), .ZN(N4221) );
  NOR4_X1 U1548 ( .A1(n1626), .A2(n1627), .A3(n1628), .A4(n1629), .ZN(n1625)
         );
  OAI221_X1 U1549 ( .B1(n890), .B2(n1148), .C1(n891), .C2(n1149), .A(n1630), 
        .ZN(n1629) );
  AOI22_X1 U1550 ( .A1(n1151), .A2(\REGISTERS[19][25] ), .B1(n1152), .B2(
        \REGISTERS[18][25] ), .ZN(n1630) );
  INV_X1 U1551 ( .A(\REGISTERS[16][25] ), .ZN(n891) );
  INV_X1 U1552 ( .A(\REGISTERS[17][25] ), .ZN(n890) );
  OAI221_X1 U1553 ( .B1(n893), .B2(n1153), .C1(n894), .C2(n1154), .A(n1631), 
        .ZN(n1628) );
  AOI22_X1 U1554 ( .A1(n1156), .A2(\REGISTERS[23][25] ), .B1(n1157), .B2(
        \REGISTERS[22][25] ), .ZN(n1631) );
  INV_X1 U1555 ( .A(\REGISTERS[20][25] ), .ZN(n894) );
  INV_X1 U1556 ( .A(\REGISTERS[21][25] ), .ZN(n893) );
  OAI221_X1 U1557 ( .B1(n896), .B2(n1158), .C1(n897), .C2(n1159), .A(n1632), 
        .ZN(n1627) );
  AOI22_X1 U1558 ( .A1(n1161), .A2(\REGISTERS[27][25] ), .B1(n1162), .B2(
        \REGISTERS[26][25] ), .ZN(n1632) );
  INV_X1 U1559 ( .A(\REGISTERS[24][25] ), .ZN(n897) );
  INV_X1 U1560 ( .A(\REGISTERS[25][25] ), .ZN(n896) );
  OAI221_X1 U1561 ( .B1(n899), .B2(n1163), .C1(n900), .C2(n1164), .A(n1633), 
        .ZN(n1626) );
  AOI22_X1 U1562 ( .A1(n1166), .A2(\REGISTERS[29][25] ), .B1(n1167), .B2(
        \REGISTERS[28][25] ), .ZN(n1633) );
  INV_X1 U1563 ( .A(\REGISTERS[30][25] ), .ZN(n900) );
  INV_X1 U1564 ( .A(\REGISTERS[31][25] ), .ZN(n899) );
  NOR4_X1 U1565 ( .A1(n1634), .A2(n1635), .A3(n1636), .A4(n1637), .ZN(n1624)
         );
  AOI22_X1 U1567 ( .A1(n1175), .A2(\REGISTERS[3][25] ), .B1(n1176), .B2(
        \REGISTERS[2][25] ), .ZN(n1638) );
  INV_X1 U1568 ( .A(\REGISTERS[1][25] ), .ZN(n906) );
  OAI221_X1 U1569 ( .B1(n909), .B2(n1177), .C1(n910), .C2(n1178), .A(n1639), 
        .ZN(n1636) );
  AOI22_X1 U1570 ( .A1(n1180), .A2(\REGISTERS[7][25] ), .B1(n1181), .B2(
        \REGISTERS[6][25] ), .ZN(n1639) );
  INV_X1 U1571 ( .A(\REGISTERS[4][25] ), .ZN(n910) );
  INV_X1 U1572 ( .A(\REGISTERS[5][25] ), .ZN(n909) );
  OAI221_X1 U1573 ( .B1(n912), .B2(n1182), .C1(n913), .C2(n1183), .A(n1640), 
        .ZN(n1635) );
  AOI22_X1 U1574 ( .A1(n1185), .A2(\REGISTERS[11][25] ), .B1(n1186), .B2(
        \REGISTERS[10][25] ), .ZN(n1640) );
  INV_X1 U1575 ( .A(\REGISTERS[8][25] ), .ZN(n913) );
  INV_X1 U1576 ( .A(\REGISTERS[9][25] ), .ZN(n912) );
  OAI221_X1 U1577 ( .B1(n915), .B2(n1187), .C1(n916), .C2(n1188), .A(n1641), 
        .ZN(n1634) );
  AOI22_X1 U1578 ( .A1(n1190), .A2(\REGISTERS[15][25] ), .B1(n1191), .B2(
        \REGISTERS[14][25] ), .ZN(n1641) );
  INV_X1 U1579 ( .A(\REGISTERS[12][25] ), .ZN(n916) );
  INV_X1 U1580 ( .A(\REGISTERS[13][25] ), .ZN(n915) );
  NAND2_X1 U1581 ( .A1(n1642), .A2(n1643), .ZN(N4220) );
  NOR4_X1 U1582 ( .A1(n1644), .A2(n1645), .A3(n1646), .A4(n1647), .ZN(n1643)
         );
  OAI221_X1 U1583 ( .B1(n924), .B2(n1148), .C1(n925), .C2(n1149), .A(n1648), 
        .ZN(n1647) );
  AOI22_X1 U1584 ( .A1(n1151), .A2(\REGISTERS[19][26] ), .B1(n1152), .B2(
        \REGISTERS[18][26] ), .ZN(n1648) );
  INV_X1 U1585 ( .A(\REGISTERS[16][26] ), .ZN(n925) );
  INV_X1 U1586 ( .A(\REGISTERS[17][26] ), .ZN(n924) );
  OAI221_X1 U1587 ( .B1(n927), .B2(n1153), .C1(n928), .C2(n1154), .A(n1649), 
        .ZN(n1646) );
  AOI22_X1 U1588 ( .A1(n1156), .A2(\REGISTERS[23][26] ), .B1(n1157), .B2(
        \REGISTERS[22][26] ), .ZN(n1649) );
  INV_X1 U1589 ( .A(\REGISTERS[20][26] ), .ZN(n928) );
  INV_X1 U1590 ( .A(\REGISTERS[21][26] ), .ZN(n927) );
  OAI221_X1 U1591 ( .B1(n930), .B2(n1158), .C1(n931), .C2(n1159), .A(n1650), 
        .ZN(n1645) );
  AOI22_X1 U1592 ( .A1(n1161), .A2(\REGISTERS[27][26] ), .B1(n1162), .B2(
        \REGISTERS[26][26] ), .ZN(n1650) );
  INV_X1 U1593 ( .A(\REGISTERS[24][26] ), .ZN(n931) );
  INV_X1 U1594 ( .A(\REGISTERS[25][26] ), .ZN(n930) );
  OAI221_X1 U1595 ( .B1(n933), .B2(n1163), .C1(n934), .C2(n1164), .A(n1651), 
        .ZN(n1644) );
  AOI22_X1 U1596 ( .A1(n1166), .A2(\REGISTERS[29][26] ), .B1(n1167), .B2(
        \REGISTERS[28][26] ), .ZN(n1651) );
  INV_X1 U1597 ( .A(\REGISTERS[30][26] ), .ZN(n934) );
  INV_X1 U1598 ( .A(\REGISTERS[31][26] ), .ZN(n933) );
  NOR4_X1 U1599 ( .A1(n1652), .A2(n1653), .A3(n1654), .A4(n1655), .ZN(n1642)
         );
  AOI22_X1 U1601 ( .A1(n1175), .A2(\REGISTERS[3][26] ), .B1(n1176), .B2(
        \REGISTERS[2][26] ), .ZN(n1656) );
  INV_X1 U1602 ( .A(\REGISTERS[1][26] ), .ZN(n940) );
  OAI221_X1 U1603 ( .B1(n943), .B2(n1177), .C1(n944), .C2(n1178), .A(n1657), 
        .ZN(n1654) );
  AOI22_X1 U1604 ( .A1(n1180), .A2(\REGISTERS[7][26] ), .B1(n1181), .B2(
        \REGISTERS[6][26] ), .ZN(n1657) );
  INV_X1 U1605 ( .A(\REGISTERS[4][26] ), .ZN(n944) );
  INV_X1 U1606 ( .A(\REGISTERS[5][26] ), .ZN(n943) );
  OAI221_X1 U1607 ( .B1(n946), .B2(n1182), .C1(n947), .C2(n1183), .A(n1658), 
        .ZN(n1653) );
  AOI22_X1 U1608 ( .A1(n1185), .A2(\REGISTERS[11][26] ), .B1(n1186), .B2(
        \REGISTERS[10][26] ), .ZN(n1658) );
  INV_X1 U1609 ( .A(\REGISTERS[8][26] ), .ZN(n947) );
  INV_X1 U1610 ( .A(\REGISTERS[9][26] ), .ZN(n946) );
  OAI221_X1 U1611 ( .B1(n949), .B2(n1187), .C1(n950), .C2(n1188), .A(n1659), 
        .ZN(n1652) );
  AOI22_X1 U1612 ( .A1(n1190), .A2(\REGISTERS[15][26] ), .B1(n1191), .B2(
        \REGISTERS[14][26] ), .ZN(n1659) );
  INV_X1 U1613 ( .A(\REGISTERS[12][26] ), .ZN(n950) );
  INV_X1 U1614 ( .A(\REGISTERS[13][26] ), .ZN(n949) );
  NAND2_X1 U1615 ( .A1(n1660), .A2(n1661), .ZN(N4219) );
  NOR4_X1 U1616 ( .A1(n1662), .A2(n1663), .A3(n1664), .A4(n1665), .ZN(n1661)
         );
  OAI221_X1 U1617 ( .B1(n958), .B2(n1148), .C1(n959), .C2(n1149), .A(n1666), 
        .ZN(n1665) );
  AOI22_X1 U1618 ( .A1(n1151), .A2(\REGISTERS[19][27] ), .B1(n1152), .B2(
        \REGISTERS[18][27] ), .ZN(n1666) );
  INV_X1 U1619 ( .A(\REGISTERS[16][27] ), .ZN(n959) );
  INV_X1 U1620 ( .A(\REGISTERS[17][27] ), .ZN(n958) );
  OAI221_X1 U1621 ( .B1(n961), .B2(n1153), .C1(n962), .C2(n1154), .A(n1667), 
        .ZN(n1664) );
  AOI22_X1 U1622 ( .A1(n1156), .A2(\REGISTERS[23][27] ), .B1(n1157), .B2(
        \REGISTERS[22][27] ), .ZN(n1667) );
  INV_X1 U1623 ( .A(\REGISTERS[20][27] ), .ZN(n962) );
  INV_X1 U1624 ( .A(\REGISTERS[21][27] ), .ZN(n961) );
  OAI221_X1 U1625 ( .B1(n964), .B2(n1158), .C1(n965), .C2(n1159), .A(n1668), 
        .ZN(n1663) );
  AOI22_X1 U1626 ( .A1(n1161), .A2(\REGISTERS[27][27] ), .B1(n1162), .B2(
        \REGISTERS[26][27] ), .ZN(n1668) );
  INV_X1 U1627 ( .A(\REGISTERS[24][27] ), .ZN(n965) );
  INV_X1 U1628 ( .A(\REGISTERS[25][27] ), .ZN(n964) );
  OAI221_X1 U1629 ( .B1(n967), .B2(n1163), .C1(n968), .C2(n1164), .A(n1669), 
        .ZN(n1662) );
  AOI22_X1 U1630 ( .A1(n1166), .A2(\REGISTERS[29][27] ), .B1(n1167), .B2(
        \REGISTERS[28][27] ), .ZN(n1669) );
  INV_X1 U1631 ( .A(\REGISTERS[30][27] ), .ZN(n968) );
  INV_X1 U1632 ( .A(\REGISTERS[31][27] ), .ZN(n967) );
  NOR4_X1 U1633 ( .A1(n1670), .A2(n1671), .A3(n1672), .A4(n1673), .ZN(n1660)
         );
  AOI22_X1 U1635 ( .A1(n1175), .A2(\REGISTERS[3][27] ), .B1(n1176), .B2(
        \REGISTERS[2][27] ), .ZN(n1674) );
  INV_X1 U1636 ( .A(\REGISTERS[1][27] ), .ZN(n974) );
  OAI221_X1 U1637 ( .B1(n977), .B2(n1177), .C1(n978), .C2(n1178), .A(n1675), 
        .ZN(n1672) );
  AOI22_X1 U1638 ( .A1(n1180), .A2(\REGISTERS[7][27] ), .B1(n1181), .B2(
        \REGISTERS[6][27] ), .ZN(n1675) );
  INV_X1 U1639 ( .A(\REGISTERS[4][27] ), .ZN(n978) );
  INV_X1 U1640 ( .A(\REGISTERS[5][27] ), .ZN(n977) );
  OAI221_X1 U1641 ( .B1(n980), .B2(n1182), .C1(n981), .C2(n1183), .A(n1676), 
        .ZN(n1671) );
  AOI22_X1 U1642 ( .A1(n1185), .A2(\REGISTERS[11][27] ), .B1(n1186), .B2(
        \REGISTERS[10][27] ), .ZN(n1676) );
  INV_X1 U1643 ( .A(\REGISTERS[8][27] ), .ZN(n981) );
  INV_X1 U1644 ( .A(\REGISTERS[9][27] ), .ZN(n980) );
  OAI221_X1 U1645 ( .B1(n983), .B2(n1187), .C1(n984), .C2(n1188), .A(n1677), 
        .ZN(n1670) );
  AOI22_X1 U1646 ( .A1(n1190), .A2(\REGISTERS[15][27] ), .B1(n1191), .B2(
        \REGISTERS[14][27] ), .ZN(n1677) );
  INV_X1 U1647 ( .A(\REGISTERS[12][27] ), .ZN(n984) );
  INV_X1 U1648 ( .A(\REGISTERS[13][27] ), .ZN(n983) );
  NAND2_X1 U1649 ( .A1(n1678), .A2(n1679), .ZN(N4218) );
  NOR4_X1 U1650 ( .A1(n1680), .A2(n1681), .A3(n1682), .A4(n1683), .ZN(n1679)
         );
  OAI221_X1 U1651 ( .B1(n992), .B2(n1148), .C1(n993), .C2(n1149), .A(n1684), 
        .ZN(n1683) );
  AOI22_X1 U1652 ( .A1(n1151), .A2(\REGISTERS[19][28] ), .B1(n1152), .B2(
        \REGISTERS[18][28] ), .ZN(n1684) );
  INV_X1 U1653 ( .A(\REGISTERS[16][28] ), .ZN(n993) );
  INV_X1 U1654 ( .A(\REGISTERS[17][28] ), .ZN(n992) );
  OAI221_X1 U1655 ( .B1(n995), .B2(n1153), .C1(n996), .C2(n1154), .A(n1685), 
        .ZN(n1682) );
  AOI22_X1 U1656 ( .A1(n1156), .A2(\REGISTERS[23][28] ), .B1(n1157), .B2(
        \REGISTERS[22][28] ), .ZN(n1685) );
  INV_X1 U1657 ( .A(\REGISTERS[20][28] ), .ZN(n996) );
  INV_X1 U1658 ( .A(\REGISTERS[21][28] ), .ZN(n995) );
  OAI221_X1 U1659 ( .B1(n998), .B2(n1158), .C1(n999), .C2(n1159), .A(n1686), 
        .ZN(n1681) );
  AOI22_X1 U1660 ( .A1(n1161), .A2(\REGISTERS[27][28] ), .B1(n1162), .B2(
        \REGISTERS[26][28] ), .ZN(n1686) );
  INV_X1 U1661 ( .A(\REGISTERS[24][28] ), .ZN(n999) );
  INV_X1 U1662 ( .A(\REGISTERS[25][28] ), .ZN(n998) );
  OAI221_X1 U1663 ( .B1(n1001), .B2(n1163), .C1(n1002), .C2(n1164), .A(n1687), 
        .ZN(n1680) );
  AOI22_X1 U1664 ( .A1(n1166), .A2(\REGISTERS[29][28] ), .B1(n1167), .B2(
        \REGISTERS[28][28] ), .ZN(n1687) );
  INV_X1 U1665 ( .A(\REGISTERS[30][28] ), .ZN(n1002) );
  INV_X1 U1666 ( .A(\REGISTERS[31][28] ), .ZN(n1001) );
  NOR4_X1 U1667 ( .A1(n1688), .A2(n1689), .A3(n1690), .A4(n1691), .ZN(n1678)
         );
  AOI22_X1 U1669 ( .A1(n1175), .A2(\REGISTERS[3][28] ), .B1(n1176), .B2(
        \REGISTERS[2][28] ), .ZN(n1692) );
  INV_X1 U1670 ( .A(\REGISTERS[1][28] ), .ZN(n1008) );
  OAI221_X1 U1671 ( .B1(n1011), .B2(n1177), .C1(n1012), .C2(n1178), .A(n1693), 
        .ZN(n1690) );
  AOI22_X1 U1672 ( .A1(n1180), .A2(\REGISTERS[7][28] ), .B1(n1181), .B2(
        \REGISTERS[6][28] ), .ZN(n1693) );
  INV_X1 U1673 ( .A(\REGISTERS[4][28] ), .ZN(n1012) );
  INV_X1 U1674 ( .A(\REGISTERS[5][28] ), .ZN(n1011) );
  OAI221_X1 U1675 ( .B1(n1014), .B2(n1182), .C1(n1015), .C2(n1183), .A(n1694), 
        .ZN(n1689) );
  AOI22_X1 U1676 ( .A1(n1185), .A2(\REGISTERS[11][28] ), .B1(n1186), .B2(
        \REGISTERS[10][28] ), .ZN(n1694) );
  INV_X1 U1677 ( .A(\REGISTERS[8][28] ), .ZN(n1015) );
  INV_X1 U1678 ( .A(\REGISTERS[9][28] ), .ZN(n1014) );
  OAI221_X1 U1679 ( .B1(n1017), .B2(n1187), .C1(n1018), .C2(n1188), .A(n1695), 
        .ZN(n1688) );
  AOI22_X1 U1680 ( .A1(n1190), .A2(\REGISTERS[15][28] ), .B1(n1191), .B2(
        \REGISTERS[14][28] ), .ZN(n1695) );
  INV_X1 U1681 ( .A(\REGISTERS[12][28] ), .ZN(n1018) );
  INV_X1 U1682 ( .A(\REGISTERS[13][28] ), .ZN(n1017) );
  NAND2_X1 U1683 ( .A1(n1696), .A2(n1697), .ZN(N4217) );
  NOR4_X1 U1684 ( .A1(n1698), .A2(n1699), .A3(n1700), .A4(n1701), .ZN(n1697)
         );
  OAI221_X1 U1685 ( .B1(n1026), .B2(n1148), .C1(n1027), .C2(n1149), .A(n1702), 
        .ZN(n1701) );
  AOI22_X1 U1686 ( .A1(n1151), .A2(\REGISTERS[19][29] ), .B1(n1152), .B2(
        \REGISTERS[18][29] ), .ZN(n1702) );
  INV_X1 U1687 ( .A(\REGISTERS[16][29] ), .ZN(n1027) );
  INV_X1 U1688 ( .A(\REGISTERS[17][29] ), .ZN(n1026) );
  OAI221_X1 U1689 ( .B1(n1029), .B2(n1153), .C1(n1030), .C2(n1154), .A(n1703), 
        .ZN(n1700) );
  AOI22_X1 U1690 ( .A1(n1156), .A2(\REGISTERS[23][29] ), .B1(n1157), .B2(
        \REGISTERS[22][29] ), .ZN(n1703) );
  INV_X1 U1691 ( .A(\REGISTERS[20][29] ), .ZN(n1030) );
  INV_X1 U1692 ( .A(\REGISTERS[21][29] ), .ZN(n1029) );
  OAI221_X1 U1693 ( .B1(n1032), .B2(n1158), .C1(n1033), .C2(n1159), .A(n1704), 
        .ZN(n1699) );
  AOI22_X1 U1694 ( .A1(n1161), .A2(\REGISTERS[27][29] ), .B1(n1162), .B2(
        \REGISTERS[26][29] ), .ZN(n1704) );
  INV_X1 U1695 ( .A(\REGISTERS[24][29] ), .ZN(n1033) );
  INV_X1 U1696 ( .A(\REGISTERS[25][29] ), .ZN(n1032) );
  OAI221_X1 U1697 ( .B1(n1035), .B2(n1163), .C1(n1036), .C2(n1164), .A(n1705), 
        .ZN(n1698) );
  AOI22_X1 U1698 ( .A1(n1166), .A2(\REGISTERS[29][29] ), .B1(n1167), .B2(
        \REGISTERS[28][29] ), .ZN(n1705) );
  INV_X1 U1699 ( .A(\REGISTERS[30][29] ), .ZN(n1036) );
  INV_X1 U1700 ( .A(\REGISTERS[31][29] ), .ZN(n1035) );
  NOR4_X1 U1701 ( .A1(n1706), .A2(n1707), .A3(n1708), .A4(n1709), .ZN(n1696)
         );
  AOI22_X1 U1703 ( .A1(n1175), .A2(\REGISTERS[3][29] ), .B1(n1176), .B2(
        \REGISTERS[2][29] ), .ZN(n1710) );
  INV_X1 U1704 ( .A(\REGISTERS[1][29] ), .ZN(n1042) );
  OAI221_X1 U1705 ( .B1(n1045), .B2(n1177), .C1(n1046), .C2(n1178), .A(n1711), 
        .ZN(n1708) );
  AOI22_X1 U1706 ( .A1(n1180), .A2(\REGISTERS[7][29] ), .B1(n1181), .B2(
        \REGISTERS[6][29] ), .ZN(n1711) );
  INV_X1 U1707 ( .A(\REGISTERS[4][29] ), .ZN(n1046) );
  INV_X1 U1708 ( .A(\REGISTERS[5][29] ), .ZN(n1045) );
  OAI221_X1 U1709 ( .B1(n1048), .B2(n1182), .C1(n1049), .C2(n1183), .A(n1712), 
        .ZN(n1707) );
  AOI22_X1 U1710 ( .A1(n1185), .A2(\REGISTERS[11][29] ), .B1(n1186), .B2(
        \REGISTERS[10][29] ), .ZN(n1712) );
  INV_X1 U1711 ( .A(\REGISTERS[8][29] ), .ZN(n1049) );
  INV_X1 U1712 ( .A(\REGISTERS[9][29] ), .ZN(n1048) );
  OAI221_X1 U1713 ( .B1(n1051), .B2(n1187), .C1(n1052), .C2(n1188), .A(n1713), 
        .ZN(n1706) );
  AOI22_X1 U1714 ( .A1(n1190), .A2(\REGISTERS[15][29] ), .B1(n1191), .B2(
        \REGISTERS[14][29] ), .ZN(n1713) );
  INV_X1 U1715 ( .A(\REGISTERS[12][29] ), .ZN(n1052) );
  INV_X1 U1716 ( .A(\REGISTERS[13][29] ), .ZN(n1051) );
  NAND2_X1 U1717 ( .A1(n1714), .A2(n1715), .ZN(N4216) );
  NOR4_X1 U1718 ( .A1(n1716), .A2(n1717), .A3(n1718), .A4(n1719), .ZN(n1715)
         );
  OAI221_X1 U1719 ( .B1(n1060), .B2(n1148), .C1(n1061), .C2(n1149), .A(n1720), 
        .ZN(n1719) );
  AOI22_X1 U1720 ( .A1(n1151), .A2(\REGISTERS[19][30] ), .B1(n1152), .B2(
        \REGISTERS[18][30] ), .ZN(n1720) );
  INV_X1 U1721 ( .A(\REGISTERS[16][30] ), .ZN(n1061) );
  INV_X1 U1722 ( .A(\REGISTERS[17][30] ), .ZN(n1060) );
  OAI221_X1 U1723 ( .B1(n1063), .B2(n1153), .C1(n1064), .C2(n1154), .A(n1721), 
        .ZN(n1718) );
  AOI22_X1 U1724 ( .A1(n1156), .A2(\REGISTERS[23][30] ), .B1(n1157), .B2(
        \REGISTERS[22][30] ), .ZN(n1721) );
  INV_X1 U1725 ( .A(\REGISTERS[20][30] ), .ZN(n1064) );
  INV_X1 U1726 ( .A(\REGISTERS[21][30] ), .ZN(n1063) );
  OAI221_X1 U1727 ( .B1(n1066), .B2(n1158), .C1(n1067), .C2(n1159), .A(n1722), 
        .ZN(n1717) );
  AOI22_X1 U1728 ( .A1(n1161), .A2(\REGISTERS[27][30] ), .B1(n1162), .B2(
        \REGISTERS[26][30] ), .ZN(n1722) );
  INV_X1 U1729 ( .A(\REGISTERS[24][30] ), .ZN(n1067) );
  INV_X1 U1730 ( .A(\REGISTERS[25][30] ), .ZN(n1066) );
  OAI221_X1 U1731 ( .B1(n1069), .B2(n1163), .C1(n1070), .C2(n1164), .A(n1723), 
        .ZN(n1716) );
  AOI22_X1 U1732 ( .A1(n1166), .A2(\REGISTERS[29][30] ), .B1(n1167), .B2(
        \REGISTERS[28][30] ), .ZN(n1723) );
  INV_X1 U1733 ( .A(\REGISTERS[30][30] ), .ZN(n1070) );
  INV_X1 U1734 ( .A(\REGISTERS[31][30] ), .ZN(n1069) );
  NOR4_X1 U1735 ( .A1(n1724), .A2(n1725), .A3(n1726), .A4(n1727), .ZN(n1714)
         );
  AOI22_X1 U1737 ( .A1(n1175), .A2(\REGISTERS[3][30] ), .B1(n1176), .B2(
        \REGISTERS[2][30] ), .ZN(n1728) );
  INV_X1 U1738 ( .A(\REGISTERS[1][30] ), .ZN(n1076) );
  OAI221_X1 U1739 ( .B1(n1079), .B2(n1177), .C1(n1080), .C2(n1178), .A(n1729), 
        .ZN(n1726) );
  AOI22_X1 U1740 ( .A1(n1180), .A2(\REGISTERS[7][30] ), .B1(n1181), .B2(
        \REGISTERS[6][30] ), .ZN(n1729) );
  INV_X1 U1741 ( .A(\REGISTERS[4][30] ), .ZN(n1080) );
  INV_X1 U1742 ( .A(\REGISTERS[5][30] ), .ZN(n1079) );
  OAI221_X1 U1743 ( .B1(n1082), .B2(n1182), .C1(n1083), .C2(n1183), .A(n1730), 
        .ZN(n1725) );
  AOI22_X1 U1744 ( .A1(n1185), .A2(\REGISTERS[11][30] ), .B1(n1186), .B2(
        \REGISTERS[10][30] ), .ZN(n1730) );
  INV_X1 U1745 ( .A(\REGISTERS[8][30] ), .ZN(n1083) );
  INV_X1 U1746 ( .A(\REGISTERS[9][30] ), .ZN(n1082) );
  OAI221_X1 U1747 ( .B1(n1085), .B2(n1187), .C1(n1086), .C2(n1188), .A(n1731), 
        .ZN(n1724) );
  AOI22_X1 U1748 ( .A1(n1190), .A2(\REGISTERS[15][30] ), .B1(n1191), .B2(
        \REGISTERS[14][30] ), .ZN(n1731) );
  INV_X1 U1749 ( .A(\REGISTERS[12][30] ), .ZN(n1086) );
  INV_X1 U1750 ( .A(\REGISTERS[13][30] ), .ZN(n1085) );
  NAND2_X1 U1751 ( .A1(n1732), .A2(n1733), .ZN(N4215) );
  NOR4_X1 U1752 ( .A1(n1734), .A2(n1735), .A3(n1736), .A4(n1737), .ZN(n1733)
         );
  OAI221_X1 U1753 ( .B1(n1094), .B2(n1148), .C1(n1095), .C2(n1149), .A(n1738), 
        .ZN(n1737) );
  AOI22_X1 U1754 ( .A1(n1151), .A2(\REGISTERS[19][31] ), .B1(n1152), .B2(
        \REGISTERS[18][31] ), .ZN(n1738) );
  INV_X1 U1758 ( .A(\REGISTERS[16][31] ), .ZN(n1095) );
  INV_X1 U1760 ( .A(\REGISTERS[17][31] ), .ZN(n1094) );
  OAI221_X1 U1761 ( .B1(n1101), .B2(n1153), .C1(n1102), .C2(n1154), .A(n1743), 
        .ZN(n1736) );
  AOI22_X1 U1762 ( .A1(n1156), .A2(\REGISTERS[23][31] ), .B1(n1157), .B2(
        \REGISTERS[22][31] ), .ZN(n1743) );
  AND2_X1 U1766 ( .A1(n1746), .A2(n1747), .ZN(n1739) );
  INV_X1 U1767 ( .A(\REGISTERS[20][31] ), .ZN(n1102) );
  AND2_X1 U1769 ( .A1(n1746), .A2(ADD_RD1[0]), .ZN(n1741) );
  AND2_X1 U1770 ( .A1(ADD_RD1[4]), .A2(n1748), .ZN(n1746) );
  INV_X1 U1771 ( .A(\REGISTERS[21][31] ), .ZN(n1101) );
  OAI221_X1 U1772 ( .B1(n1109), .B2(n1158), .C1(n1110), .C2(n1159), .A(n1749), 
        .ZN(n1735) );
  AOI22_X1 U1773 ( .A1(n1161), .A2(\REGISTERS[27][31] ), .B1(n1162), .B2(
        \REGISTERS[26][31] ), .ZN(n1749) );
  INV_X1 U1777 ( .A(\REGISTERS[24][31] ), .ZN(n1110) );
  INV_X1 U1779 ( .A(\REGISTERS[25][31] ), .ZN(n1109) );
  OAI221_X1 U1780 ( .B1(n1114), .B2(n1163), .C1(n1115), .C2(n1164), .A(n1752), 
        .ZN(n1734) );
  AOI22_X1 U1781 ( .A1(n1166), .A2(\REGISTERS[29][31] ), .B1(n1167), .B2(
        \REGISTERS[28][31] ), .ZN(n1752) );
  AND2_X1 U1785 ( .A1(n1753), .A2(n1747), .ZN(n1750) );
  INV_X1 U1786 ( .A(\REGISTERS[30][31] ), .ZN(n1115) );
  AND2_X1 U1788 ( .A1(ADD_RD1[0]), .A2(n1753), .ZN(n1751) );
  AND2_X1 U1789 ( .A1(ADD_RD1[4]), .A2(ADD_RD1[3]), .ZN(n1753) );
  INV_X1 U1790 ( .A(\REGISTERS[31][31] ), .ZN(n1114) );
  NOR4_X1 U1791 ( .A1(n1754), .A2(n1755), .A3(n1756), .A4(n1757), .ZN(n1732)
         );
  AOI22_X1 U1793 ( .A1(n1175), .A2(\REGISTERS[3][31] ), .B1(n1176), .B2(
        \REGISTERS[2][31] ), .ZN(n1758) );
  INV_X1 U1798 ( .A(\REGISTERS[1][31] ), .ZN(n1122) );
  OAI221_X1 U1799 ( .B1(n1127), .B2(n1177), .C1(n1128), .C2(n1178), .A(n1761), 
        .ZN(n1756) );
  AOI22_X1 U1800 ( .A1(n1180), .A2(\REGISTERS[7][31] ), .B1(n1181), .B2(
        \REGISTERS[6][31] ), .ZN(n1761) );
  AND2_X1 U1804 ( .A1(n1762), .A2(n1747), .ZN(n1759) );
  INV_X1 U1805 ( .A(\REGISTERS[4][31] ), .ZN(n1128) );
  AND2_X1 U1807 ( .A1(n1762), .A2(ADD_RD1[0]), .ZN(n1760) );
  NOR2_X1 U1808 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[4]), .ZN(n1762) );
  INV_X1 U1809 ( .A(\REGISTERS[5][31] ), .ZN(n1127) );
  OAI221_X1 U1810 ( .B1(n1131), .B2(n1182), .C1(n1132), .C2(n1183), .A(n1763), 
        .ZN(n1755) );
  AOI22_X1 U1811 ( .A1(n1185), .A2(\REGISTERS[11][31] ), .B1(n1186), .B2(
        \REGISTERS[10][31] ), .ZN(n1763) );
  NOR2_X1 U1814 ( .A1(n1766), .A2(ADD_RD1[2]), .ZN(n1740) );
  INV_X1 U1816 ( .A(\REGISTERS[8][31] ), .ZN(n1132) );
  NOR2_X1 U1818 ( .A1(ADD_RD1[1]), .A2(ADD_RD1[2]), .ZN(n1742) );
  INV_X1 U1819 ( .A(\REGISTERS[9][31] ), .ZN(n1131) );
  OAI221_X1 U1820 ( .B1(n1137), .B2(n1187), .C1(n1138), .C2(n1188), .A(n1767), 
        .ZN(n1754) );
  AOI22_X1 U1821 ( .A1(n1190), .A2(\REGISTERS[15][31] ), .B1(n1191), .B2(
        \REGISTERS[14][31] ), .ZN(n1767) );
  NOR2_X1 U1824 ( .A1(n1768), .A2(n1766), .ZN(n1744) );
  INV_X1 U1825 ( .A(ADD_RD1[1]), .ZN(n1766) );
  AND2_X1 U1827 ( .A1(n1769), .A2(n1747), .ZN(n1764) );
  INV_X1 U1828 ( .A(ADD_RD1[0]), .ZN(n1747) );
  INV_X1 U1829 ( .A(\REGISTERS[12][31] ), .ZN(n1138) );
  INV_X1 U1832 ( .A(ADD_RD1[2]), .ZN(n1768) );
  AND2_X1 U1833 ( .A1(n1769), .A2(ADD_RD1[0]), .ZN(n1765) );
  NOR2_X1 U1834 ( .A1(n1748), .A2(ADD_RD1[4]), .ZN(n1769) );
  INV_X1 U1835 ( .A(ADD_RD1[3]), .ZN(n1748) );
  INV_X1 U1836 ( .A(\REGISTERS[13][31] ), .ZN(n1137) );
  NAND2_X1 U1837 ( .A1(n1770), .A2(n193), .ZN(N4083) );
  NAND3_X1 U1838 ( .A1(n1771), .A2(n1), .A3(n1773), .ZN(n1770) );
  NAND2_X1 U1839 ( .A1(n1774), .A2(n193), .ZN(N4019) );
  NAND3_X1 U1840 ( .A1(n1773), .A2(n1772), .A3(n1775), .ZN(n1774) );
  NAND2_X1 U1841 ( .A1(n1776), .A2(n193), .ZN(N3955) );
  NAND3_X1 U1842 ( .A1(n1773), .A2(n1772), .A3(n1777), .ZN(n1776) );
  NAND2_X1 U1843 ( .A1(n1778), .A2(n193), .ZN(N3891) );
  NAND3_X1 U1844 ( .A1(n1773), .A2(n1772), .A3(n1779), .ZN(n1778) );
  NAND2_X1 U1845 ( .A1(n1780), .A2(n193), .ZN(N3827) );
  NAND3_X1 U1846 ( .A1(n1773), .A2(n1772), .A3(n1781), .ZN(n1780) );
  NAND2_X1 U1847 ( .A1(n1782), .A2(n193), .ZN(N3763) );
  NAND3_X1 U1848 ( .A1(n1773), .A2(n1772), .A3(n1783), .ZN(n1782) );
  NAND2_X1 U1849 ( .A1(n1784), .A2(n193), .ZN(N3699) );
  NAND3_X1 U1850 ( .A1(n1773), .A2(n1772), .A3(n1785), .ZN(n1784) );
  NOR2_X1 U1851 ( .A1(ADD_WR[3]), .A2(ADD_WR[4]), .ZN(n1773) );
  NAND2_X1 U1852 ( .A1(n1786), .A2(n193), .ZN(N3635) );
  NAND3_X1 U1853 ( .A1(n1787), .A2(n1772), .A3(n1788), .ZN(n1786) );
  NAND2_X1 U1854 ( .A1(n1789), .A2(n193), .ZN(N3571) );
  NAND3_X1 U1855 ( .A1(n1771), .A2(n1772), .A3(n1787), .ZN(n1789) );
  NAND2_X1 U1856 ( .A1(n1790), .A2(n193), .ZN(N3507) );
  NAND3_X1 U1857 ( .A1(n1775), .A2(n1772), .A3(n1787), .ZN(n1790) );
  NAND2_X1 U1858 ( .A1(n1791), .A2(n193), .ZN(N3443) );
  NAND3_X1 U1859 ( .A1(n1777), .A2(n1772), .A3(n1787), .ZN(n1791) );
  NAND2_X1 U1860 ( .A1(n1792), .A2(n193), .ZN(N3379) );
  NAND3_X1 U1861 ( .A1(n1779), .A2(n1772), .A3(n1787), .ZN(n1792) );
  NAND2_X1 U1862 ( .A1(n1793), .A2(n227), .ZN(N3315) );
  NAND3_X1 U1863 ( .A1(n1781), .A2(n1772), .A3(n1787), .ZN(n1793) );
  NAND2_X1 U1864 ( .A1(n1794), .A2(n227), .ZN(N3251) );
  NAND3_X1 U1865 ( .A1(n1783), .A2(n1772), .A3(n1787), .ZN(n1794) );
  NAND2_X1 U1866 ( .A1(n1795), .A2(n227), .ZN(N3187) );
  NAND3_X1 U1867 ( .A1(n1785), .A2(n1772), .A3(n1787), .ZN(n1795) );
  NOR2_X1 U1868 ( .A1(n1796), .A2(ADD_WR[4]), .ZN(n1787) );
  NAND2_X1 U1869 ( .A1(n1797), .A2(n227), .ZN(N3123) );
  NAND3_X1 U1870 ( .A1(n1788), .A2(n1772), .A3(n1798), .ZN(n1797) );
  NAND2_X1 U1871 ( .A1(n1799), .A2(n227), .ZN(N3059) );
  NAND3_X1 U1872 ( .A1(n1771), .A2(n1772), .A3(n1798), .ZN(n1799) );
  NAND2_X1 U1873 ( .A1(n1800), .A2(n227), .ZN(N2995) );
  NAND3_X1 U1874 ( .A1(n1775), .A2(n1772), .A3(n1798), .ZN(n1800) );
  NAND2_X1 U1875 ( .A1(n1801), .A2(n227), .ZN(N2931) );
  NAND3_X1 U1876 ( .A1(n1777), .A2(n1772), .A3(n1798), .ZN(n1801) );
  NAND2_X1 U1877 ( .A1(n1802), .A2(n227), .ZN(N2867) );
  NAND3_X1 U1878 ( .A1(n1779), .A2(n1772), .A3(n1798), .ZN(n1802) );
  NAND2_X1 U1879 ( .A1(n1803), .A2(n227), .ZN(N2803) );
  NAND3_X1 U1880 ( .A1(n1781), .A2(n1772), .A3(n1798), .ZN(n1803) );
  NAND2_X1 U1881 ( .A1(n1804), .A2(n227), .ZN(N2739) );
  NAND3_X1 U1882 ( .A1(n1783), .A2(n1772), .A3(n1798), .ZN(n1804) );
  NAND2_X1 U1883 ( .A1(n1805), .A2(n227), .ZN(N2675) );
  NAND3_X1 U1884 ( .A1(n1785), .A2(n1772), .A3(n1798), .ZN(n1805) );
  AND2_X1 U1885 ( .A1(ADD_WR[4]), .A2(n1796), .ZN(n1798) );
  INV_X1 U1886 ( .A(ADD_WR[3]), .ZN(n1796) );
  NAND2_X1 U1887 ( .A1(n1806), .A2(n227), .ZN(N2611) );
  NAND3_X1 U1888 ( .A1(n1788), .A2(n1772), .A3(n1807), .ZN(n1806) );
  NOR3_X1 U1889 ( .A1(ADD_WR[1]), .A2(ADD_WR[2]), .A3(ADD_WR[0]), .ZN(n1788)
         );
  NAND2_X1 U1890 ( .A1(n1808), .A2(n261), .ZN(N2547) );
  NAND3_X1 U1891 ( .A1(n1771), .A2(n1772), .A3(n1807), .ZN(n1808) );
  NOR3_X1 U1892 ( .A1(ADD_WR[1]), .A2(ADD_WR[2]), .A3(n1809), .ZN(n1771) );
  NAND2_X1 U1893 ( .A1(n1810), .A2(n261), .ZN(N2483) );
  NAND3_X1 U1894 ( .A1(n1775), .A2(n1772), .A3(n1807), .ZN(n1810) );
  NOR3_X1 U1895 ( .A1(ADD_WR[0]), .A2(ADD_WR[2]), .A3(n1811), .ZN(n1775) );
  NAND2_X1 U1896 ( .A1(n1812), .A2(n261), .ZN(N2419) );
  NAND3_X1 U1897 ( .A1(n1777), .A2(n1), .A3(n1807), .ZN(n1812) );
  NOR3_X1 U1898 ( .A1(n1809), .A2(ADD_WR[2]), .A3(n1811), .ZN(n1777) );
  NAND2_X1 U1899 ( .A1(n1813), .A2(n261), .ZN(N2355) );
  NAND3_X1 U1900 ( .A1(n1779), .A2(n1), .A3(n1807), .ZN(n1813) );
  NOR3_X1 U1901 ( .A1(ADD_WR[0]), .A2(ADD_WR[1]), .A3(n1814), .ZN(n1779) );
  NAND2_X1 U1902 ( .A1(n1815), .A2(n261), .ZN(N2291) );
  NAND3_X1 U1903 ( .A1(n1781), .A2(n1), .A3(n1807), .ZN(n1815) );
  NOR3_X1 U1904 ( .A1(n1809), .A2(ADD_WR[1]), .A3(n1814), .ZN(n1781) );
  NAND2_X1 U1905 ( .A1(n1816), .A2(n261), .ZN(N2227) );
  NAND3_X1 U1906 ( .A1(n1783), .A2(n1), .A3(n1807), .ZN(n1816) );
  NOR3_X1 U1907 ( .A1(n1811), .A2(ADD_WR[0]), .A3(n1814), .ZN(n1783) );
  AND2_X1 U1908 ( .A1(DATAIN[31]), .A2(n261), .ZN(N4148) );
  AND2_X1 U1909 ( .A1(DATAIN[30]), .A2(n329), .ZN(N4146) );
  AND2_X1 U1910 ( .A1(DATAIN[29]), .A2(n329), .ZN(N4144) );
  AND2_X1 U1911 ( .A1(DATAIN[28]), .A2(n329), .ZN(N4142) );
  AND2_X1 U1912 ( .A1(DATAIN[27]), .A2(n329), .ZN(N4140) );
  AND2_X1 U1913 ( .A1(DATAIN[26]), .A2(n329), .ZN(N4138) );
  AND2_X1 U1914 ( .A1(DATAIN[25]), .A2(n329), .ZN(N4136) );
  AND2_X1 U1915 ( .A1(DATAIN[24]), .A2(n329), .ZN(N4134) );
  AND2_X1 U1916 ( .A1(DATAIN[23]), .A2(n329), .ZN(N4132) );
  AND2_X1 U1917 ( .A1(DATAIN[22]), .A2(n329), .ZN(N4130) );
  AND2_X1 U1918 ( .A1(DATAIN[21]), .A2(n329), .ZN(N4128) );
  AND2_X1 U1919 ( .A1(DATAIN[20]), .A2(n295), .ZN(N4126) );
  AND2_X1 U1920 ( .A1(DATAIN[19]), .A2(n295), .ZN(N4124) );
  AND2_X1 U1921 ( .A1(DATAIN[18]), .A2(n295), .ZN(N4122) );
  AND2_X1 U1922 ( .A1(DATAIN[17]), .A2(n295), .ZN(N4120) );
  AND2_X1 U1923 ( .A1(DATAIN[16]), .A2(n295), .ZN(N4118) );
  AND2_X1 U1924 ( .A1(DATAIN[15]), .A2(n295), .ZN(N4116) );
  AND2_X1 U1925 ( .A1(DATAIN[14]), .A2(n295), .ZN(N4114) );
  AND2_X1 U1926 ( .A1(DATAIN[13]), .A2(n295), .ZN(N4112) );
  AND2_X1 U1927 ( .A1(DATAIN[12]), .A2(n295), .ZN(N4110) );
  AND2_X1 U1928 ( .A1(DATAIN[11]), .A2(n295), .ZN(N4108) );
  AND2_X1 U1929 ( .A1(DATAIN[10]), .A2(n295), .ZN(N4106) );
  AND2_X1 U1930 ( .A1(DATAIN[9]), .A2(n295), .ZN(N4104) );
  AND2_X1 U1931 ( .A1(DATAIN[8]), .A2(n295), .ZN(N4102) );
  AND2_X1 U1932 ( .A1(DATAIN[7]), .A2(n295), .ZN(N4100) );
  AND2_X1 U1933 ( .A1(DATAIN[6]), .A2(n295), .ZN(N4098) );
  AND2_X1 U1934 ( .A1(DATAIN[5]), .A2(n295), .ZN(N4096) );
  AND2_X1 U1935 ( .A1(DATAIN[4]), .A2(n261), .ZN(N4094) );
  AND2_X1 U1936 ( .A1(DATAIN[3]), .A2(n261), .ZN(N4092) );
  AND2_X1 U1937 ( .A1(DATAIN[2]), .A2(n261), .ZN(N4090) );
  AND2_X1 U1938 ( .A1(DATAIN[1]), .A2(n261), .ZN(N4088) );
  AND2_X1 U1939 ( .A1(DATAIN[0]), .A2(n261), .ZN(N4086) );
  NAND2_X1 U1940 ( .A1(n1817), .A2(n261), .ZN(N2163) );
  NAND3_X1 U1941 ( .A1(n1785), .A2(n1), .A3(n1807), .ZN(n1817) );
  AND2_X1 U1942 ( .A1(ADD_WR[4]), .A2(ADD_WR[3]), .ZN(n1807) );
  AND2_X1 U1943 ( .A1(WR), .A2(ENABLE), .ZN(n1772) );
  NOR3_X1 U1944 ( .A1(n1811), .A2(n1809), .A3(n1814), .ZN(n1785) );
  INV_X1 U1945 ( .A(ADD_WR[2]), .ZN(n1814) );
  INV_X1 U1946 ( .A(ADD_WR[0]), .ZN(n1809) );
  INV_X1 U1947 ( .A(ADD_WR[1]), .ZN(n1811) );
  NOR2_X2 U3 ( .A1(n1140), .A2(ADD_RD2[1]), .ZN(n1105) );
  NOR2_X2 U4 ( .A1(n1768), .A2(ADD_RD1[1]), .ZN(n1745) );
  CLKBUF_X1 U5 ( .A(n1772), .Z(n1) );
  AND2_X2 U6 ( .A1(n1759), .A2(n1744), .ZN(n1181) );
  AND2_X2 U7 ( .A1(n1764), .A2(n1744), .ZN(n1191) );
  AND2_X2 U8 ( .A1(n1739), .A2(n1740), .ZN(n1152) );
  AND2_X2 U9 ( .A1(n1745), .A2(n1750), .ZN(n1167) );
  AND2_X2 U10 ( .A1(n1740), .A2(n1750), .ZN(n1162) );
  AND2_X2 U11 ( .A1(n1759), .A2(n1740), .ZN(n1176) );
  AND2_X2 U12 ( .A1(n1764), .A2(n1740), .ZN(n1186) );
  NAND2_X2 U13 ( .A1(n1125), .A2(n1105), .ZN(n49) );
  AND2_X2 U14 ( .A1(n1739), .A2(n1744), .ZN(n1157) );
  NAND2_X2 U15 ( .A1(n1097), .A2(n1105), .ZN(n17) );
  NAND2_X2 U16 ( .A1(n1100), .A2(n1112), .ZN(n24) );
  NAND2_X2 U17 ( .A1(n1134), .A2(n1105), .ZN(n63) );
  NAND2_X2 U18 ( .A1(n1112), .A2(n1104), .ZN(n31) );
  NAND2_X2 U19 ( .A1(n1134), .A2(n1100), .ZN(n56) );
  NAND2_X2 U20 ( .A1(n1097), .A2(n1100), .ZN(n10) );
  NAND2_X2 U21 ( .A1(n1760), .A2(n1742), .ZN(n1172) );
  NAND2_X2 U22 ( .A1(n1759), .A2(n1745), .ZN(n1178) );
  NAND2_X2 U23 ( .A1(n1750), .A2(n1744), .ZN(n1164) );
  NAND2_X2 U24 ( .A1(n1742), .A2(n1750), .ZN(n1159) );
  NAND2_X2 U25 ( .A1(n1764), .A2(n1742), .ZN(n1183) );
  NAND2_X2 U26 ( .A1(n1739), .A2(n1742), .ZN(n1149) );
  NAND2_X2 U27 ( .A1(n1764), .A2(n1745), .ZN(n1188) );
  NAND2_X2 U28 ( .A1(n1739), .A2(n1745), .ZN(n1154) );
  AND2_X2 U29 ( .A1(n1097), .A2(n1098), .ZN(n14) );
  AND2_X2 U30 ( .A1(n1125), .A2(n1098), .ZN(n46) );
  AND2_X2 U31 ( .A1(n1097), .A2(n1104), .ZN(n21) );
  AND2_X2 U32 ( .A1(n1134), .A2(n1104), .ZN(n67) );
  AND2_X2 U33 ( .A1(n1105), .A2(n1112), .ZN(n35) );
  AND2_X2 U34 ( .A1(n1134), .A2(n1098), .ZN(n60) );
  AND2_X2 U47 ( .A1(n1098), .A2(n1112), .ZN(n28) );
  NAND2_X2 U66 ( .A1(n1765), .A2(n1745), .ZN(n1187) );
  AND2_X2 U85 ( .A1(n1125), .A2(n1104), .ZN(n53) );
  NAND2_X2 U104 ( .A1(n1741), .A2(n1742), .ZN(n1148) );
  NAND2_X2 U123 ( .A1(n1744), .A2(n1751), .ZN(n1163) );
  NAND2_X2 U142 ( .A1(n1765), .A2(n1742), .ZN(n1182) );
  NAND2_X2 U161 ( .A1(n1760), .A2(n1745), .ZN(n1177) );
  NAND2_X2 U180 ( .A1(n1741), .A2(n1745), .ZN(n1153) );
  NAND2_X2 U199 ( .A1(n1742), .A2(n1751), .ZN(n1158) );
  AND2_X2 U218 ( .A1(n1740), .A2(n1751), .ZN(n1161) );
  AND2_X2 U237 ( .A1(n1745), .A2(n1751), .ZN(n1166) );
  AND2_X2 U256 ( .A1(n1760), .A2(n1740), .ZN(n1175) );
  AND2_X2 U275 ( .A1(n1741), .A2(n1744), .ZN(n1156) );
  AND2_X2 U294 ( .A1(n1741), .A2(n1740), .ZN(n1151) );
  AND2_X2 U313 ( .A1(n1760), .A2(n1744), .ZN(n1180) );
  AND2_X2 U332 ( .A1(n1765), .A2(n1740), .ZN(n1185) );
  AND2_X2 U351 ( .A1(n1765), .A2(n1744), .ZN(n1190) );
  AND2_X2 U370 ( .A1(n1126), .A2(n1104), .ZN(n52) );
  AND2_X2 U389 ( .A1(n1099), .A2(n1098), .ZN(n13) );
  AND2_X2 U408 ( .A1(n1099), .A2(n1104), .ZN(n20) );
  AND2_X2 U427 ( .A1(n1126), .A2(n1098), .ZN(n45) );
  AND2_X2 U446 ( .A1(n1135), .A2(n1098), .ZN(n59) );
  AND2_X2 U465 ( .A1(n1135), .A2(n1104), .ZN(n66) );
  AND2_X2 U484 ( .A1(n1098), .A2(n1113), .ZN(n27) );
  AND2_X2 U503 ( .A1(n1105), .A2(n1113), .ZN(n34) );
  NAND2_X2 U522 ( .A1(n1104), .A2(n1113), .ZN(n29) );
  NAND2_X2 U541 ( .A1(n1126), .A2(n1105), .ZN(n47) );
  NAND2_X2 U560 ( .A1(n1135), .A2(n1100), .ZN(n54) );
  NAND2_X2 U579 ( .A1(n1100), .A2(n1113), .ZN(n22) );
  NAND2_X2 U598 ( .A1(n1099), .A2(n1105), .ZN(n15) );
  NAND2_X2 U617 ( .A1(n1135), .A2(n1105), .ZN(n61) );
  NAND2_X2 U629 ( .A1(n1126), .A2(n1100), .ZN(n40) );
  NAND2_X2 U630 ( .A1(n1099), .A2(n1100), .ZN(n8) );
  OAI21_X1 U639 ( .B1(n40), .B2(n41), .A(n44), .ZN(n39) );
  OAI21_X1 U644 ( .B1(n40), .B2(n90), .A(n92), .ZN(n89) );
  OAI21_X1 U645 ( .B1(n40), .B2(n124), .A(n126), .ZN(n123) );
  OAI21_X1 U646 ( .B1(n40), .B2(n158), .A(n160), .ZN(n157) );
  OAI21_X1 U647 ( .B1(n40), .B2(n192), .A(n194), .ZN(n191) );
  OAI21_X1 U650 ( .B1(n40), .B2(n226), .A(n228), .ZN(n225) );
  OAI21_X1 U651 ( .B1(n40), .B2(n260), .A(n262), .ZN(n259) );
  OAI21_X1 U652 ( .B1(n40), .B2(n294), .A(n296), .ZN(n293) );
  OAI21_X1 U654 ( .B1(n40), .B2(n328), .A(n330), .ZN(n327) );
  OAI21_X1 U658 ( .B1(n40), .B2(n362), .A(n364), .ZN(n361) );
  OAI21_X1 U660 ( .B1(n40), .B2(n396), .A(n398), .ZN(n395) );
  OAI21_X1 U661 ( .B1(n40), .B2(n430), .A(n432), .ZN(n429) );
  OAI21_X1 U662 ( .B1(n40), .B2(n464), .A(n466), .ZN(n463) );
  OAI21_X1 U663 ( .B1(n40), .B2(n498), .A(n500), .ZN(n497) );
  OAI21_X1 U666 ( .B1(n40), .B2(n532), .A(n534), .ZN(n531) );
  OAI21_X1 U667 ( .B1(n40), .B2(n566), .A(n568), .ZN(n565) );
  OAI21_X1 U668 ( .B1(n40), .B2(n600), .A(n602), .ZN(n599) );
  OAI21_X1 U670 ( .B1(n40), .B2(n634), .A(n636), .ZN(n633) );
  OAI21_X1 U675 ( .B1(n40), .B2(n668), .A(n670), .ZN(n667) );
  OAI21_X1 U676 ( .B1(n40), .B2(n702), .A(n704), .ZN(n701) );
  OAI21_X1 U678 ( .B1(n40), .B2(n736), .A(n738), .ZN(n735) );
  OAI21_X1 U679 ( .B1(n40), .B2(n770), .A(n772), .ZN(n769) );
  OAI21_X1 U683 ( .B1(n40), .B2(n804), .A(n806), .ZN(n803) );
  OAI21_X1 U684 ( .B1(n40), .B2(n838), .A(n840), .ZN(n837) );
  OAI21_X1 U687 ( .B1(n40), .B2(n872), .A(n874), .ZN(n871) );
  OAI21_X1 U690 ( .B1(n40), .B2(n906), .A(n908), .ZN(n905) );
  OAI21_X1 U691 ( .B1(n40), .B2(n940), .A(n942), .ZN(n939) );
  OAI21_X1 U716 ( .B1(n40), .B2(n974), .A(n976), .ZN(n973) );
  OAI21_X1 U750 ( .B1(n40), .B2(n1008), .A(n1010), .ZN(n1007) );
  OAI21_X1 U784 ( .B1(n40), .B2(n1042), .A(n1044), .ZN(n1041) );
  OAI21_X1 U818 ( .B1(n40), .B2(n1076), .A(n1078), .ZN(n1075) );
  OAI21_X1 U852 ( .B1(n40), .B2(n1122), .A(n1124), .ZN(n1121) );
  OAI21_X1 U886 ( .B1(n41), .B2(n1172), .A(n1174), .ZN(n1171) );
  OAI21_X1 U920 ( .B1(n90), .B2(n1172), .A(n1206), .ZN(n1205) );
  OAI21_X1 U954 ( .B1(n124), .B2(n1172), .A(n1224), .ZN(n1223) );
  OAI21_X1 U988 ( .B1(n158), .B2(n1172), .A(n1242), .ZN(n1241) );
  OAI21_X1 U1022 ( .B1(n192), .B2(n1172), .A(n1260), .ZN(n1259) );
  OAI21_X1 U1056 ( .B1(n226), .B2(n1172), .A(n1278), .ZN(n1277) );
  OAI21_X1 U1090 ( .B1(n260), .B2(n1172), .A(n1296), .ZN(n1295) );
  OAI21_X1 U1124 ( .B1(n294), .B2(n1172), .A(n1314), .ZN(n1313) );
  OAI21_X1 U1158 ( .B1(n328), .B2(n1172), .A(n1332), .ZN(n1331) );
  OAI21_X1 U1192 ( .B1(n362), .B2(n1172), .A(n1350), .ZN(n1349) );
  OAI21_X1 U1226 ( .B1(n396), .B2(n1172), .A(n1368), .ZN(n1367) );
  OAI21_X1 U1260 ( .B1(n430), .B2(n1172), .A(n1386), .ZN(n1385) );
  OAI21_X1 U1294 ( .B1(n464), .B2(n1172), .A(n1404), .ZN(n1403) );
  OAI21_X1 U1328 ( .B1(n498), .B2(n1172), .A(n1422), .ZN(n1421) );
  OAI21_X1 U1362 ( .B1(n532), .B2(n1172), .A(n1440), .ZN(n1439) );
  OAI21_X1 U1396 ( .B1(n566), .B2(n1172), .A(n1458), .ZN(n1457) );
  OAI21_X1 U1430 ( .B1(n600), .B2(n1172), .A(n1476), .ZN(n1475) );
  OAI21_X1 U1464 ( .B1(n634), .B2(n1172), .A(n1494), .ZN(n1493) );
  OAI21_X1 U1498 ( .B1(n668), .B2(n1172), .A(n1512), .ZN(n1511) );
  OAI21_X1 U1532 ( .B1(n702), .B2(n1172), .A(n1530), .ZN(n1529) );
  OAI21_X1 U1566 ( .B1(n736), .B2(n1172), .A(n1548), .ZN(n1547) );
  OAI21_X1 U1600 ( .B1(n770), .B2(n1172), .A(n1566), .ZN(n1565) );
  OAI21_X1 U1634 ( .B1(n804), .B2(n1172), .A(n1584), .ZN(n1583) );
  OAI21_X1 U1668 ( .B1(n838), .B2(n1172), .A(n1602), .ZN(n1601) );
  OAI21_X1 U1702 ( .B1(n872), .B2(n1172), .A(n1620), .ZN(n1619) );
  OAI21_X1 U1736 ( .B1(n906), .B2(n1172), .A(n1638), .ZN(n1637) );
  OAI21_X1 U1755 ( .B1(n940), .B2(n1172), .A(n1656), .ZN(n1655) );
  OAI21_X1 U1756 ( .B1(n974), .B2(n1172), .A(n1674), .ZN(n1673) );
  OAI21_X1 U1757 ( .B1(n1008), .B2(n1172), .A(n1692), .ZN(n1691) );
  OAI21_X1 U1759 ( .B1(n1042), .B2(n1172), .A(n1710), .ZN(n1709) );
  OAI21_X1 U1763 ( .B1(n1076), .B2(n1172), .A(n1728), .ZN(n1727) );
  OAI21_X1 U1764 ( .B1(n1122), .B2(n1172), .A(n1758), .ZN(n1757) );
  CLKBUF_X1 U631 ( .A(RESET), .Z(n193) );
  CLKBUF_X1 U632 ( .A(RESET), .Z(n227) );
  CLKBUF_X1 U635 ( .A(RESET), .Z(n261) );
  CLKBUF_X1 U636 ( .A(RESET), .Z(n295) );
  CLKBUF_X1 U637 ( .A(RESET), .Z(n329) );
endmodule


module alu_NUMBIT32 ( DATA1, DATA2, .FUNC({\FUNC[4] , \FUNC[3] , \FUNC[2] , 
        \FUNC[1] , \FUNC[0] }), OUTALU );
  input [31:0] DATA1;
  input [31:0] DATA2;
  output [31:0] OUTALU;
  input \FUNC[4] , \FUNC[3] , \FUNC[2] , \FUNC[1] , \FUNC[0] ;
  wire   sub_add, \Sel[2] , sign_unsign, \CU_OUT[0] , Adder_Cout, n104, n205,
         n305, n306, n308, n310, n311, n312, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n352, n353, n355,
         n356, n360, n359, n358, n357, n354, n349, n313, n309, n307, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379;
  wire   [1:0] Conf;
  wire   [2:0] Comp_OP;
  wire   [31:0] OUT_adder;
  wire   [31:0] LU_out;
  wire   [31:0] SHIFT_OUT;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30;

  CLKBUF_X2 U233 ( .A(n104), .Z(n306) );
  INV_X1 U241 ( .A(n315), .ZN(OUTALU[9]) );
  AOI222_X1 U242 ( .A1(OUT_adder[9]), .A2(n316), .B1(LU_out[9]), .B2(n317), 
        .C1(SHIFT_OUT[9]), .C2(n318), .ZN(n315) );
  INV_X1 U243 ( .A(n319), .ZN(OUTALU[8]) );
  AOI222_X1 U244 ( .A1(OUT_adder[8]), .A2(n316), .B1(LU_out[8]), .B2(n317), 
        .C1(SHIFT_OUT[8]), .C2(n318), .ZN(n319) );
  INV_X1 U245 ( .A(n320), .ZN(OUTALU[7]) );
  AOI222_X1 U246 ( .A1(OUT_adder[7]), .A2(n316), .B1(LU_out[7]), .B2(n317), 
        .C1(SHIFT_OUT[7]), .C2(n318), .ZN(n320) );
  INV_X1 U247 ( .A(n321), .ZN(OUTALU[6]) );
  AOI222_X1 U248 ( .A1(OUT_adder[6]), .A2(n316), .B1(LU_out[6]), .B2(n317), 
        .C1(SHIFT_OUT[6]), .C2(n318), .ZN(n321) );
  INV_X1 U249 ( .A(n322), .ZN(OUTALU[5]) );
  AOI222_X1 U250 ( .A1(OUT_adder[5]), .A2(n316), .B1(LU_out[5]), .B2(n317), 
        .C1(SHIFT_OUT[5]), .C2(n318), .ZN(n322) );
  INV_X1 U251 ( .A(n323), .ZN(OUTALU[4]) );
  AOI222_X1 U252 ( .A1(OUT_adder[4]), .A2(n316), .B1(LU_out[4]), .B2(n317), 
        .C1(SHIFT_OUT[4]), .C2(n318), .ZN(n323) );
  INV_X1 U253 ( .A(n324), .ZN(OUTALU[3]) );
  AOI222_X1 U254 ( .A1(n368), .A2(n316), .B1(LU_out[3]), .B2(n317), .C1(
        SHIFT_OUT[3]), .C2(n318), .ZN(n324) );
  INV_X1 U255 ( .A(n325), .ZN(OUTALU[31]) );
  AOI222_X1 U256 ( .A1(OUT_adder[31]), .A2(n316), .B1(LU_out[31]), .B2(n317), 
        .C1(SHIFT_OUT[31]), .C2(n318), .ZN(n325) );
  INV_X1 U257 ( .A(n326), .ZN(OUTALU[30]) );
  INV_X1 U259 ( .A(n327), .ZN(OUTALU[2]) );
  AOI222_X1 U260 ( .A1(OUT_adder[2]), .A2(n316), .B1(LU_out[2]), .B2(n317), 
        .C1(SHIFT_OUT[2]), .C2(n318), .ZN(n327) );
  INV_X1 U261 ( .A(n328), .ZN(OUTALU[29]) );
  INV_X1 U263 ( .A(n329), .ZN(OUTALU[28]) );
  INV_X1 U265 ( .A(n330), .ZN(OUTALU[27]) );
  AOI222_X1 U266 ( .A1(n378), .A2(n316), .B1(LU_out[27]), .B2(n317), .C1(
        SHIFT_OUT[27]), .C2(n318), .ZN(n330) );
  INV_X1 U267 ( .A(n331), .ZN(OUTALU[26]) );
  INV_X1 U269 ( .A(n332), .ZN(OUTALU[25]) );
  AOI222_X1 U270 ( .A1(OUT_adder[25]), .A2(n316), .B1(LU_out[25]), .B2(n317), 
        .C1(SHIFT_OUT[25]), .C2(n318), .ZN(n332) );
  INV_X1 U271 ( .A(n333), .ZN(OUTALU[24]) );
  INV_X1 U273 ( .A(n334), .ZN(OUTALU[23]) );
  AOI222_X1 U274 ( .A1(OUT_adder[23]), .A2(n316), .B1(LU_out[23]), .B2(n317), 
        .C1(SHIFT_OUT[23]), .C2(n318), .ZN(n334) );
  INV_X1 U275 ( .A(n335), .ZN(OUTALU[22]) );
  AOI222_X1 U276 ( .A1(OUT_adder[22]), .A2(n316), .B1(LU_out[22]), .B2(n317), 
        .C1(SHIFT_OUT[22]), .C2(n318), .ZN(n335) );
  INV_X1 U277 ( .A(n336), .ZN(OUTALU[21]) );
  INV_X1 U279 ( .A(n337), .ZN(OUTALU[20]) );
  INV_X1 U281 ( .A(n338), .ZN(OUTALU[1]) );
  AOI222_X1 U282 ( .A1(OUT_adder[1]), .A2(n316), .B1(LU_out[1]), .B2(n317), 
        .C1(SHIFT_OUT[1]), .C2(n318), .ZN(n338) );
  INV_X1 U283 ( .A(n339), .ZN(OUTALU[19]) );
  AOI222_X1 U284 ( .A1(OUT_adder[19]), .A2(n316), .B1(LU_out[19]), .B2(n317), 
        .C1(SHIFT_OUT[19]), .C2(n318), .ZN(n339) );
  INV_X1 U285 ( .A(n340), .ZN(OUTALU[18]) );
  AOI222_X1 U286 ( .A1(OUT_adder[18]), .A2(n316), .B1(LU_out[18]), .B2(n317), 
        .C1(SHIFT_OUT[18]), .C2(n318), .ZN(n340) );
  INV_X1 U287 ( .A(n341), .ZN(OUTALU[17]) );
  AOI222_X1 U288 ( .A1(OUT_adder[17]), .A2(n316), .B1(LU_out[17]), .B2(n317), 
        .C1(SHIFT_OUT[17]), .C2(n318), .ZN(n341) );
  INV_X1 U289 ( .A(n342), .ZN(OUTALU[16]) );
  INV_X1 U291 ( .A(n343), .ZN(OUTALU[15]) );
  AOI222_X1 U292 ( .A1(OUT_adder[15]), .A2(n316), .B1(LU_out[15]), .B2(n317), 
        .C1(SHIFT_OUT[15]), .C2(n318), .ZN(n343) );
  INV_X1 U293 ( .A(n344), .ZN(OUTALU[14]) );
  AOI222_X1 U294 ( .A1(OUT_adder[14]), .A2(n316), .B1(LU_out[14]), .B2(n317), 
        .C1(SHIFT_OUT[14]), .C2(n318), .ZN(n344) );
  INV_X1 U295 ( .A(n345), .ZN(OUTALU[13]) );
  AOI222_X1 U296 ( .A1(OUT_adder[13]), .A2(n316), .B1(LU_out[13]), .B2(n317), 
        .C1(SHIFT_OUT[13]), .C2(n318), .ZN(n345) );
  INV_X1 U297 ( .A(n346), .ZN(OUTALU[12]) );
  AOI222_X1 U298 ( .A1(OUT_adder[12]), .A2(n316), .B1(LU_out[12]), .B2(n317), 
        .C1(SHIFT_OUT[12]), .C2(n318), .ZN(n346) );
  INV_X1 U299 ( .A(n347), .ZN(OUTALU[11]) );
  AOI222_X1 U300 ( .A1(OUT_adder[11]), .A2(n316), .B1(LU_out[11]), .B2(n317), 
        .C1(SHIFT_OUT[11]), .C2(n318), .ZN(n347) );
  INV_X1 U301 ( .A(n348), .ZN(OUTALU[10]) );
  AOI222_X1 U302 ( .A1(OUT_adder[10]), .A2(n316), .B1(LU_out[10]), .B2(n317), 
        .C1(SHIFT_OUT[10]), .C2(n318), .ZN(n348) );
  NAND3_X1 U305 ( .A1(n352), .A2(n308), .A3(n353), .ZN(n314) );
  OAI21_X1 U309 ( .B1(n311), .B2(n312), .A(n356), .ZN(n205) );
  INV_X1 U310 ( .A(n352), .ZN(n311) );
  NOR2_X1 U318 ( .A1(FUNC[4]), .A2(FUNC[3]), .ZN(n353) );
  AOI21_X1 U321 ( .B1(n312), .B2(n356), .A(n308), .ZN(Comp_OP[0]) );
  NOR2_X1 U327 ( .A1(n360), .A2(FUNC[4]), .ZN(n355) );
  INV_X1 U328 ( .A(FUNC[3]), .ZN(n360) );
  P4addersub_N32 P4addersub_0 ( .A({DATA1[31:29], n367, DATA1[27:0]}), .B(
        DATA2), .sub_add(n305), .Y(OUT_adder), .Cout(Adder_Cout) );
  logicunit logicunit_0 ( .A({DATA1[31:29], n367, DATA1[27:24], n366, 
        DATA1[22:16], n375, DATA1[14], n369, DATA1[12], n373, DATA1[10], n374, 
        DATA1[8], n370, DATA1[6], n372, DATA1[4], n376, DATA1[2], n371, n377}), 
        .B(DATA2), .SEL({\Sel[2] , n306, n306}), .LU_OUT(LU_out) );
  ComparatorUnit ComparatorUnit_0 ( .A_MSB(DATA1[31]), .B_MSB(DATA2[31]), 
        .SUBIN(OUT_adder), .COUT(Adder_Cout), .SIGN_UNSIGN(sign_unsign), .OP({
        n205, Comp_OP[1:0]}), .CU_OUT({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, SYNOPSYS_UNCONNECTED__22, 
        SYNOPSYS_UNCONNECTED__23, SYNOPSYS_UNCONNECTED__24, 
        SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, SYNOPSYS_UNCONNECTED__28, 
        SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, \CU_OUT[0] }) );
  shifter shifter_0 ( .R({DATA1[31:29], n367, DATA1[27:24], n366, DATA1[22:16], 
        n375, DATA1[14], n369, DATA1[12], n373, DATA1[10], n374, DATA1[8], 
        n370, DATA1[6], n372, DATA1[4], n376, DATA1[2], n371, n377}), .Offset(
        DATA2[4:0]), .Conf(Conf), .Shift_OUT(SHIFT_OUT) );
  INV_X1 U326 ( .A(n355), .ZN(n312) );
  NAND2_X1 U320 ( .A1(FUNC[1]), .A2(n355), .ZN(n310) );
  INV_X1 U240 ( .A(n313), .ZN(\Sel[2] ) );
  OAI21_X1 U239 ( .B1(n308), .B2(n313), .A(n314), .ZN(n104) );
  INV_X1 U322 ( .A(FUNC[0]), .ZN(n308) );
  NAND3_X1 U317 ( .A1(n353), .A2(FUNC[2]), .A3(FUNC[1]), .ZN(n358) );
  OAI22_X1 U238 ( .A1(FUNC[2]), .A2(n310), .B1(n311), .B2(n312), .ZN(
        sign_unsign) );
  NOR2_X1 U315 ( .A1(n308), .A2(n358), .ZN(Conf[1]) );
  NOR2_X1 U316 ( .A1(FUNC[0]), .A2(n358), .ZN(Conf[0]) );
  NOR2_X1 U308 ( .A1(n355), .A2(n205), .ZN(n309) );
  NAND2_X2 U235 ( .A1(n313), .A2(n314), .ZN(n317) );
  INV_X1 U325 ( .A(FUNC[1]), .ZN(n357) );
  NAND3_X1 U306 ( .A1(n353), .A2(n354), .A3(FUNC[1]), .ZN(n313) );
  NOR2_X1 U311 ( .A1(n354), .A2(FUNC[1]), .ZN(n352) );
  NAND4_X1 U323 ( .A1(FUNC[4]), .A2(n357), .A3(n354), .A4(n360), .ZN(n356) );
  INV_X1 U324 ( .A(FUNC[2]), .ZN(n354) );
  OAI21_X1 U237 ( .B1(n307), .B2(n308), .A(n309), .ZN(sub_add) );
  NAND3_X1 U313 ( .A1(n357), .A2(n354), .A3(n353), .ZN(n307) );
  NAND3_X1 U314 ( .A1(n353), .A2(FUNC[2]), .A3(FUNC[0]), .ZN(n359) );
  NAND2_X2 U234 ( .A1(n358), .A2(n359), .ZN(n318) );
  INV_X2 U236 ( .A(n307), .ZN(n316) );
  AOI22_X1 U312 ( .A1(SHIFT_OUT[0]), .A2(n318), .B1(OUT_adder[0]), .B2(n316), 
        .ZN(n349) );
  AOI222_X4 U232 ( .A1(OUT_adder[28]), .A2(n316), .B1(LU_out[28]), .B2(n317), 
        .C1(SHIFT_OUT[28]), .C2(n318), .ZN(n329) );
  CLKBUF_X1 U258 ( .A(OUT_adder[26]), .Z(n364) );
  OAI221_X1 U262 ( .B1(n361), .B2(n362), .C1(n363), .C2(n309), .A(n349), .ZN(
        OUTALU[0]) );
  INV_X1 U264 ( .A(LU_out[0]), .ZN(n361) );
  INV_X1 U268 ( .A(n317), .ZN(n362) );
  INV_X1 U272 ( .A(\CU_OUT[0] ), .ZN(n363) );
  CLKBUF_X1 U278 ( .A(OUT_adder[16]), .Z(n365) );
  AOI222_X4 U280 ( .A1(n364), .A2(n316), .B1(LU_out[26]), .B2(n317), .C1(
        SHIFT_OUT[26]), .C2(n318), .ZN(n331) );
  AOI222_X4 U290 ( .A1(n365), .A2(n316), .B1(LU_out[16]), .B2(n317), .C1(
        SHIFT_OUT[16]), .C2(n318), .ZN(n342) );
  CLKBUF_X1 U303 ( .A(DATA1[23]), .Z(n366) );
  BUF_X2 U304 ( .A(DATA1[28]), .Z(n367) );
  AOI222_X4 U307 ( .A1(OUT_adder[21]), .A2(n316), .B1(LU_out[21]), .B2(n317), 
        .C1(SHIFT_OUT[21]), .C2(n318), .ZN(n336) );
  AOI222_X4 U319 ( .A1(OUT_adder[29]), .A2(n316), .B1(LU_out[29]), .B2(n317), 
        .C1(SHIFT_OUT[29]), .C2(n318), .ZN(n328) );
  CLKBUF_X1 U329 ( .A(OUT_adder[30]), .Z(n379) );
  CLKBUF_X1 U330 ( .A(OUT_adder[3]), .Z(n368) );
  CLKBUF_X1 U331 ( .A(DATA1[13]), .Z(n369) );
  CLKBUF_X1 U332 ( .A(DATA1[7]), .Z(n370) );
  CLKBUF_X1 U333 ( .A(DATA1[1]), .Z(n371) );
  CLKBUF_X1 U334 ( .A(DATA1[5]), .Z(n372) );
  CLKBUF_X1 U335 ( .A(DATA1[11]), .Z(n373) );
  CLKBUF_X1 U336 ( .A(DATA1[9]), .Z(n374) );
  CLKBUF_X1 U337 ( .A(DATA1[15]), .Z(n375) );
  CLKBUF_X1 U338 ( .A(DATA1[3]), .Z(n376) );
  INV_X2 U339 ( .A(n310), .ZN(Comp_OP[1]) );
  CLKBUF_X1 U340 ( .A(DATA1[0]), .Z(n377) );
  AOI222_X4 U341 ( .A1(OUT_adder[24]), .A2(n316), .B1(LU_out[24]), .B2(n317), 
        .C1(SHIFT_OUT[24]), .C2(n318), .ZN(n333) );
  AOI222_X4 U342 ( .A1(OUT_adder[20]), .A2(n316), .B1(LU_out[20]), .B2(n317), 
        .C1(SHIFT_OUT[20]), .C2(n318), .ZN(n337) );
  CLKBUF_X1 U343 ( .A(OUT_adder[27]), .Z(n378) );
  AOI222_X4 U344 ( .A1(n379), .A2(n316), .B1(LU_out[30]), .B2(n317), .C1(
        SHIFT_OUT[30]), .C2(n318), .ZN(n326) );
  BUF_X8 U345 ( .A(sub_add), .Z(n305) );
endmodule


module P4addersub_N32 ( A, B, sub_add, Y, Cout );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input sub_add;
  output Cout;
  wire   net6007, net6009, net6012, net6021, net6024, n1, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n13, n14, n15, n16, n19, n21, n22, n25, n26,
         n38, n23, n24, n27, n28, n29, n30, n31, n32, n33, n34, n35, n43, n44,
         n45, n46, n47, n48, n49, n50, n51;
  wire   [31:0] B_subadd;
  wire   [7:1] carry;
  assign n23 = sub_add;
  assign n24 = A[5];
  assign n27 = A[19];
  assign n28 = A[9];
  assign n29 = A[11];
  assign n30 = A[28];
  assign n31 = A[23];
  assign n32 = A[7];
  assign n33 = A[3];
  assign n34 = A[13];
  assign n35 = A[15];

  XOR2_X1 U65 ( .A(n23), .B(B[13]), .Z(net6024) );
  XOR2_X1 U66 ( .A(n23), .B(B[23]), .Z(net6021) );
  XOR2_X1 U67 ( .A(n23), .B(B[7]), .Z(net6012) );
  XOR2_X1 U68 ( .A(n23), .B(B[11]), .Z(net6009) );
  XOR2_X1 U69 ( .A(n23), .B(B[15]), .Z(net6007) );
  XOR2_X1 U70 ( .A(n23), .B(B[17]), .Z(n9) );
  XOR2_X1 U71 ( .A(n23), .B(B[20]), .Z(n8) );
  XOR2_X1 U72 ( .A(n23), .B(B[1]), .Z(n7) );
  XOR2_X1 U73 ( .A(n23), .B(B[22]), .Z(n6) );
  XOR2_X1 U74 ( .A(n23), .B(B[8]), .Z(n5) );
  XOR2_X1 U75 ( .A(n23), .B(B[14]), .Z(n4) );
  XOR2_X1 U76 ( .A(n23), .B(B[0]), .Z(n38) );
  XOR2_X1 U77 ( .A(n23), .B(B[10]), .Z(n3) );
  XOR2_X1 U78 ( .A(n23), .B(B[19]), .Z(n26) );
  XOR2_X1 U79 ( .A(n23), .B(B[16]), .Z(n25) );
  XOR2_X1 U80 ( .A(n23), .B(B[5]), .Z(n22) );
  XOR2_X1 U81 ( .A(n23), .B(B[9]), .Z(n21) );
  XOR2_X1 U82 ( .A(n23), .B(B[6]), .Z(n2) );
  XOR2_X1 U83 ( .A(n23), .B(B[27]), .Z(n19) );
  XOR2_X1 U84 ( .A(n23), .B(B[3]), .Z(n16) );
  XOR2_X1 U85 ( .A(n23), .B(B[2]), .Z(n15) );
  XOR2_X1 U86 ( .A(n23), .B(B[24]), .Z(n14) );
  XOR2_X1 U87 ( .A(n23), .B(B[18]), .Z(n13) );
  XOR2_X1 U88 ( .A(n23), .B(B[21]), .Z(n11) );
  XOR2_X1 U89 ( .A(n23), .B(B[12]), .Z(n10) );
  XOR2_X1 U90 ( .A(n23), .B(B[28]), .Z(n1) );
  XOR2_X1 U91 ( .A(n23), .B(B[4]), .Z(B_subadd[4]) );
  XOR2_X1 U92 ( .A(n23), .B(B[31]), .Z(B_subadd[31]) );
  XOR2_X1 U93 ( .A(n23), .B(B[30]), .Z(B_subadd[30]) );
  XOR2_X1 U94 ( .A(n23), .B(B[29]), .Z(B_subadd[29]) );
  XOR2_X1 U95 ( .A(n23), .B(B[26]), .Z(B_subadd[26]) );
  XOR2_X1 U96 ( .A(n23), .B(B[25]), .Z(B_subadd[25]) );
  STCG_N32_L5 STCG_1 ( .A({A[31:29], n30, A[27:24], n31, A[22:20], n27, 
        A[18:16], n35, A[14], n34, A[12], n29, A[10], n28, A[8], n32, A[6], 
        n24, A[4], n33, A[2:0]}), .B({B_subadd[31:29], n1, n19, 
        B_subadd[26:25], n14, net6021, n6, n11, n8, n26, n13, n9, n25, net6007, 
        n4, net6024, n10, net6009, n3, n21, n5, net6012, n2, n22, B_subadd[4], 
        n16, n15, n7, n38}), .cin(n23), .cout({Cout, carry}) );
  sumgen_N_blocks8 sumgen_1 ( .A({A[31:29], n30, A[27:24], n31, A[22:20], n27, 
        A[18:16], n50, A[14], n46, A[12], n47, A[10], n45, A[8], n49, A[6], 
        n44, A[4], n48, A[2], n43, n51}), .B({B_subadd[31:29], n1, n19, 
        B_subadd[26:25], n14, net6021, n6, n11, n8, n26, n13, n9, n25, net6007, 
        n4, net6024, n10, net6009, n3, n21, n5, net6012, n2, n22, B_subadd[4], 
        n16, n15, n7, n38}), .Ci({carry, n23}), .S(Y) );
  BUF_X2 U97 ( .A(n28), .Z(n45) );
  CLKBUF_X1 U98 ( .A(A[1]), .Z(n43) );
  CLKBUF_X1 U99 ( .A(n24), .Z(n44) );
  CLKBUF_X1 U100 ( .A(n34), .Z(n46) );
  CLKBUF_X1 U101 ( .A(n29), .Z(n47) );
  BUF_X2 U102 ( .A(A[0]), .Z(n51) );
  CLKBUF_X1 U103 ( .A(n33), .Z(n48) );
  CLKBUF_X1 U104 ( .A(n32), .Z(n49) );
  CLKBUF_X1 U105 ( .A(n35), .Z(n50) );
endmodule


module HazardUnit_NUMBIT32_ADDRESS_WIDTH_RF5_OP_CODE_SIZE6 ( CLK, RST, RS1, 
        RS2, REGWRITE_DX, MEMREAD_DX, RD, OPCODE, STALL );
  input [4:0] RS1;
  input [4:0] RS2;
  input [4:0] RD;
  input [5:0] OPCODE;
  input CLK, RST, REGWRITE_DX, MEMREAD_DX;
  output STALL;
  wire   N9, N10, N11, N12, N13, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24;

  DFF_X1 \RD_DX_reg[4]  ( .D(N13), .CK(CLK), .QN(n6) );
  DFF_X1 \RD_DX_reg[3]  ( .D(N12), .CK(CLK), .QN(n5) );
  DFF_X1 \RD_DX_reg[2]  ( .D(N11), .CK(CLK), .QN(n9) );
  DFF_X1 \RD_DX_reg[1]  ( .D(N10), .CK(CLK), .QN(n8) );
  DFF_X1 \RD_DX_reg[0]  ( .D(N9), .CK(CLK), .QN(n7) );
  AND2_X1 U3 ( .A1(n3), .A2(n4), .ZN(n18) );
  XOR2_X1 U4 ( .A(n6), .B(RS1[4]), .Z(n3) );
  XOR2_X1 U5 ( .A(RS1[2]), .B(n9), .Z(n4) );
  AND4_X2 U6 ( .A1(n15), .A2(n16), .A3(n17), .A4(n18), .ZN(n12) );
  NAND2_X1 U7 ( .A1(n10), .A2(n11), .ZN(STALL) );
  NAND4_X1 U8 ( .A1(OPCODE[2]), .A2(n12), .A3(REGWRITE_DX), .A4(n13), .ZN(n11)
         );
  NOR4_X1 U9 ( .A1(OPCODE[5]), .A2(OPCODE[4]), .A3(OPCODE[3]), .A4(OPCODE[1]), 
        .ZN(n13) );
  OAI21_X1 U10 ( .B1(n14), .B2(n12), .A(MEMREAD_DX), .ZN(n10) );
  XOR2_X1 U11 ( .A(n7), .B(RS1[0]), .Z(n17) );
  XOR2_X1 U12 ( .A(n8), .B(RS1[1]), .Z(n16) );
  XOR2_X1 U13 ( .A(n5), .B(RS1[3]), .Z(n15) );
  NOR3_X1 U14 ( .A1(n19), .A2(n20), .A3(n21), .ZN(n14) );
  XNOR2_X1 U15 ( .A(n6), .B(RS2[4]), .ZN(n21) );
  XNOR2_X1 U16 ( .A(n9), .B(RS2[2]), .ZN(n20) );
  NAND3_X1 U17 ( .A1(n22), .A2(n23), .A3(n24), .ZN(n19) );
  XOR2_X1 U18 ( .A(n7), .B(RS2[0]), .Z(n24) );
  XOR2_X1 U19 ( .A(n8), .B(RS2[1]), .Z(n23) );
  XOR2_X1 U20 ( .A(n5), .B(RS2[3]), .Z(n22) );
  AND2_X1 U21 ( .A1(RST), .A2(RD[0]), .ZN(N9) );
  AND2_X1 U22 ( .A1(RD[4]), .A2(RST), .ZN(N13) );
  AND2_X1 U23 ( .A1(RD[3]), .A2(RST), .ZN(N12) );
  AND2_X1 U24 ( .A1(RD[2]), .A2(RST), .ZN(N11) );
  AND2_X1 U25 ( .A1(RD[1]), .A2(RST), .ZN(N10) );
endmodule


module BTB_PC_SIZE32_BTBSIZE5 ( Reset, Clk, Enable, PC_read, WR, PC_write, 
        SetT_NT, Set_target, OUT_PC_target, OUTT_NT, prevT_NT );
  input [31:0] PC_read;
  input [31:0] PC_write;
  input [31:0] Set_target;
  output [31:0] OUT_PC_target;
  input Reset, Clk, Enable, WR, SetT_NT;
  output OUTT_NT, prevT_NT;
  wire   \pc_target[2][31] , \pc_target[2][30] , \pc_target[2][29] ,
         \pc_target[2][28] , \pc_target[2][27] , \pc_target[2][26] ,
         \pc_target[2][25] , \pc_target[2][24] , \pc_target[2][23] ,
         \pc_target[2][22] , \pc_target[2][21] , \pc_target[2][20] ,
         \pc_target[2][19] , \pc_target[2][18] , \pc_target[2][17] ,
         \pc_target[2][16] , \pc_target[2][15] , \pc_target[2][14] ,
         \pc_target[2][13] , \pc_target[2][12] , \pc_target[2][11] ,
         \pc_target[2][10] , \pc_target[2][9] , \pc_target[2][8] ,
         \pc_target[2][7] , \pc_target[2][6] , \pc_target[2][5] ,
         \pc_target[2][4] , \pc_target[2][3] , \pc_target[2][2] ,
         \pc_target[2][1] , \pc_target[2][0] , \pc_target[3][31] ,
         \pc_target[3][30] , \pc_target[3][29] , \pc_target[3][28] ,
         \pc_target[3][27] , \pc_target[3][26] , \pc_target[3][25] ,
         \pc_target[3][24] , \pc_target[3][23] , \pc_target[3][22] ,
         \pc_target[3][21] , \pc_target[3][20] , \pc_target[3][19] ,
         \pc_target[3][18] , \pc_target[3][17] , \pc_target[3][16] ,
         \pc_target[3][15] , \pc_target[3][14] , \pc_target[3][13] ,
         \pc_target[3][12] , \pc_target[3][11] , \pc_target[3][10] ,
         \pc_target[3][9] , \pc_target[3][8] , \pc_target[3][7] ,
         \pc_target[3][6] , \pc_target[3][5] , \pc_target[3][4] ,
         \pc_target[3][3] , \pc_target[3][2] , \pc_target[3][1] ,
         \pc_target[3][0] , \pc_target[6][31] , \pc_target[6][30] ,
         \pc_target[6][29] , \pc_target[6][28] , \pc_target[6][27] ,
         \pc_target[6][26] , \pc_target[6][25] , \pc_target[6][24] ,
         \pc_target[6][23] , \pc_target[6][22] , \pc_target[6][21] ,
         \pc_target[6][20] , \pc_target[6][19] , \pc_target[6][18] ,
         \pc_target[6][17] , \pc_target[6][16] , \pc_target[6][15] ,
         \pc_target[6][14] , \pc_target[6][13] , \pc_target[6][12] ,
         \pc_target[6][11] , \pc_target[6][10] , \pc_target[6][9] ,
         \pc_target[6][8] , \pc_target[6][7] , \pc_target[6][6] ,
         \pc_target[6][5] , \pc_target[6][4] , \pc_target[6][3] ,
         \pc_target[6][2] , \pc_target[6][1] , \pc_target[6][0] ,
         \pc_target[7][31] , \pc_target[7][30] , \pc_target[7][29] ,
         \pc_target[7][28] , \pc_target[7][27] , \pc_target[7][26] ,
         \pc_target[7][25] , \pc_target[7][24] , \pc_target[7][23] ,
         \pc_target[7][22] , \pc_target[7][21] , \pc_target[7][20] ,
         \pc_target[7][19] , \pc_target[7][18] , \pc_target[7][17] ,
         \pc_target[7][16] , \pc_target[7][15] , \pc_target[7][14] ,
         \pc_target[7][13] , \pc_target[7][12] , \pc_target[7][11] ,
         \pc_target[7][10] , \pc_target[7][9] , \pc_target[7][8] ,
         \pc_target[7][7] , \pc_target[7][6] , \pc_target[7][5] ,
         \pc_target[7][4] , \pc_target[7][3] , \pc_target[7][2] ,
         \pc_target[7][1] , \pc_target[7][0] , \pc_target[10][31] ,
         \pc_target[10][30] , \pc_target[10][29] , \pc_target[10][28] ,
         \pc_target[10][27] , \pc_target[10][26] , \pc_target[10][25] ,
         \pc_target[10][24] , \pc_target[10][23] , \pc_target[10][22] ,
         \pc_target[10][21] , \pc_target[10][20] , \pc_target[10][19] ,
         \pc_target[10][18] , \pc_target[10][17] , \pc_target[10][16] ,
         \pc_target[10][15] , \pc_target[10][14] , \pc_target[10][13] ,
         \pc_target[10][12] , \pc_target[10][11] , \pc_target[10][10] ,
         \pc_target[10][9] , \pc_target[10][8] , \pc_target[10][7] ,
         \pc_target[10][6] , \pc_target[10][5] , \pc_target[10][4] ,
         \pc_target[10][3] , \pc_target[10][2] , \pc_target[10][1] ,
         \pc_target[10][0] , \pc_target[11][31] , \pc_target[11][30] ,
         \pc_target[11][29] , \pc_target[11][28] , \pc_target[11][27] ,
         \pc_target[11][26] , \pc_target[11][25] , \pc_target[11][24] ,
         \pc_target[11][23] , \pc_target[11][22] , \pc_target[11][21] ,
         \pc_target[11][20] , \pc_target[11][19] , \pc_target[11][18] ,
         \pc_target[11][17] , \pc_target[11][16] , \pc_target[11][15] ,
         \pc_target[11][14] , \pc_target[11][13] , \pc_target[11][12] ,
         \pc_target[11][11] , \pc_target[11][10] , \pc_target[11][9] ,
         \pc_target[11][8] , \pc_target[11][7] , \pc_target[11][6] ,
         \pc_target[11][5] , \pc_target[11][4] , \pc_target[11][3] ,
         \pc_target[11][2] , \pc_target[11][1] , \pc_target[11][0] ,
         \pc_target[14][31] , \pc_target[14][30] , \pc_target[14][29] ,
         \pc_target[14][28] , \pc_target[14][27] , \pc_target[14][26] ,
         \pc_target[14][25] , \pc_target[14][24] , \pc_target[14][23] ,
         \pc_target[14][22] , \pc_target[14][21] , \pc_target[14][20] ,
         \pc_target[14][19] , \pc_target[14][18] , \pc_target[14][17] ,
         \pc_target[14][16] , \pc_target[14][15] , \pc_target[14][14] ,
         \pc_target[14][13] , \pc_target[14][12] , \pc_target[14][11] ,
         \pc_target[14][10] , \pc_target[14][9] , \pc_target[14][8] ,
         \pc_target[14][7] , \pc_target[14][6] , \pc_target[14][5] ,
         \pc_target[14][4] , \pc_target[14][3] , \pc_target[14][2] ,
         \pc_target[14][1] , \pc_target[14][0] , \pc_target[15][31] ,
         \pc_target[15][30] , \pc_target[15][29] , \pc_target[15][28] ,
         \pc_target[15][27] , \pc_target[15][26] , \pc_target[15][25] ,
         \pc_target[15][24] , \pc_target[15][23] , \pc_target[15][22] ,
         \pc_target[15][21] , \pc_target[15][20] , \pc_target[15][19] ,
         \pc_target[15][18] , \pc_target[15][17] , \pc_target[15][16] ,
         \pc_target[15][15] , \pc_target[15][14] , \pc_target[15][13] ,
         \pc_target[15][12] , \pc_target[15][11] , \pc_target[15][10] ,
         \pc_target[15][9] , \pc_target[15][8] , \pc_target[15][7] ,
         \pc_target[15][6] , \pc_target[15][5] , \pc_target[15][4] ,
         \pc_target[15][3] , \pc_target[15][2] , \pc_target[15][1] ,
         \pc_target[15][0] , \pc_target[16][22] , \pc_target[18][31] ,
         \pc_target[18][30] , \pc_target[18][29] , \pc_target[18][28] ,
         \pc_target[18][27] , \pc_target[18][26] , \pc_target[18][25] ,
         \pc_target[18][24] , \pc_target[18][23] , \pc_target[18][22] ,
         \pc_target[18][21] , \pc_target[18][20] , \pc_target[18][19] ,
         \pc_target[18][18] , \pc_target[18][17] , \pc_target[18][16] ,
         \pc_target[18][15] , \pc_target[18][14] , \pc_target[18][13] ,
         \pc_target[18][12] , \pc_target[18][11] , \pc_target[18][10] ,
         \pc_target[18][9] , \pc_target[18][8] , \pc_target[18][7] ,
         \pc_target[18][6] , \pc_target[18][5] , \pc_target[18][4] ,
         \pc_target[18][3] , \pc_target[18][2] , \pc_target[18][1] ,
         \pc_target[18][0] , \pc_target[19][31] , \pc_target[19][30] ,
         \pc_target[19][29] , \pc_target[19][28] , \pc_target[19][27] ,
         \pc_target[19][26] , \pc_target[19][25] , \pc_target[19][24] ,
         \pc_target[19][23] , \pc_target[19][22] , \pc_target[19][21] ,
         \pc_target[19][20] , \pc_target[19][19] , \pc_target[19][18] ,
         \pc_target[19][17] , \pc_target[19][16] , \pc_target[19][15] ,
         \pc_target[19][14] , \pc_target[19][13] , \pc_target[19][12] ,
         \pc_target[19][11] , \pc_target[19][10] , \pc_target[19][9] ,
         \pc_target[19][8] , \pc_target[19][7] , \pc_target[19][6] ,
         \pc_target[19][5] , \pc_target[19][4] , \pc_target[19][3] ,
         \pc_target[19][2] , \pc_target[19][1] , \pc_target[19][0] ,
         \pc_target[20][31] , \pc_target[20][30] , \pc_target[20][29] ,
         \pc_target[20][28] , \pc_target[20][27] , \pc_target[20][26] ,
         \pc_target[20][25] , \pc_target[20][24] , \pc_target[20][23] ,
         \pc_target[20][22] , \pc_target[20][21] , \pc_target[20][20] ,
         \pc_target[20][19] , \pc_target[20][18] , \pc_target[20][17] ,
         \pc_target[20][16] , \pc_target[20][15] , \pc_target[20][14] ,
         \pc_target[20][13] , \pc_target[20][12] , \pc_target[20][11] ,
         \pc_target[20][10] , \pc_target[20][9] , \pc_target[20][8] ,
         \pc_target[20][7] , \pc_target[20][6] , \pc_target[20][5] ,
         \pc_target[20][4] , \pc_target[20][3] , \pc_target[20][2] ,
         \pc_target[20][1] , \pc_target[20][0] , \pc_target[21][31] ,
         \pc_target[21][30] , \pc_target[21][29] , \pc_target[21][28] ,
         \pc_target[21][27] , \pc_target[21][26] , \pc_target[21][25] ,
         \pc_target[21][24] , \pc_target[21][23] , \pc_target[21][22] ,
         \pc_target[21][21] , \pc_target[21][20] , \pc_target[21][19] ,
         \pc_target[21][18] , \pc_target[21][17] , \pc_target[21][16] ,
         \pc_target[21][15] , \pc_target[21][14] , \pc_target[21][13] ,
         \pc_target[21][12] , \pc_target[21][11] , \pc_target[21][10] ,
         \pc_target[21][9] , \pc_target[21][8] , \pc_target[21][7] ,
         \pc_target[21][6] , \pc_target[21][5] , \pc_target[21][4] ,
         \pc_target[21][3] , \pc_target[21][2] , \pc_target[21][1] ,
         \pc_target[21][0] , \pc_target[26][31] , \pc_target[26][30] ,
         \pc_target[26][29] , \pc_target[26][28] , \pc_target[26][27] ,
         \pc_target[26][26] , \pc_target[26][25] , \pc_target[26][24] ,
         \pc_target[26][23] , \pc_target[26][22] , \pc_target[26][21] ,
         \pc_target[26][20] , \pc_target[26][19] , \pc_target[26][18] ,
         \pc_target[26][17] , \pc_target[26][16] , \pc_target[26][15] ,
         \pc_target[26][14] , \pc_target[26][13] , \pc_target[26][12] ,
         \pc_target[26][11] , \pc_target[26][10] , \pc_target[26][9] ,
         \pc_target[26][8] , \pc_target[26][7] , \pc_target[26][6] ,
         \pc_target[26][5] , \pc_target[26][4] , \pc_target[26][3] ,
         \pc_target[26][2] , \pc_target[26][1] , \pc_target[26][0] ,
         \pc_target[27][31] , \pc_target[27][30] , \pc_target[27][29] ,
         \pc_target[27][28] , \pc_target[27][27] , \pc_target[27][26] ,
         \pc_target[27][25] , \pc_target[27][24] , \pc_target[27][23] ,
         \pc_target[27][22] , \pc_target[27][21] , \pc_target[27][20] ,
         \pc_target[27][19] , \pc_target[27][18] , \pc_target[27][17] ,
         \pc_target[27][16] , \pc_target[27][15] , \pc_target[27][14] ,
         \pc_target[27][13] , \pc_target[27][12] , \pc_target[27][11] ,
         \pc_target[27][10] , \pc_target[27][9] , \pc_target[27][8] ,
         \pc_target[27][7] , \pc_target[27][6] , \pc_target[27][5] ,
         \pc_target[27][4] , \pc_target[27][3] , \pc_target[27][2] ,
         \pc_target[27][1] , \pc_target[27][0] , \pc_target[30][31] ,
         \pc_target[30][30] , \pc_target[30][29] , \pc_target[30][28] ,
         \pc_target[30][27] , \pc_target[30][26] , \pc_target[30][25] ,
         \pc_target[30][24] , \pc_target[30][23] , \pc_target[30][22] ,
         \pc_target[30][21] , \pc_target[30][20] , \pc_target[30][19] ,
         \pc_target[30][18] , \pc_target[30][17] , \pc_target[30][16] ,
         \pc_target[30][15] , \pc_target[30][14] , \pc_target[30][13] ,
         \pc_target[30][12] , \pc_target[30][11] , \pc_target[30][10] ,
         \pc_target[30][9] , \pc_target[30][8] , \pc_target[30][7] ,
         \pc_target[30][6] , \pc_target[30][5] , \pc_target[30][4] ,
         \pc_target[30][3] , \pc_target[30][2] , \pc_target[30][1] ,
         \pc_target[30][0] , \pc_target[31][31] , \pc_target[31][30] ,
         \pc_target[31][29] , \pc_target[31][28] , \pc_target[31][27] ,
         \pc_target[31][26] , \pc_target[31][25] , \pc_target[31][24] ,
         \pc_target[31][23] , \pc_target[31][22] , \pc_target[31][21] ,
         \pc_target[31][20] , \pc_target[31][19] , \pc_target[31][18] ,
         \pc_target[31][17] , \pc_target[31][16] , \pc_target[31][15] ,
         \pc_target[31][14] , \pc_target[31][13] , \pc_target[31][12] ,
         \pc_target[31][11] , \pc_target[31][10] , \pc_target[31][9] ,
         \pc_target[31][8] , \pc_target[31][7] , \pc_target[31][6] ,
         \pc_target[31][5] , \pc_target[31][4] , \pc_target[31][3] ,
         \pc_target[31][2] , \pc_target[31][1] , \pc_target[31][0] , N96, N97,
         N98, N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N109,
         N110, N111, N112, N113, N114, N115, N116, N117, N118, N119, N120,
         N121, N122, N123, N124, N125, N126, N127, \pc_lut[2][31] ,
         \pc_lut[2][30] , \pc_lut[2][29] , \pc_lut[2][28] , \pc_lut[2][27] ,
         \pc_lut[2][26] , \pc_lut[2][25] , \pc_lut[2][24] , \pc_lut[2][23] ,
         \pc_lut[2][22] , \pc_lut[2][21] , \pc_lut[2][20] , \pc_lut[2][19] ,
         \pc_lut[2][18] , \pc_lut[2][17] , \pc_lut[2][16] , \pc_lut[2][15] ,
         \pc_lut[2][14] , \pc_lut[2][13] , \pc_lut[2][12] , \pc_lut[2][11] ,
         \pc_lut[2][10] , \pc_lut[2][9] , \pc_lut[2][8] , \pc_lut[2][7] ,
         \pc_lut[2][6] , \pc_lut[2][5] , \pc_lut[2][1] , \pc_lut[3][31] ,
         \pc_lut[3][30] , \pc_lut[3][29] , \pc_lut[3][28] , \pc_lut[3][27] ,
         \pc_lut[3][26] , \pc_lut[3][25] , \pc_lut[3][24] , \pc_lut[3][23] ,
         \pc_lut[3][22] , \pc_lut[3][21] , \pc_lut[3][20] , \pc_lut[3][19] ,
         \pc_lut[3][18] , \pc_lut[3][17] , \pc_lut[3][16] , \pc_lut[3][15] ,
         \pc_lut[3][14] , \pc_lut[3][13] , \pc_lut[3][12] , \pc_lut[3][11] ,
         \pc_lut[3][10] , \pc_lut[3][9] , \pc_lut[3][8] , \pc_lut[3][7] ,
         \pc_lut[3][6] , \pc_lut[3][5] , \pc_lut[3][1] , \pc_lut[3][0] ,
         \pc_lut[6][31] , \pc_lut[6][30] , \pc_lut[6][29] , \pc_lut[6][28] ,
         \pc_lut[6][27] , \pc_lut[6][26] , \pc_lut[6][25] , \pc_lut[6][24] ,
         \pc_lut[6][23] , \pc_lut[6][22] , \pc_lut[6][21] , \pc_lut[6][20] ,
         \pc_lut[6][19] , \pc_lut[6][18] , \pc_lut[6][17] , \pc_lut[6][16] ,
         \pc_lut[6][15] , \pc_lut[6][14] , \pc_lut[6][13] , \pc_lut[6][12] ,
         \pc_lut[6][11] , \pc_lut[6][10] , \pc_lut[6][9] , \pc_lut[6][8] ,
         \pc_lut[6][7] , \pc_lut[6][6] , \pc_lut[6][5] , \pc_lut[6][2] ,
         \pc_lut[6][1] , \pc_lut[7][31] , \pc_lut[7][30] , \pc_lut[7][29] ,
         \pc_lut[7][28] , \pc_lut[7][27] , \pc_lut[7][26] , \pc_lut[7][25] ,
         \pc_lut[7][24] , \pc_lut[7][23] , \pc_lut[7][22] , \pc_lut[7][21] ,
         \pc_lut[7][20] , \pc_lut[7][19] , \pc_lut[7][18] , \pc_lut[7][17] ,
         \pc_lut[7][16] , \pc_lut[7][15] , \pc_lut[7][14] , \pc_lut[7][13] ,
         \pc_lut[7][12] , \pc_lut[7][11] , \pc_lut[7][10] , \pc_lut[7][9] ,
         \pc_lut[7][8] , \pc_lut[7][7] , \pc_lut[7][6] , \pc_lut[7][5] ,
         \pc_lut[7][2] , \pc_lut[7][1] , \pc_lut[7][0] , \pc_lut[10][31] ,
         \pc_lut[10][30] , \pc_lut[10][29] , \pc_lut[10][28] ,
         \pc_lut[10][27] , \pc_lut[10][26] , \pc_lut[10][25] ,
         \pc_lut[10][24] , \pc_lut[10][23] , \pc_lut[10][22] ,
         \pc_lut[10][21] , \pc_lut[10][20] , \pc_lut[10][19] ,
         \pc_lut[10][18] , \pc_lut[10][17] , \pc_lut[10][16] ,
         \pc_lut[10][15] , \pc_lut[10][14] , \pc_lut[10][13] ,
         \pc_lut[10][12] , \pc_lut[10][11] , \pc_lut[10][10] , \pc_lut[10][9] ,
         \pc_lut[10][8] , \pc_lut[10][7] , \pc_lut[10][6] , \pc_lut[10][5] ,
         \pc_lut[10][3] , \pc_lut[10][1] , \pc_lut[11][31] , \pc_lut[11][30] ,
         \pc_lut[11][29] , \pc_lut[11][28] , \pc_lut[11][27] ,
         \pc_lut[11][26] , \pc_lut[11][25] , \pc_lut[11][24] ,
         \pc_lut[11][23] , \pc_lut[11][22] , \pc_lut[11][21] ,
         \pc_lut[11][20] , \pc_lut[11][19] , \pc_lut[11][18] ,
         \pc_lut[11][17] , \pc_lut[11][16] , \pc_lut[11][15] ,
         \pc_lut[11][14] , \pc_lut[11][13] , \pc_lut[11][12] ,
         \pc_lut[11][11] , \pc_lut[11][10] , \pc_lut[11][9] , \pc_lut[11][8] ,
         \pc_lut[11][7] , \pc_lut[11][6] , \pc_lut[11][5] , \pc_lut[11][3] ,
         \pc_lut[11][1] , \pc_lut[11][0] , \pc_lut[14][31] , \pc_lut[14][30] ,
         \pc_lut[14][29] , \pc_lut[14][28] , \pc_lut[14][27] ,
         \pc_lut[14][26] , \pc_lut[14][25] , \pc_lut[14][24] ,
         \pc_lut[14][23] , \pc_lut[14][22] , \pc_lut[14][21] ,
         \pc_lut[14][20] , \pc_lut[14][19] , \pc_lut[14][18] ,
         \pc_lut[14][17] , \pc_lut[14][16] , \pc_lut[14][15] ,
         \pc_lut[14][14] , \pc_lut[14][13] , \pc_lut[14][12] ,
         \pc_lut[14][11] , \pc_lut[14][10] , \pc_lut[14][9] , \pc_lut[14][8] ,
         \pc_lut[14][7] , \pc_lut[14][6] , \pc_lut[14][5] , \pc_lut[14][3] ,
         \pc_lut[14][2] , \pc_lut[14][1] , \pc_lut[15][31] , \pc_lut[15][30] ,
         \pc_lut[15][29] , \pc_lut[15][28] , \pc_lut[15][27] ,
         \pc_lut[15][26] , \pc_lut[15][25] , \pc_lut[15][24] ,
         \pc_lut[15][23] , \pc_lut[15][22] , \pc_lut[15][21] ,
         \pc_lut[15][20] , \pc_lut[15][19] , \pc_lut[15][18] ,
         \pc_lut[15][17] , \pc_lut[15][16] , \pc_lut[15][15] ,
         \pc_lut[15][14] , \pc_lut[15][13] , \pc_lut[15][12] ,
         \pc_lut[15][11] , \pc_lut[15][10] , \pc_lut[15][9] , \pc_lut[15][8] ,
         \pc_lut[15][7] , \pc_lut[15][6] , \pc_lut[15][5] , \pc_lut[15][3] ,
         \pc_lut[15][2] , \pc_lut[15][1] , \pc_lut[15][0] , \pc_lut[18][31] ,
         \pc_lut[18][30] , \pc_lut[18][29] , \pc_lut[18][28] ,
         \pc_lut[18][27] , \pc_lut[18][26] , \pc_lut[18][25] ,
         \pc_lut[18][24] , \pc_lut[18][23] , \pc_lut[18][22] ,
         \pc_lut[18][21] , \pc_lut[18][20] , \pc_lut[18][19] ,
         \pc_lut[18][18] , \pc_lut[18][17] , \pc_lut[18][16] ,
         \pc_lut[18][15] , \pc_lut[18][14] , \pc_lut[18][13] ,
         \pc_lut[18][12] , \pc_lut[18][11] , \pc_lut[18][10] , \pc_lut[18][9] ,
         \pc_lut[18][8] , \pc_lut[18][7] , \pc_lut[18][6] , \pc_lut[18][5] ,
         \pc_lut[18][4] , \pc_lut[18][1] , \pc_lut[19][31] , \pc_lut[19][30] ,
         \pc_lut[19][29] , \pc_lut[19][28] , \pc_lut[19][27] ,
         \pc_lut[19][26] , \pc_lut[19][25] , \pc_lut[19][24] ,
         \pc_lut[19][23] , \pc_lut[19][22] , \pc_lut[19][21] ,
         \pc_lut[19][20] , \pc_lut[19][19] , \pc_lut[19][18] ,
         \pc_lut[19][17] , \pc_lut[19][16] , \pc_lut[19][15] ,
         \pc_lut[19][14] , \pc_lut[19][13] , \pc_lut[19][12] ,
         \pc_lut[19][11] , \pc_lut[19][10] , \pc_lut[19][9] , \pc_lut[19][8] ,
         \pc_lut[19][7] , \pc_lut[19][6] , \pc_lut[19][5] , \pc_lut[19][4] ,
         \pc_lut[19][1] , \pc_lut[19][0] , \pc_lut[20][31] , \pc_lut[20][30] ,
         \pc_lut[20][29] , \pc_lut[20][28] , \pc_lut[20][27] ,
         \pc_lut[20][26] , \pc_lut[20][25] , \pc_lut[20][24] ,
         \pc_lut[20][23] , \pc_lut[20][22] , \pc_lut[20][21] ,
         \pc_lut[20][20] , \pc_lut[20][19] , \pc_lut[20][18] ,
         \pc_lut[20][17] , \pc_lut[20][16] , \pc_lut[20][15] ,
         \pc_lut[20][14] , \pc_lut[20][13] , \pc_lut[20][12] ,
         \pc_lut[20][11] , \pc_lut[20][10] , \pc_lut[20][9] , \pc_lut[20][8] ,
         \pc_lut[20][7] , \pc_lut[20][6] , \pc_lut[20][5] , \pc_lut[20][4] ,
         \pc_lut[20][2] , \pc_lut[21][31] , \pc_lut[21][30] , \pc_lut[21][29] ,
         \pc_lut[21][28] , \pc_lut[21][27] , \pc_lut[21][26] ,
         \pc_lut[21][25] , \pc_lut[21][24] , \pc_lut[21][23] ,
         \pc_lut[21][22] , \pc_lut[21][21] , \pc_lut[21][20] ,
         \pc_lut[21][19] , \pc_lut[21][18] , \pc_lut[21][17] ,
         \pc_lut[21][16] , \pc_lut[21][15] , \pc_lut[21][14] ,
         \pc_lut[21][13] , \pc_lut[21][12] , \pc_lut[21][11] ,
         \pc_lut[21][10] , \pc_lut[21][9] , \pc_lut[21][8] , \pc_lut[21][7] ,
         \pc_lut[21][6] , \pc_lut[21][5] , \pc_lut[21][4] , \pc_lut[21][2] ,
         \pc_lut[21][0] , \pc_lut[26][31] , \pc_lut[26][30] , \pc_lut[26][29] ,
         \pc_lut[26][28] , \pc_lut[26][27] , \pc_lut[26][26] ,
         \pc_lut[26][25] , \pc_lut[26][24] , \pc_lut[26][23] ,
         \pc_lut[26][22] , \pc_lut[26][21] , \pc_lut[26][20] ,
         \pc_lut[26][19] , \pc_lut[26][18] , \pc_lut[26][17] ,
         \pc_lut[26][16] , \pc_lut[26][15] , \pc_lut[26][14] ,
         \pc_lut[26][13] , \pc_lut[26][12] , \pc_lut[26][11] ,
         \pc_lut[26][10] , \pc_lut[26][9] , \pc_lut[26][8] , \pc_lut[26][7] ,
         \pc_lut[26][6] , \pc_lut[26][5] , \pc_lut[26][4] , \pc_lut[26][3] ,
         \pc_lut[26][1] , \pc_lut[27][31] , \pc_lut[27][30] , \pc_lut[27][29] ,
         \pc_lut[27][28] , \pc_lut[27][27] , \pc_lut[27][26] ,
         \pc_lut[27][25] , \pc_lut[27][24] , \pc_lut[27][23] ,
         \pc_lut[27][22] , \pc_lut[27][21] , \pc_lut[27][20] ,
         \pc_lut[27][19] , \pc_lut[27][18] , \pc_lut[27][17] ,
         \pc_lut[27][16] , \pc_lut[27][15] , \pc_lut[27][14] ,
         \pc_lut[27][13] , \pc_lut[27][12] , \pc_lut[27][11] ,
         \pc_lut[27][10] , \pc_lut[27][9] , \pc_lut[27][8] , \pc_lut[27][7] ,
         \pc_lut[27][6] , \pc_lut[27][5] , \pc_lut[27][4] , \pc_lut[27][3] ,
         \pc_lut[27][1] , \pc_lut[27][0] , \pc_lut[30][31] , \pc_lut[30][30] ,
         \pc_lut[30][29] , \pc_lut[30][28] , \pc_lut[30][27] ,
         \pc_lut[30][26] , \pc_lut[30][25] , \pc_lut[30][24] ,
         \pc_lut[30][23] , \pc_lut[30][22] , \pc_lut[30][21] ,
         \pc_lut[30][20] , \pc_lut[30][19] , \pc_lut[30][18] ,
         \pc_lut[30][17] , \pc_lut[30][16] , \pc_lut[30][15] ,
         \pc_lut[30][14] , \pc_lut[30][13] , \pc_lut[30][12] ,
         \pc_lut[30][11] , \pc_lut[30][10] , \pc_lut[30][9] , \pc_lut[30][8] ,
         \pc_lut[30][7] , \pc_lut[30][6] , \pc_lut[30][5] , \pc_lut[30][4] ,
         \pc_lut[30][3] , \pc_lut[30][2] , \pc_lut[30][1] , \pc_lut[31][31] ,
         \pc_lut[31][30] , \pc_lut[31][29] , \pc_lut[31][28] ,
         \pc_lut[31][27] , \pc_lut[31][26] , \pc_lut[31][25] ,
         \pc_lut[31][24] , \pc_lut[31][23] , \pc_lut[31][22] ,
         \pc_lut[31][21] , \pc_lut[31][20] , \pc_lut[31][19] ,
         \pc_lut[31][18] , \pc_lut[31][17] , \pc_lut[31][16] ,
         \pc_lut[31][15] , \pc_lut[31][14] , \pc_lut[31][13] ,
         \pc_lut[31][12] , \pc_lut[31][11] , \pc_lut[31][10] , \pc_lut[31][9] ,
         \pc_lut[31][8] , \pc_lut[31][7] , \pc_lut[31][6] , \pc_lut[31][5] ,
         \pc_lut[31][4] , \pc_lut[31][3] , \pc_lut[31][2] , \pc_lut[31][1] ,
         \pc_lut[31][0] , N188, N189, N190, N191, N192, N193, N194, N195, N196,
         N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207,
         N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218,
         N219, N220, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1257, n1258, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1393, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1497, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1657, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1791, n1792, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1825,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1927, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2014, n2015, n2016,
         n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
         n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
         n2058, n2059, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2092, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2191, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2386,
         n2389, n2391, n2392, n2394, n2397, n2399, n2400, n2401, n2404, n2405,
         n2406, n2407, n2412, n2413, n2414, n2415, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
         n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
         n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
         n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
         n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
         n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
         n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
         n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
         n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
         n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
         n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
         n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
         n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
         n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
         n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
         n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
         n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
         n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6721, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6818, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6913, n6914, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6946, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6977, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7072,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7104,
         n7105, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7136,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7233, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7296, n7297, n7298, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7328, n7330, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7360, n7361, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7392, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7425, n7426, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7458,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7489, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n2, n3,
         n283, n525, n558, n768, n802, n871, n973, n1240, n1256, n1259, n1275,
         n1292, n1293, n1344, n1392, n1394, n1426, n1427, n1428, n1446, n1463,
         n1481, n1496, n1498, n1611, n1656, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976;

  DFFR_X1 prevT_NTs_reg ( .D(OUTT_NT), .CK(Clk), .RN(n3894), .Q(prevT_NT) );
  DFFR_X1 \pc_lut_reg[0][31]  ( .D(n7537), .CK(Clk), .RN(n3895), .QN(n2241) );
  DFFR_X1 \pc_lut_reg[0][29]  ( .D(n7536), .CK(Clk), .RN(n3895), .QN(n2240) );
  DFFR_X1 \pc_lut_reg[0][27]  ( .D(n7535), .CK(Clk), .RN(n3895), .QN(n2239) );
  DFFR_X1 \pc_lut_reg[0][25]  ( .D(n7534), .CK(Clk), .RN(n3895), .QN(n2238) );
  DFFR_X1 \pc_lut_reg[0][23]  ( .D(n7533), .CK(Clk), .RN(n3895), .QN(n2237) );
  DFFR_X1 \pc_lut_reg[0][21]  ( .D(n7532), .CK(Clk), .RN(n3895), .QN(n2236) );
  DFFR_X1 \pc_lut_reg[0][19]  ( .D(n7531), .CK(Clk), .RN(n3895), .QN(n2235) );
  DFFR_X1 \pc_lut_reg[0][17]  ( .D(n7530), .CK(Clk), .RN(n3895), .QN(n2234) );
  DFFR_X1 \pc_lut_reg[0][15]  ( .D(n7529), .CK(Clk), .RN(n3895), .QN(n2233) );
  DFFR_X1 \pc_lut_reg[0][13]  ( .D(n7528), .CK(Clk), .RN(n3895), .QN(n2232) );
  DFFR_X1 \pc_lut_reg[0][11]  ( .D(n7527), .CK(Clk), .RN(n3895), .QN(n2231) );
  DFFR_X1 \pc_lut_reg[0][9]  ( .D(n7526), .CK(Clk), .RN(n3895), .QN(n2230) );
  DFFR_X1 \pc_lut_reg[0][7]  ( .D(n7525), .CK(Clk), .RN(n3895), .QN(n2229) );
  DFFR_X1 \pc_lut_reg[0][5]  ( .D(n7524), .CK(Clk), .RN(n3858), .QN(n2228) );
  DFFR_X1 \pc_lut_reg[0][6]  ( .D(n7518), .CK(Clk), .RN(n3895), .QN(n2222) );
  DFFR_X1 \pc_lut_reg[0][8]  ( .D(n7517), .CK(Clk), .RN(n3895), .QN(n2221) );
  DFFR_X1 \pc_lut_reg[0][10]  ( .D(n7516), .CK(Clk), .RN(n3896), .QN(n2220) );
  DFFR_X1 \pc_lut_reg[0][12]  ( .D(n7515), .CK(Clk), .RN(n3896), .QN(n2219) );
  DFFR_X1 \pc_lut_reg[0][14]  ( .D(n7514), .CK(Clk), .RN(n3896), .QN(n2218) );
  DFFR_X1 \pc_lut_reg[0][16]  ( .D(n7513), .CK(Clk), .RN(n3896), .QN(n2217) );
  DFFR_X1 \pc_lut_reg[0][18]  ( .D(n7512), .CK(Clk), .RN(n3861), .QN(n2216) );
  DFFR_X1 \pc_lut_reg[0][20]  ( .D(n7511), .CK(Clk), .RN(n3896), .QN(n2215) );
  DFFR_X1 \pc_lut_reg[0][22]  ( .D(n7510), .CK(Clk), .RN(n3896), .QN(n2214) );
  DFFR_X1 \pc_lut_reg[0][24]  ( .D(n7509), .CK(Clk), .RN(n3896), .QN(n2213) );
  DFFR_X1 \pc_lut_reg[0][26]  ( .D(n7508), .CK(Clk), .RN(n3916), .QN(n2212) );
  DFFR_X1 \pc_lut_reg[0][28]  ( .D(n7507), .CK(Clk), .RN(n3912), .QN(n2211) );
  DFFR_X1 \pc_lut_reg[0][30]  ( .D(n7506), .CK(Clk), .RN(n3912), .QN(n2209) );
  DFFR_X1 \pc_lut_reg[1][31]  ( .D(n7505), .CK(Clk), .RN(n3913), .QN(n2207) );
  DFFR_X1 \pc_lut_reg[1][29]  ( .D(n7504), .CK(Clk), .RN(n3913), .QN(n2206) );
  DFFR_X1 \pc_lut_reg[1][27]  ( .D(n7503), .CK(Clk), .RN(n3913), .QN(n2205) );
  DFFR_X1 \pc_lut_reg[1][25]  ( .D(n7502), .CK(Clk), .RN(n3913), .QN(n2204) );
  DFFR_X1 \pc_lut_reg[1][23]  ( .D(n7501), .CK(Clk), .RN(n3913), .QN(n2203) );
  DFFR_X1 \pc_lut_reg[1][21]  ( .D(n7500), .CK(Clk), .RN(n3913), .QN(n2202) );
  DFFR_X1 \pc_lut_reg[1][19]  ( .D(n7499), .CK(Clk), .RN(n3913), .QN(n2201) );
  DFFR_X1 \pc_lut_reg[1][17]  ( .D(n7498), .CK(Clk), .RN(n3913), .QN(n2200) );
  DFFR_X1 \pc_lut_reg[1][15]  ( .D(n7497), .CK(Clk), .RN(n3913), .QN(n2199) );
  DFFR_X1 \pc_lut_reg[1][13]  ( .D(n7496), .CK(Clk), .RN(n3913), .QN(n2198) );
  DFFR_X1 \pc_lut_reg[1][11]  ( .D(n7495), .CK(Clk), .RN(n3913), .QN(n2197) );
  DFFR_X1 \pc_lut_reg[1][9]  ( .D(n7494), .CK(Clk), .RN(n3913), .QN(n2196) );
  DFFR_X1 \pc_lut_reg[1][7]  ( .D(n7493), .CK(Clk), .RN(n3913), .QN(n2195) );
  DFFR_X1 \pc_lut_reg[1][5]  ( .D(n7492), .CK(Clk), .RN(n3858), .QN(n2194) );
  DFFR_X1 \pc_lut_reg[1][0]  ( .D(n7489), .CK(Clk), .RN(n3913), .QN(n2191) );
  DFFR_X1 \pc_lut_reg[1][6]  ( .D(n7486), .CK(Clk), .RN(n3913), .QN(n2188) );
  DFFR_X1 \pc_lut_reg[1][8]  ( .D(n7485), .CK(Clk), .RN(n3914), .QN(n2187) );
  DFFR_X1 \pc_lut_reg[1][10]  ( .D(n7484), .CK(Clk), .RN(n3914), .QN(n2186) );
  DFFR_X1 \pc_lut_reg[1][12]  ( .D(n7483), .CK(Clk), .RN(n3914), .QN(n2185) );
  DFFR_X1 \pc_lut_reg[1][14]  ( .D(n7482), .CK(Clk), .RN(n3914), .QN(n2184) );
  DFFR_X1 \pc_lut_reg[1][16]  ( .D(n7481), .CK(Clk), .RN(n3914), .QN(n2183) );
  DFFR_X1 \pc_lut_reg[1][18]  ( .D(n7480), .CK(Clk), .RN(n3861), .QN(n2182) );
  DFFR_X1 \pc_lut_reg[1][20]  ( .D(n7479), .CK(Clk), .RN(n3914), .QN(n2181) );
  DFFR_X1 \pc_lut_reg[1][22]  ( .D(n7478), .CK(Clk), .RN(n3914), .QN(n2180) );
  DFFR_X1 \pc_lut_reg[1][24]  ( .D(n7477), .CK(Clk), .RN(n3914), .QN(n2179) );
  DFFR_X1 \pc_lut_reg[1][26]  ( .D(n7476), .CK(Clk), .RN(n3914), .QN(n2178) );
  DFFR_X1 \pc_lut_reg[1][28]  ( .D(n7475), .CK(Clk), .RN(n3914), .QN(n2177) );
  DFFR_X1 \pc_lut_reg[1][30]  ( .D(n7474), .CK(Clk), .RN(n3914), .QN(n2175) );
  DFFR_X1 \pc_lut_reg[2][31]  ( .D(n7473), .CK(Clk), .RN(n3914), .Q(
        \pc_lut[2][31] ), .QN(n2173) );
  DFFR_X1 \pc_lut_reg[2][29]  ( .D(n7472), .CK(Clk), .RN(n3914), .Q(
        \pc_lut[2][29] ), .QN(n2172) );
  DFFR_X1 \pc_lut_reg[2][27]  ( .D(n7471), .CK(Clk), .RN(n3914), .Q(
        \pc_lut[2][27] ), .QN(n2171) );
  DFFR_X1 \pc_lut_reg[2][25]  ( .D(n7470), .CK(Clk), .RN(n3914), .Q(
        \pc_lut[2][25] ), .QN(n2170) );
  DFFR_X1 \pc_lut_reg[2][23]  ( .D(n7469), .CK(Clk), .RN(n3915), .Q(
        \pc_lut[2][23] ), .QN(n2169) );
  DFFR_X1 \pc_lut_reg[2][21]  ( .D(n7468), .CK(Clk), .RN(n3915), .Q(
        \pc_lut[2][21] ), .QN(n2168) );
  DFFR_X1 \pc_lut_reg[2][19]  ( .D(n7467), .CK(Clk), .RN(n3915), .Q(
        \pc_lut[2][19] ), .QN(n2167) );
  DFFR_X1 \pc_lut_reg[2][17]  ( .D(n7466), .CK(Clk), .RN(n3915), .Q(
        \pc_lut[2][17] ), .QN(n2166) );
  DFFR_X1 \pc_lut_reg[2][15]  ( .D(n7465), .CK(Clk), .RN(n3915), .Q(
        \pc_lut[2][15] ), .QN(n2165) );
  DFFR_X1 \pc_lut_reg[2][13]  ( .D(n7464), .CK(Clk), .RN(n3915), .Q(
        \pc_lut[2][13] ), .QN(n2164) );
  DFFR_X1 \pc_lut_reg[2][11]  ( .D(n7463), .CK(Clk), .RN(n3915), .Q(
        \pc_lut[2][11] ), .QN(n2163) );
  DFFR_X1 \pc_lut_reg[2][9]  ( .D(n7462), .CK(Clk), .RN(n3915), .Q(
        \pc_lut[2][9] ), .QN(n2162) );
  DFFR_X1 \pc_lut_reg[2][7]  ( .D(n7461), .CK(Clk), .RN(n3915), .Q(
        \pc_lut[2][7] ), .QN(n2161) );
  DFFR_X1 \pc_lut_reg[2][5]  ( .D(n7460), .CK(Clk), .RN(n3858), .Q(
        \pc_lut[2][5] ), .QN(n2160) );
  DFFR_X1 \pc_lut_reg[2][1]  ( .D(n7458), .CK(Clk), .RN(n3915), .Q(
        \pc_lut[2][1] ) );
  DFFR_X1 \pc_lut_reg[2][6]  ( .D(n7454), .CK(Clk), .RN(n3915), .Q(
        \pc_lut[2][6] ), .QN(n2158) );
  DFFR_X1 \pc_lut_reg[2][8]  ( .D(n7453), .CK(Clk), .RN(n3915), .Q(
        \pc_lut[2][8] ), .QN(n2157) );
  DFFR_X1 \pc_lut_reg[2][10]  ( .D(n7452), .CK(Clk), .RN(n3915), .Q(
        \pc_lut[2][10] ), .QN(n2156) );
  DFFR_X1 \pc_lut_reg[2][12]  ( .D(n7451), .CK(Clk), .RN(n3915), .Q(
        \pc_lut[2][12] ), .QN(n2155) );
  DFFR_X1 \pc_lut_reg[2][14]  ( .D(n7450), .CK(Clk), .RN(n3915), .Q(
        \pc_lut[2][14] ), .QN(n2154) );
  DFFR_X1 \pc_lut_reg[2][16]  ( .D(n7449), .CK(Clk), .RN(n3916), .Q(
        \pc_lut[2][16] ), .QN(n2153) );
  DFFR_X1 \pc_lut_reg[2][18]  ( .D(n7448), .CK(Clk), .RN(n3861), .Q(
        \pc_lut[2][18] ), .QN(n2152) );
  DFFR_X1 \pc_lut_reg[2][20]  ( .D(n7447), .CK(Clk), .RN(n3916), .Q(
        \pc_lut[2][20] ), .QN(n2151) );
  DFFR_X1 \pc_lut_reg[2][22]  ( .D(n7446), .CK(Clk), .RN(n3916), .Q(
        \pc_lut[2][22] ), .QN(n2150) );
  DFFR_X1 \pc_lut_reg[2][24]  ( .D(n7445), .CK(Clk), .RN(n3916), .Q(
        \pc_lut[2][24] ), .QN(n2149) );
  DFFR_X1 \pc_lut_reg[2][26]  ( .D(n7444), .CK(Clk), .RN(n3916), .Q(
        \pc_lut[2][26] ), .QN(n2148) );
  DFFR_X1 \pc_lut_reg[2][28]  ( .D(n7443), .CK(Clk), .RN(n3916), .Q(
        \pc_lut[2][28] ), .QN(n2147) );
  DFFR_X1 \pc_lut_reg[2][30]  ( .D(n7442), .CK(Clk), .RN(n3916), .Q(
        \pc_lut[2][30] ), .QN(n2145) );
  DFFR_X1 \pc_lut_reg[3][31]  ( .D(n7441), .CK(Clk), .RN(n3916), .Q(
        \pc_lut[3][31] ), .QN(n2140) );
  DFFR_X1 \pc_lut_reg[3][29]  ( .D(n7440), .CK(Clk), .RN(n3916), .Q(
        \pc_lut[3][29] ), .QN(n2139) );
  DFFR_X1 \pc_lut_reg[3][27]  ( .D(n7439), .CK(Clk), .RN(n3916), .Q(
        \pc_lut[3][27] ), .QN(n2138) );
  DFFR_X1 \pc_lut_reg[3][25]  ( .D(n7438), .CK(Clk), .RN(n3916), .Q(
        \pc_lut[3][25] ), .QN(n2137) );
  DFFR_X1 \pc_lut_reg[3][23]  ( .D(n7437), .CK(Clk), .RN(n3916), .Q(
        \pc_lut[3][23] ), .QN(n2136) );
  DFFR_X1 \pc_lut_reg[3][21]  ( .D(n7436), .CK(Clk), .RN(n3916), .Q(
        \pc_lut[3][21] ), .QN(n2135) );
  DFFR_X1 \pc_lut_reg[3][19]  ( .D(n7435), .CK(Clk), .RN(n3916), .Q(
        \pc_lut[3][19] ), .QN(n2134) );
  DFFR_X1 \pc_lut_reg[3][17]  ( .D(n7434), .CK(Clk), .RN(n3917), .Q(
        \pc_lut[3][17] ), .QN(n2133) );
  DFFR_X1 \pc_lut_reg[3][15]  ( .D(n7433), .CK(Clk), .RN(n3917), .Q(
        \pc_lut[3][15] ), .QN(n2132) );
  DFFR_X1 \pc_lut_reg[3][13]  ( .D(n7432), .CK(Clk), .RN(n3917), .Q(
        \pc_lut[3][13] ), .QN(n2131) );
  DFFR_X1 \pc_lut_reg[3][11]  ( .D(n7431), .CK(Clk), .RN(n3917), .Q(
        \pc_lut[3][11] ), .QN(n2130) );
  DFFR_X1 \pc_lut_reg[3][9]  ( .D(n7430), .CK(Clk), .RN(n3917), .Q(
        \pc_lut[3][9] ), .QN(n2129) );
  DFFR_X1 \pc_lut_reg[3][7]  ( .D(n7429), .CK(Clk), .RN(n3917), .Q(
        \pc_lut[3][7] ), .QN(n2128) );
  DFFR_X1 \pc_lut_reg[3][5]  ( .D(n7428), .CK(Clk), .RN(n3858), .Q(
        \pc_lut[3][5] ), .QN(n2127) );
  DFFR_X1 \pc_lut_reg[3][1]  ( .D(n7426), .CK(Clk), .RN(n3917), .Q(
        \pc_lut[3][1] ) );
  DFFR_X1 \pc_lut_reg[3][0]  ( .D(n7425), .CK(Clk), .RN(n3917), .Q(
        \pc_lut[3][0] ) );
  DFFR_X1 \pc_lut_reg[3][6]  ( .D(n7422), .CK(Clk), .RN(n3917), .Q(
        \pc_lut[3][6] ), .QN(n2124) );
  DFFR_X1 \pc_lut_reg[3][8]  ( .D(n7421), .CK(Clk), .RN(n3917), .Q(
        \pc_lut[3][8] ), .QN(n2123) );
  DFFR_X1 \pc_lut_reg[3][10]  ( .D(n7420), .CK(Clk), .RN(n3917), .Q(
        \pc_lut[3][10] ), .QN(n2122) );
  DFFR_X1 \pc_lut_reg[3][12]  ( .D(n7419), .CK(Clk), .RN(n3917), .Q(
        \pc_lut[3][12] ), .QN(n2121) );
  DFFR_X1 \pc_lut_reg[3][14]  ( .D(n7418), .CK(Clk), .RN(n3917), .Q(
        \pc_lut[3][14] ), .QN(n2120) );
  DFFR_X1 \pc_lut_reg[3][16]  ( .D(n7417), .CK(Clk), .RN(n3917), .Q(
        \pc_lut[3][16] ), .QN(n2119) );
  DFFR_X1 \pc_lut_reg[3][18]  ( .D(n7416), .CK(Clk), .RN(n3861), .Q(
        \pc_lut[3][18] ), .QN(n2118) );
  DFFR_X1 \pc_lut_reg[3][20]  ( .D(n7415), .CK(Clk), .RN(n3917), .Q(
        \pc_lut[3][20] ), .QN(n2117) );
  DFFR_X1 \pc_lut_reg[3][22]  ( .D(n7414), .CK(Clk), .RN(n3918), .Q(
        \pc_lut[3][22] ), .QN(n2116) );
  DFFR_X1 \pc_lut_reg[3][24]  ( .D(n7413), .CK(Clk), .RN(n3918), .Q(
        \pc_lut[3][24] ), .QN(n2115) );
  DFFR_X1 \pc_lut_reg[3][26]  ( .D(n7412), .CK(Clk), .RN(n3918), .Q(
        \pc_lut[3][26] ), .QN(n2114) );
  DFFR_X1 \pc_lut_reg[3][28]  ( .D(n7411), .CK(Clk), .RN(n3918), .Q(
        \pc_lut[3][28] ), .QN(n2113) );
  DFFR_X1 \pc_lut_reg[3][30]  ( .D(n7410), .CK(Clk), .RN(n3918), .Q(
        \pc_lut[3][30] ), .QN(n2111) );
  DFFR_X1 \pc_lut_reg[4][31]  ( .D(n7409), .CK(Clk), .RN(n3918), .QN(n2109) );
  DFFR_X1 \pc_lut_reg[4][29]  ( .D(n7408), .CK(Clk), .RN(n3918), .QN(n2108) );
  DFFR_X1 \pc_lut_reg[4][27]  ( .D(n7407), .CK(Clk), .RN(n3918), .QN(n2107) );
  DFFR_X1 \pc_lut_reg[4][25]  ( .D(n7406), .CK(Clk), .RN(n3918), .QN(n2106) );
  DFFR_X1 \pc_lut_reg[4][23]  ( .D(n7405), .CK(Clk), .RN(n3918), .QN(n2105) );
  DFFR_X1 \pc_lut_reg[4][21]  ( .D(n7404), .CK(Clk), .RN(n3918), .QN(n2104) );
  DFFR_X1 \pc_lut_reg[4][19]  ( .D(n7403), .CK(Clk), .RN(n3918), .QN(n2103) );
  DFFR_X1 \pc_lut_reg[4][17]  ( .D(n7402), .CK(Clk), .RN(n3918), .QN(n2102) );
  DFFR_X1 \pc_lut_reg[4][15]  ( .D(n7401), .CK(Clk), .RN(n3918), .QN(n2101) );
  DFFR_X1 \pc_lut_reg[4][13]  ( .D(n7400), .CK(Clk), .RN(n3918), .QN(n2100) );
  DFFR_X1 \pc_lut_reg[4][11]  ( .D(n7399), .CK(Clk), .RN(n3919), .QN(n2099) );
  DFFR_X1 \pc_lut_reg[4][9]  ( .D(n7398), .CK(Clk), .RN(n3919), .QN(n2098) );
  DFFR_X1 \pc_lut_reg[4][7]  ( .D(n7397), .CK(Clk), .RN(n3919), .QN(n2097) );
  DFFR_X1 \pc_lut_reg[4][5]  ( .D(n7396), .CK(Clk), .RN(n3859), .QN(n2096) );
  DFFR_X1 \pc_lut_reg[4][2]  ( .D(n7392), .CK(Clk), .RN(n3919), .QN(n2092) );
  DFFR_X1 \pc_lut_reg[4][6]  ( .D(n7390), .CK(Clk), .RN(n3919), .QN(n2090) );
  DFFR_X1 \pc_lut_reg[4][8]  ( .D(n7389), .CK(Clk), .RN(n3919), .QN(n2089) );
  DFFR_X1 \pc_lut_reg[4][10]  ( .D(n7388), .CK(Clk), .RN(n3919), .QN(n2088) );
  DFFR_X1 \pc_lut_reg[4][12]  ( .D(n7387), .CK(Clk), .RN(n3919), .QN(n2087) );
  DFFR_X1 \pc_lut_reg[4][14]  ( .D(n7386), .CK(Clk), .RN(n3919), .QN(n2086) );
  DFFR_X1 \pc_lut_reg[4][16]  ( .D(n7385), .CK(Clk), .RN(n3919), .QN(n2085) );
  DFFR_X1 \pc_lut_reg[4][18]  ( .D(n7384), .CK(Clk), .RN(n3862), .QN(n2084) );
  DFFR_X1 \pc_lut_reg[4][20]  ( .D(n7383), .CK(Clk), .RN(n3919), .QN(n2083) );
  DFFR_X1 \pc_lut_reg[4][22]  ( .D(n7382), .CK(Clk), .RN(n3919), .QN(n2082) );
  DFFR_X1 \pc_lut_reg[4][24]  ( .D(n7381), .CK(Clk), .RN(n3919), .QN(n2081) );
  DFFR_X1 \pc_lut_reg[4][26]  ( .D(n7380), .CK(Clk), .RN(n3919), .QN(n2080) );
  DFFR_X1 \pc_lut_reg[4][28]  ( .D(n7379), .CK(Clk), .RN(n3920), .QN(n2079) );
  DFFR_X1 \pc_lut_reg[4][30]  ( .D(n7378), .CK(Clk), .RN(n3920), .QN(n2077) );
  DFFR_X1 \pc_lut_reg[5][31]  ( .D(n7377), .CK(Clk), .RN(n3919), .QN(n2075) );
  DFFR_X1 \pc_lut_reg[5][29]  ( .D(n7376), .CK(Clk), .RN(n3920), .QN(n2074) );
  DFFR_X1 \pc_lut_reg[5][27]  ( .D(n7375), .CK(Clk), .RN(n3920), .QN(n2073) );
  DFFR_X1 \pc_lut_reg[5][25]  ( .D(n7374), .CK(Clk), .RN(n3920), .QN(n2072) );
  DFFR_X1 \pc_lut_reg[5][23]  ( .D(n7373), .CK(Clk), .RN(n3920), .QN(n2071) );
  DFFR_X1 \pc_lut_reg[5][21]  ( .D(n7372), .CK(Clk), .RN(n3920), .QN(n2070) );
  DFFR_X1 \pc_lut_reg[5][19]  ( .D(n7371), .CK(Clk), .RN(n3920), .QN(n2069) );
  DFFR_X1 \pc_lut_reg[5][17]  ( .D(n7370), .CK(Clk), .RN(n3920), .QN(n2068) );
  DFFR_X1 \pc_lut_reg[5][15]  ( .D(n7369), .CK(Clk), .RN(n3920), .QN(n2067) );
  DFFR_X1 \pc_lut_reg[5][13]  ( .D(n7368), .CK(Clk), .RN(n3920), .QN(n2066) );
  DFFR_X1 \pc_lut_reg[5][11]  ( .D(n7367), .CK(Clk), .RN(n3920), .QN(n2065) );
  DFFR_X1 \pc_lut_reg[5][9]  ( .D(n7366), .CK(Clk), .RN(n3920), .QN(n2064) );
  DFFR_X1 \pc_lut_reg[5][7]  ( .D(n7365), .CK(Clk), .RN(n3920), .QN(n2063) );
  DFFR_X1 \pc_lut_reg[5][5]  ( .D(n7364), .CK(Clk), .RN(n3859), .QN(n2062) );
  DFFR_X1 \pc_lut_reg[5][0]  ( .D(n7361), .CK(Clk), .RN(n3920), .QN(n2059) );
  DFFR_X1 \pc_lut_reg[5][2]  ( .D(n7360), .CK(Clk), .RN(n3908), .QN(n2058) );
  DFFR_X1 \pc_lut_reg[5][6]  ( .D(n7358), .CK(Clk), .RN(n3904), .QN(n2056) );
  DFFR_X1 \pc_lut_reg[5][8]  ( .D(n7357), .CK(Clk), .RN(n3904), .QN(n2055) );
  DFFR_X1 \pc_lut_reg[5][10]  ( .D(n7356), .CK(Clk), .RN(n3904), .QN(n2054) );
  DFFR_X1 \pc_lut_reg[5][12]  ( .D(n7355), .CK(Clk), .RN(n3904), .QN(n2053) );
  DFFR_X1 \pc_lut_reg[5][14]  ( .D(n7354), .CK(Clk), .RN(n3904), .QN(n2052) );
  DFFR_X1 \pc_lut_reg[5][16]  ( .D(n7353), .CK(Clk), .RN(n3905), .QN(n2051) );
  DFFR_X1 \pc_lut_reg[5][18]  ( .D(n7352), .CK(Clk), .RN(n3862), .QN(n2050) );
  DFFR_X1 \pc_lut_reg[5][20]  ( .D(n7351), .CK(Clk), .RN(n3905), .QN(n2049) );
  DFFR_X1 \pc_lut_reg[5][22]  ( .D(n7350), .CK(Clk), .RN(n3905), .QN(n2048) );
  DFFR_X1 \pc_lut_reg[5][24]  ( .D(n7349), .CK(Clk), .RN(n3905), .QN(n2047) );
  DFFR_X1 \pc_lut_reg[5][26]  ( .D(n7348), .CK(Clk), .RN(n3905), .QN(n2046) );
  DFFR_X1 \pc_lut_reg[5][28]  ( .D(n7347), .CK(Clk), .RN(n3905), .QN(n2045) );
  DFFR_X1 \pc_lut_reg[5][30]  ( .D(n7346), .CK(Clk), .RN(n3905), .QN(n2043) );
  DFFR_X1 \pc_lut_reg[6][31]  ( .D(n7345), .CK(Clk), .RN(n3905), .Q(
        \pc_lut[6][31] ), .QN(n2041) );
  DFFR_X1 \pc_lut_reg[6][29]  ( .D(n7344), .CK(Clk), .RN(n3905), .Q(
        \pc_lut[6][29] ), .QN(n2040) );
  DFFR_X1 \pc_lut_reg[6][27]  ( .D(n7343), .CK(Clk), .RN(n3905), .Q(
        \pc_lut[6][27] ), .QN(n2039) );
  DFFR_X1 \pc_lut_reg[6][25]  ( .D(n7342), .CK(Clk), .RN(n3905), .Q(
        \pc_lut[6][25] ), .QN(n2038) );
  DFFR_X1 \pc_lut_reg[6][23]  ( .D(n7341), .CK(Clk), .RN(n3905), .Q(
        \pc_lut[6][23] ), .QN(n2037) );
  DFFR_X1 \pc_lut_reg[6][21]  ( .D(n7340), .CK(Clk), .RN(n3905), .Q(
        \pc_lut[6][21] ), .QN(n2036) );
  DFFR_X1 \pc_lut_reg[6][19]  ( .D(n7339), .CK(Clk), .RN(n3905), .Q(
        \pc_lut[6][19] ), .QN(n2035) );
  DFFR_X1 \pc_lut_reg[6][17]  ( .D(n7338), .CK(Clk), .RN(n3905), .Q(
        \pc_lut[6][17] ), .QN(n2034) );
  DFFR_X1 \pc_lut_reg[6][15]  ( .D(n7337), .CK(Clk), .RN(n3906), .Q(
        \pc_lut[6][15] ), .QN(n2033) );
  DFFR_X1 \pc_lut_reg[6][13]  ( .D(n7336), .CK(Clk), .RN(n3906), .Q(
        \pc_lut[6][13] ), .QN(n2032) );
  DFFR_X1 \pc_lut_reg[6][11]  ( .D(n7335), .CK(Clk), .RN(n3906), .Q(
        \pc_lut[6][11] ), .QN(n2031) );
  DFFR_X1 \pc_lut_reg[6][9]  ( .D(n7334), .CK(Clk), .RN(n3906), .Q(
        \pc_lut[6][9] ), .QN(n2030) );
  DFFR_X1 \pc_lut_reg[6][7]  ( .D(n7333), .CK(Clk), .RN(n3906), .Q(
        \pc_lut[6][7] ), .QN(n2029) );
  DFFR_X1 \pc_lut_reg[6][5]  ( .D(n7332), .CK(Clk), .RN(n3859), .Q(
        \pc_lut[6][5] ), .QN(n2028) );
  DFFR_X1 \pc_lut_reg[6][1]  ( .D(n7330), .CK(Clk), .RN(n3906), .Q(
        \pc_lut[6][1] ) );
  DFFR_X1 \pc_lut_reg[6][2]  ( .D(n7328), .CK(Clk), .RN(n3906), .Q(
        \pc_lut[6][2] ) );
  DFFR_X1 \pc_lut_reg[6][6]  ( .D(n7326), .CK(Clk), .RN(n3906), .Q(
        \pc_lut[6][6] ), .QN(n2025) );
  DFFR_X1 \pc_lut_reg[6][8]  ( .D(n7325), .CK(Clk), .RN(n3906), .Q(
        \pc_lut[6][8] ), .QN(n2024) );
  DFFR_X1 \pc_lut_reg[6][10]  ( .D(n7324), .CK(Clk), .RN(n3906), .Q(
        \pc_lut[6][10] ), .QN(n2023) );
  DFFR_X1 \pc_lut_reg[6][12]  ( .D(n7323), .CK(Clk), .RN(n3906), .Q(
        \pc_lut[6][12] ), .QN(n2022) );
  DFFR_X1 \pc_lut_reg[6][14]  ( .D(n7322), .CK(Clk), .RN(n3906), .Q(
        \pc_lut[6][14] ), .QN(n2021) );
  DFFR_X1 \pc_lut_reg[6][16]  ( .D(n7321), .CK(Clk), .RN(n3906), .Q(
        \pc_lut[6][16] ), .QN(n2020) );
  DFFR_X1 \pc_lut_reg[6][18]  ( .D(n7320), .CK(Clk), .RN(n3862), .Q(
        \pc_lut[6][18] ), .QN(n2019) );
  DFFR_X1 \pc_lut_reg[6][20]  ( .D(n7319), .CK(Clk), .RN(n3906), .Q(
        \pc_lut[6][20] ), .QN(n2018) );
  DFFR_X1 \pc_lut_reg[6][22]  ( .D(n7318), .CK(Clk), .RN(n3906), .Q(
        \pc_lut[6][22] ), .QN(n2017) );
  DFFR_X1 \pc_lut_reg[6][24]  ( .D(n7317), .CK(Clk), .RN(n3907), .Q(
        \pc_lut[6][24] ), .QN(n2016) );
  DFFR_X1 \pc_lut_reg[6][26]  ( .D(n7316), .CK(Clk), .RN(n3907), .Q(
        \pc_lut[6][26] ), .QN(n2015) );
  DFFR_X1 \pc_lut_reg[6][28]  ( .D(n7315), .CK(Clk), .RN(n3907), .Q(
        \pc_lut[6][28] ), .QN(n2014) );
  DFFR_X1 \pc_lut_reg[6][30]  ( .D(n7314), .CK(Clk), .RN(n3907), .Q(
        \pc_lut[6][30] ), .QN(n2012) );
  DFFR_X1 \pc_lut_reg[7][31]  ( .D(n7313), .CK(Clk), .RN(n3907), .Q(
        \pc_lut[7][31] ), .QN(n2009) );
  DFFR_X1 \pc_lut_reg[7][29]  ( .D(n7312), .CK(Clk), .RN(n3907), .Q(
        \pc_lut[7][29] ), .QN(n2008) );
  DFFR_X1 \pc_lut_reg[7][27]  ( .D(n7311), .CK(Clk), .RN(n3907), .Q(
        \pc_lut[7][27] ), .QN(n2007) );
  DFFR_X1 \pc_lut_reg[7][25]  ( .D(n7310), .CK(Clk), .RN(n3907), .Q(
        \pc_lut[7][25] ), .QN(n2006) );
  DFFR_X1 \pc_lut_reg[7][23]  ( .D(n7309), .CK(Clk), .RN(n3907), .Q(
        \pc_lut[7][23] ), .QN(n2005) );
  DFFR_X1 \pc_lut_reg[7][21]  ( .D(n7308), .CK(Clk), .RN(n3907), .Q(
        \pc_lut[7][21] ), .QN(n2004) );
  DFFR_X1 \pc_lut_reg[7][19]  ( .D(n7307), .CK(Clk), .RN(n3907), .Q(
        \pc_lut[7][19] ), .QN(n2003) );
  DFFR_X1 \pc_lut_reg[7][17]  ( .D(n7306), .CK(Clk), .RN(n3907), .Q(
        \pc_lut[7][17] ), .QN(n2002) );
  DFFR_X1 \pc_lut_reg[7][15]  ( .D(n7305), .CK(Clk), .RN(n3907), .Q(
        \pc_lut[7][15] ), .QN(n2001) );
  DFFR_X1 \pc_lut_reg[7][13]  ( .D(n7304), .CK(Clk), .RN(n3907), .Q(
        \pc_lut[7][13] ), .QN(n2000) );
  DFFR_X1 \pc_lut_reg[7][11]  ( .D(n7303), .CK(Clk), .RN(n3907), .Q(
        \pc_lut[7][11] ), .QN(n1999) );
  DFFR_X1 \pc_lut_reg[7][9]  ( .D(n7302), .CK(Clk), .RN(n3908), .Q(
        \pc_lut[7][9] ), .QN(n1998) );
  DFFR_X1 \pc_lut_reg[7][7]  ( .D(n7301), .CK(Clk), .RN(n3908), .Q(
        \pc_lut[7][7] ), .QN(n1997) );
  DFFR_X1 \pc_lut_reg[7][5]  ( .D(n7300), .CK(Clk), .RN(n3859), .Q(
        \pc_lut[7][5] ), .QN(n1996) );
  DFFR_X1 \pc_lut_reg[7][1]  ( .D(n7298), .CK(Clk), .RN(n3908), .Q(
        \pc_lut[7][1] ) );
  DFFR_X1 \pc_lut_reg[7][0]  ( .D(n7297), .CK(Clk), .RN(n3908), .Q(
        \pc_lut[7][0] ) );
  DFFR_X1 \pc_lut_reg[7][2]  ( .D(n7296), .CK(Clk), .RN(n3908), .Q(
        \pc_lut[7][2] ) );
  DFFR_X1 \pc_lut_reg[7][6]  ( .D(n7294), .CK(Clk), .RN(n3908), .Q(
        \pc_lut[7][6] ), .QN(n1992) );
  DFFR_X1 \pc_lut_reg[7][8]  ( .D(n7293), .CK(Clk), .RN(n3908), .Q(
        \pc_lut[7][8] ), .QN(n1991) );
  DFFR_X1 \pc_lut_reg[7][10]  ( .D(n7292), .CK(Clk), .RN(n3908), .Q(
        \pc_lut[7][10] ), .QN(n1990) );
  DFFR_X1 \pc_lut_reg[7][12]  ( .D(n7291), .CK(Clk), .RN(n3897), .Q(
        \pc_lut[7][12] ), .QN(n1989) );
  DFFR_X1 \pc_lut_reg[7][14]  ( .D(n7290), .CK(Clk), .RN(n3897), .Q(
        \pc_lut[7][14] ), .QN(n1988) );
  DFFR_X1 \pc_lut_reg[7][16]  ( .D(n7289), .CK(Clk), .RN(n3897), .Q(
        \pc_lut[7][16] ), .QN(n1987) );
  DFFR_X1 \pc_lut_reg[7][18]  ( .D(n7288), .CK(Clk), .RN(n3862), .Q(
        \pc_lut[7][18] ), .QN(n1986) );
  DFFR_X1 \pc_lut_reg[7][20]  ( .D(n7287), .CK(Clk), .RN(n3897), .Q(
        \pc_lut[7][20] ), .QN(n1985) );
  DFFR_X1 \pc_lut_reg[7][22]  ( .D(n7286), .CK(Clk), .RN(n3897), .Q(
        \pc_lut[7][22] ), .QN(n1984) );
  DFFR_X1 \pc_lut_reg[7][24]  ( .D(n7285), .CK(Clk), .RN(n3897), .Q(
        \pc_lut[7][24] ), .QN(n1983) );
  DFFR_X1 \pc_lut_reg[7][26]  ( .D(n7284), .CK(Clk), .RN(n3897), .Q(
        \pc_lut[7][26] ), .QN(n1982) );
  DFFR_X1 \pc_lut_reg[7][28]  ( .D(n7283), .CK(Clk), .RN(n3897), .Q(
        \pc_lut[7][28] ), .QN(n1981) );
  DFFR_X1 \pc_lut_reg[7][30]  ( .D(n7282), .CK(Clk), .RN(n3897), .Q(
        \pc_lut[7][30] ), .QN(n1979) );
  DFFR_X1 \pc_lut_reg[8][31]  ( .D(n7281), .CK(Clk), .RN(n3897), .QN(n1977) );
  DFFR_X1 \pc_lut_reg[8][29]  ( .D(n7280), .CK(Clk), .RN(n3897), .QN(n1976) );
  DFFR_X1 \pc_lut_reg[8][27]  ( .D(n7279), .CK(Clk), .RN(n3897), .QN(n1975) );
  DFFR_X1 \pc_lut_reg[8][25]  ( .D(n7278), .CK(Clk), .RN(n3897), .QN(n1974) );
  DFFR_X1 \pc_lut_reg[8][23]  ( .D(n7277), .CK(Clk), .RN(n3898), .QN(n1973) );
  DFFR_X1 \pc_lut_reg[8][21]  ( .D(n7276), .CK(Clk), .RN(n3898), .QN(n1972) );
  DFFR_X1 \pc_lut_reg[8][19]  ( .D(n7275), .CK(Clk), .RN(n3898), .QN(n1971) );
  DFFR_X1 \pc_lut_reg[8][17]  ( .D(n7274), .CK(Clk), .RN(n3898), .QN(n1970) );
  DFFR_X1 \pc_lut_reg[8][15]  ( .D(n7273), .CK(Clk), .RN(n3898), .QN(n1969) );
  DFFR_X1 \pc_lut_reg[8][13]  ( .D(n7272), .CK(Clk), .RN(n3898), .QN(n1968) );
  DFFR_X1 \pc_lut_reg[8][11]  ( .D(n7271), .CK(Clk), .RN(n3898), .QN(n1967) );
  DFFR_X1 \pc_lut_reg[8][9]  ( .D(n7270), .CK(Clk), .RN(n3898), .QN(n1966) );
  DFFR_X1 \pc_lut_reg[8][7]  ( .D(n7269), .CK(Clk), .RN(n3898), .QN(n1965) );
  DFFR_X1 \pc_lut_reg[8][5]  ( .D(n7268), .CK(Clk), .RN(n3859), .QN(n1964) );
  DFFR_X1 \pc_lut_reg[8][3]  ( .D(n7267), .CK(Clk), .RN(n3898), .QN(n1963) );
  DFFR_X1 \pc_lut_reg[8][6]  ( .D(n7262), .CK(Clk), .RN(n3898), .QN(n1958) );
  DFFR_X1 \pc_lut_reg[8][8]  ( .D(n7261), .CK(Clk), .RN(n3898), .QN(n1957) );
  DFFR_X1 \pc_lut_reg[8][10]  ( .D(n7260), .CK(Clk), .RN(n3898), .QN(n1956) );
  DFFR_X1 \pc_lut_reg[8][12]  ( .D(n7259), .CK(Clk), .RN(n3898), .QN(n1955) );
  DFFR_X1 \pc_lut_reg[8][14]  ( .D(n7258), .CK(Clk), .RN(n3899), .QN(n1954) );
  DFFR_X1 \pc_lut_reg[8][16]  ( .D(n7257), .CK(Clk), .RN(n3899), .QN(n1953) );
  DFFR_X1 \pc_lut_reg[8][18]  ( .D(n7256), .CK(Clk), .RN(n3862), .QN(n1952) );
  DFFR_X1 \pc_lut_reg[8][20]  ( .D(n7255), .CK(Clk), .RN(n3899), .QN(n1951) );
  DFFR_X1 \pc_lut_reg[8][22]  ( .D(n7254), .CK(Clk), .RN(n3899), .QN(n1950) );
  DFFR_X1 \pc_lut_reg[8][24]  ( .D(n7253), .CK(Clk), .RN(n3899), .QN(n1949) );
  DFFR_X1 \pc_lut_reg[8][26]  ( .D(n7252), .CK(Clk), .RN(n3899), .QN(n1948) );
  DFFR_X1 \pc_lut_reg[8][28]  ( .D(n7251), .CK(Clk), .RN(n3899), .QN(n1947) );
  DFFR_X1 \pc_lut_reg[8][30]  ( .D(n7250), .CK(Clk), .RN(n3899), .QN(n1945) );
  DFFR_X1 \pc_lut_reg[9][31]  ( .D(n7249), .CK(Clk), .RN(n3898), .QN(n1943) );
  DFFR_X1 \pc_lut_reg[9][29]  ( .D(n7248), .CK(Clk), .RN(n3899), .QN(n1942) );
  DFFR_X1 \pc_lut_reg[9][27]  ( .D(n7247), .CK(Clk), .RN(n3899), .QN(n1941) );
  DFFR_X1 \pc_lut_reg[9][25]  ( .D(n7246), .CK(Clk), .RN(n3899), .QN(n1940) );
  DFFR_X1 \pc_lut_reg[9][23]  ( .D(n7245), .CK(Clk), .RN(n3899), .QN(n1939) );
  DFFR_X1 \pc_lut_reg[9][21]  ( .D(n7244), .CK(Clk), .RN(n3899), .QN(n1938) );
  DFFR_X1 \pc_lut_reg[9][19]  ( .D(n7243), .CK(Clk), .RN(n3899), .QN(n1937) );
  DFFR_X1 \pc_lut_reg[9][17]  ( .D(n7242), .CK(Clk), .RN(n3899), .QN(n1936) );
  DFFR_X1 \pc_lut_reg[9][15]  ( .D(n7241), .CK(Clk), .RN(n3900), .QN(n1935) );
  DFFR_X1 \pc_lut_reg[9][13]  ( .D(n7240), .CK(Clk), .RN(n3900), .QN(n1934) );
  DFFR_X1 \pc_lut_reg[9][11]  ( .D(n7239), .CK(Clk), .RN(n3900), .QN(n1933) );
  DFFR_X1 \pc_lut_reg[9][9]  ( .D(n7238), .CK(Clk), .RN(n3900), .QN(n1932) );
  DFFR_X1 \pc_lut_reg[9][7]  ( .D(n7237), .CK(Clk), .RN(n3900), .QN(n1931) );
  DFFR_X1 \pc_lut_reg[9][5]  ( .D(n7236), .CK(Clk), .RN(n3859), .QN(n1930) );
  DFFR_X1 \pc_lut_reg[9][3]  ( .D(n7235), .CK(Clk), .RN(n3900), .QN(n1929) );
  DFFR_X1 \pc_lut_reg[9][0]  ( .D(n7233), .CK(Clk), .RN(n3900), .QN(n1927) );
  DFFR_X1 \pc_lut_reg[9][6]  ( .D(n7230), .CK(Clk), .RN(n3900), .QN(n1924) );
  DFFR_X1 \pc_lut_reg[9][8]  ( .D(n7229), .CK(Clk), .RN(n3900), .QN(n1923) );
  DFFR_X1 \pc_lut_reg[9][10]  ( .D(n7228), .CK(Clk), .RN(n3900), .QN(n1922) );
  DFFR_X1 \pc_lut_reg[9][12]  ( .D(n7227), .CK(Clk), .RN(n3900), .QN(n1921) );
  DFFR_X1 \pc_lut_reg[9][14]  ( .D(n7226), .CK(Clk), .RN(n3900), .QN(n1920) );
  DFFR_X1 \pc_lut_reg[9][16]  ( .D(n7225), .CK(Clk), .RN(n3900), .QN(n1919) );
  DFFR_X1 \pc_lut_reg[9][18]  ( .D(n7224), .CK(Clk), .RN(n3862), .QN(n1918) );
  DFFR_X1 \pc_lut_reg[9][20]  ( .D(n7223), .CK(Clk), .RN(n3900), .QN(n1917) );
  DFFR_X1 \pc_lut_reg[9][22]  ( .D(n7222), .CK(Clk), .RN(n3901), .QN(n1916) );
  DFFR_X1 \pc_lut_reg[9][24]  ( .D(n7221), .CK(Clk), .RN(n3901), .QN(n1915) );
  DFFR_X1 \pc_lut_reg[9][26]  ( .D(n7220), .CK(Clk), .RN(n3901), .QN(n1914) );
  DFFR_X1 \pc_lut_reg[9][28]  ( .D(n7219), .CK(Clk), .RN(n3901), .QN(n1913) );
  DFFR_X1 \pc_lut_reg[9][30]  ( .D(n7218), .CK(Clk), .RN(n3901), .QN(n1911) );
  DFFR_X1 \pc_lut_reg[10][31]  ( .D(n7217), .CK(Clk), .RN(n3901), .Q(
        \pc_lut[10][31] ), .QN(n1909) );
  DFFR_X1 \pc_lut_reg[10][29]  ( .D(n7216), .CK(Clk), .RN(n3901), .Q(
        \pc_lut[10][29] ), .QN(n1908) );
  DFFR_X1 \pc_lut_reg[10][27]  ( .D(n7215), .CK(Clk), .RN(n3901), .Q(
        \pc_lut[10][27] ), .QN(n1907) );
  DFFR_X1 \pc_lut_reg[10][25]  ( .D(n7214), .CK(Clk), .RN(n3901), .Q(
        \pc_lut[10][25] ), .QN(n1906) );
  DFFR_X1 \pc_lut_reg[10][23]  ( .D(n7213), .CK(Clk), .RN(n3901), .Q(
        \pc_lut[10][23] ), .QN(n1905) );
  DFFR_X1 \pc_lut_reg[10][21]  ( .D(n7212), .CK(Clk), .RN(n3901), .Q(
        \pc_lut[10][21] ), .QN(n1904) );
  DFFR_X1 \pc_lut_reg[10][19]  ( .D(n7211), .CK(Clk), .RN(n3901), .Q(
        \pc_lut[10][19] ), .QN(n1903) );
  DFFR_X1 \pc_lut_reg[10][17]  ( .D(n7210), .CK(Clk), .RN(n3901), .Q(
        \pc_lut[10][17] ), .QN(n1902) );
  DFFR_X1 \pc_lut_reg[10][15]  ( .D(n7209), .CK(Clk), .RN(n3901), .Q(
        \pc_lut[10][15] ), .QN(n1901) );
  DFFR_X1 \pc_lut_reg[10][13]  ( .D(n7208), .CK(Clk), .RN(n3901), .Q(
        \pc_lut[10][13] ), .QN(n1900) );
  DFFR_X1 \pc_lut_reg[10][11]  ( .D(n7207), .CK(Clk), .RN(n3902), .Q(
        \pc_lut[10][11] ), .QN(n1899) );
  DFFR_X1 \pc_lut_reg[10][9]  ( .D(n7206), .CK(Clk), .RN(n3902), .Q(
        \pc_lut[10][9] ), .QN(n1898) );
  DFFR_X1 \pc_lut_reg[10][7]  ( .D(n7205), .CK(Clk), .RN(n3902), .Q(
        \pc_lut[10][7] ), .QN(n1897) );
  DFFR_X1 \pc_lut_reg[10][5]  ( .D(n7204), .CK(Clk), .RN(n3859), .Q(
        \pc_lut[10][5] ), .QN(n1896) );
  DFFR_X1 \pc_lut_reg[10][3]  ( .D(n7203), .CK(Clk), .RN(n3902), .Q(
        \pc_lut[10][3] ) );
  DFFR_X1 \pc_lut_reg[10][1]  ( .D(n7202), .CK(Clk), .RN(n3902), .Q(
        \pc_lut[10][1] ) );
  DFFR_X1 \pc_lut_reg[10][6]  ( .D(n7198), .CK(Clk), .RN(n3902), .Q(
        \pc_lut[10][6] ), .QN(n1893) );
  DFFR_X1 \pc_lut_reg[10][8]  ( .D(n7197), .CK(Clk), .RN(n3902), .Q(
        \pc_lut[10][8] ), .QN(n1892) );
  DFFR_X1 \pc_lut_reg[10][10]  ( .D(n7196), .CK(Clk), .RN(n3902), .Q(
        \pc_lut[10][10] ), .QN(n1891) );
  DFFR_X1 \pc_lut_reg[10][12]  ( .D(n7195), .CK(Clk), .RN(n3902), .Q(
        \pc_lut[10][12] ), .QN(n1890) );
  DFFR_X1 \pc_lut_reg[10][14]  ( .D(n7194), .CK(Clk), .RN(n3902), .Q(
        \pc_lut[10][14] ), .QN(n1889) );
  DFFR_X1 \pc_lut_reg[10][16]  ( .D(n7193), .CK(Clk), .RN(n3902), .Q(
        \pc_lut[10][16] ), .QN(n1888) );
  DFFR_X1 \pc_lut_reg[10][18]  ( .D(n7192), .CK(Clk), .RN(n3862), .Q(
        \pc_lut[10][18] ), .QN(n1887) );
  DFFR_X1 \pc_lut_reg[10][20]  ( .D(n7191), .CK(Clk), .RN(n3902), .Q(
        \pc_lut[10][20] ), .QN(n1886) );
  DFFR_X1 \pc_lut_reg[10][22]  ( .D(n7190), .CK(Clk), .RN(n3902), .Q(
        \pc_lut[10][22] ), .QN(n1885) );
  DFFR_X1 \pc_lut_reg[10][24]  ( .D(n7189), .CK(Clk), .RN(n3902), .Q(
        \pc_lut[10][24] ), .QN(n1884) );
  DFFR_X1 \pc_lut_reg[10][26]  ( .D(n7188), .CK(Clk), .RN(n3902), .Q(
        \pc_lut[10][26] ), .QN(n1883) );
  DFFR_X1 \pc_lut_reg[10][28]  ( .D(n7187), .CK(Clk), .RN(n3903), .Q(
        \pc_lut[10][28] ), .QN(n1882) );
  DFFR_X1 \pc_lut_reg[10][30]  ( .D(n7186), .CK(Clk), .RN(n3903), .Q(
        \pc_lut[10][30] ), .QN(n1880) );
  DFFR_X1 \pc_lut_reg[11][31]  ( .D(n7185), .CK(Clk), .RN(n3903), .Q(
        \pc_lut[11][31] ), .QN(n1877) );
  DFFR_X1 \pc_lut_reg[11][29]  ( .D(n7184), .CK(Clk), .RN(n3903), .Q(
        \pc_lut[11][29] ), .QN(n1876) );
  DFFR_X1 \pc_lut_reg[11][27]  ( .D(n7183), .CK(Clk), .RN(n3903), .Q(
        \pc_lut[11][27] ), .QN(n1875) );
  DFFR_X1 \pc_lut_reg[11][25]  ( .D(n7182), .CK(Clk), .RN(n3903), .Q(
        \pc_lut[11][25] ), .QN(n1874) );
  DFFR_X1 \pc_lut_reg[11][23]  ( .D(n7181), .CK(Clk), .RN(n3903), .Q(
        \pc_lut[11][23] ), .QN(n1873) );
  DFFR_X1 \pc_lut_reg[11][21]  ( .D(n7180), .CK(Clk), .RN(n3903), .Q(
        \pc_lut[11][21] ), .QN(n1872) );
  DFFR_X1 \pc_lut_reg[11][19]  ( .D(n7179), .CK(Clk), .RN(n3903), .Q(
        \pc_lut[11][19] ), .QN(n1871) );
  DFFR_X1 \pc_lut_reg[11][17]  ( .D(n7178), .CK(Clk), .RN(n3903), .Q(
        \pc_lut[11][17] ), .QN(n1870) );
  DFFR_X1 \pc_lut_reg[11][15]  ( .D(n7177), .CK(Clk), .RN(n3903), .Q(
        \pc_lut[11][15] ), .QN(n1869) );
  DFFR_X1 \pc_lut_reg[11][13]  ( .D(n7176), .CK(Clk), .RN(n3903), .Q(
        \pc_lut[11][13] ), .QN(n1868) );
  DFFR_X1 \pc_lut_reg[11][11]  ( .D(n7175), .CK(Clk), .RN(n3903), .Q(
        \pc_lut[11][11] ), .QN(n1867) );
  DFFR_X1 \pc_lut_reg[11][9]  ( .D(n7174), .CK(Clk), .RN(n3903), .Q(
        \pc_lut[11][9] ), .QN(n1866) );
  DFFR_X1 \pc_lut_reg[11][7]  ( .D(n7173), .CK(Clk), .RN(n3903), .Q(
        \pc_lut[11][7] ), .QN(n1865) );
  DFFR_X1 \pc_lut_reg[11][5]  ( .D(n7172), .CK(Clk), .RN(n3859), .Q(
        \pc_lut[11][5] ), .QN(n1864) );
  DFFR_X1 \pc_lut_reg[11][3]  ( .D(n7171), .CK(Clk), .RN(n3904), .Q(
        \pc_lut[11][3] ) );
  DFFR_X1 \pc_lut_reg[11][1]  ( .D(n7170), .CK(Clk), .RN(n3904), .Q(
        \pc_lut[11][1] ) );
  DFFR_X1 \pc_lut_reg[11][0]  ( .D(n7169), .CK(Clk), .RN(n3904), .Q(
        \pc_lut[11][0] ) );
  DFFR_X1 \pc_lut_reg[11][6]  ( .D(n7166), .CK(Clk), .RN(n3904), .Q(
        \pc_lut[11][6] ), .QN(n1860) );
  DFFR_X1 \pc_lut_reg[11][8]  ( .D(n7165), .CK(Clk), .RN(n3904), .Q(
        \pc_lut[11][8] ), .QN(n1859) );
  DFFR_X1 \pc_lut_reg[11][10]  ( .D(n7164), .CK(Clk), .RN(n3904), .Q(
        \pc_lut[11][10] ), .QN(n1858) );
  DFFR_X1 \pc_lut_reg[11][12]  ( .D(n7163), .CK(Clk), .RN(n3904), .Q(
        \pc_lut[11][12] ), .QN(n1857) );
  DFFR_X1 \pc_lut_reg[11][14]  ( .D(n7162), .CK(Clk), .RN(n3904), .Q(
        \pc_lut[11][14] ), .QN(n1856) );
  DFFR_X1 \pc_lut_reg[11][16]  ( .D(n7161), .CK(Clk), .RN(n3904), .Q(
        \pc_lut[11][16] ), .QN(n1855) );
  DFFR_X1 \pc_lut_reg[11][18]  ( .D(n7160), .CK(Clk), .RN(n3862), .Q(
        \pc_lut[11][18] ), .QN(n1854) );
  DFFR_X1 \pc_lut_reg[11][20]  ( .D(n7159), .CK(Clk), .RN(n3892), .Q(
        \pc_lut[11][20] ), .QN(n1853) );
  DFFR_X1 \pc_lut_reg[11][22]  ( .D(n7158), .CK(Clk), .RN(n3888), .Q(
        \pc_lut[11][22] ), .QN(n1852) );
  DFFR_X1 \pc_lut_reg[11][24]  ( .D(n7157), .CK(Clk), .RN(n3888), .Q(
        \pc_lut[11][24] ), .QN(n1851) );
  DFFR_X1 \pc_lut_reg[11][26]  ( .D(n7156), .CK(Clk), .RN(n3888), .Q(
        \pc_lut[11][26] ), .QN(n1850) );
  DFFR_X1 \pc_lut_reg[11][28]  ( .D(n7155), .CK(Clk), .RN(n3888), .Q(
        \pc_lut[11][28] ), .QN(n1849) );
  DFFR_X1 \pc_lut_reg[11][30]  ( .D(n7154), .CK(Clk), .RN(n3888), .Q(
        \pc_lut[11][30] ), .QN(n1847) );
  DFFR_X1 \pc_lut_reg[12][31]  ( .D(n7153), .CK(Clk), .RN(n3888), .QN(n1842)
         );
  DFFR_X1 \pc_lut_reg[12][29]  ( .D(n7152), .CK(Clk), .RN(n3888), .QN(n1841)
         );
  DFFR_X1 \pc_lut_reg[12][27]  ( .D(n7151), .CK(Clk), .RN(n3888), .QN(n1840)
         );
  DFFR_X1 \pc_lut_reg[12][25]  ( .D(n7150), .CK(Clk), .RN(n3888), .QN(n1839)
         );
  DFFR_X1 \pc_lut_reg[12][23]  ( .D(n7149), .CK(Clk), .RN(n3888), .QN(n1838)
         );
  DFFR_X1 \pc_lut_reg[12][21]  ( .D(n7148), .CK(Clk), .RN(n3888), .QN(n1837)
         );
  DFFR_X1 \pc_lut_reg[12][19]  ( .D(n7147), .CK(Clk), .RN(n3889), .QN(n1836)
         );
  DFFR_X1 \pc_lut_reg[12][17]  ( .D(n7146), .CK(Clk), .RN(n3889), .QN(n1835)
         );
  DFFR_X1 \pc_lut_reg[12][15]  ( .D(n7145), .CK(Clk), .RN(n3889), .QN(n1834)
         );
  DFFR_X1 \pc_lut_reg[12][13]  ( .D(n7144), .CK(Clk), .RN(n3889), .QN(n1833)
         );
  DFFR_X1 \pc_lut_reg[12][11]  ( .D(n7143), .CK(Clk), .RN(n3889), .QN(n1832)
         );
  DFFR_X1 \pc_lut_reg[12][9]  ( .D(n7142), .CK(Clk), .RN(n3889), .QN(n1831) );
  DFFR_X1 \pc_lut_reg[12][7]  ( .D(n7141), .CK(Clk), .RN(n3889), .QN(n1830) );
  DFFR_X1 \pc_lut_reg[12][5]  ( .D(n7140), .CK(Clk), .RN(n3859), .QN(n1829) );
  DFFR_X1 \pc_lut_reg[12][3]  ( .D(n7139), .CK(Clk), .RN(n3889), .QN(n1828) );
  DFFR_X1 \pc_lut_reg[12][2]  ( .D(n7136), .CK(Clk), .RN(n3889), .QN(n1825) );
  DFFR_X1 \pc_lut_reg[12][6]  ( .D(n7134), .CK(Clk), .RN(n3889), .QN(n1823) );
  DFFR_X1 \pc_lut_reg[12][8]  ( .D(n7133), .CK(Clk), .RN(n3889), .QN(n1822) );
  DFFR_X1 \pc_lut_reg[12][10]  ( .D(n7132), .CK(Clk), .RN(n3889), .QN(n1821)
         );
  DFFR_X1 \pc_lut_reg[12][12]  ( .D(n7131), .CK(Clk), .RN(n3889), .QN(n1820)
         );
  DFFR_X1 \pc_lut_reg[12][14]  ( .D(n7130), .CK(Clk), .RN(n3889), .QN(n1819)
         );
  DFFR_X1 \pc_lut_reg[12][16]  ( .D(n7129), .CK(Clk), .RN(n3889), .QN(n1818)
         );
  DFFR_X1 \pc_lut_reg[12][18]  ( .D(n7128), .CK(Clk), .RN(n3862), .QN(n1817)
         );
  DFFR_X1 \pc_lut_reg[12][20]  ( .D(n7127), .CK(Clk), .RN(n3890), .QN(n1816)
         );
  DFFR_X1 \pc_lut_reg[12][22]  ( .D(n7126), .CK(Clk), .RN(n3890), .QN(n1815)
         );
  DFFR_X1 \pc_lut_reg[12][24]  ( .D(n7125), .CK(Clk), .RN(n3890), .QN(n1814)
         );
  DFFR_X1 \pc_lut_reg[12][26]  ( .D(n7124), .CK(Clk), .RN(n3890), .QN(n1813)
         );
  DFFR_X1 \pc_lut_reg[12][28]  ( .D(n7123), .CK(Clk), .RN(n3890), .QN(n1812)
         );
  DFFR_X1 \pc_lut_reg[12][30]  ( .D(n7122), .CK(Clk), .RN(n3890), .QN(n1810)
         );
  DFFR_X1 \pc_lut_reg[13][31]  ( .D(n7121), .CK(Clk), .RN(n3890), .QN(n1808)
         );
  DFFR_X1 \pc_lut_reg[13][29]  ( .D(n7120), .CK(Clk), .RN(n3890), .QN(n1807)
         );
  DFFR_X1 \pc_lut_reg[13][27]  ( .D(n7119), .CK(Clk), .RN(n3890), .QN(n1806)
         );
  DFFR_X1 \pc_lut_reg[13][25]  ( .D(n7118), .CK(Clk), .RN(n3890), .QN(n1805)
         );
  DFFR_X1 \pc_lut_reg[13][23]  ( .D(n7117), .CK(Clk), .RN(n3890), .QN(n1804)
         );
  DFFR_X1 \pc_lut_reg[13][21]  ( .D(n7116), .CK(Clk), .RN(n3890), .QN(n1803)
         );
  DFFR_X1 \pc_lut_reg[13][19]  ( .D(n7115), .CK(Clk), .RN(n3890), .QN(n1802)
         );
  DFFR_X1 \pc_lut_reg[13][17]  ( .D(n7114), .CK(Clk), .RN(n3890), .QN(n1801)
         );
  DFFR_X1 \pc_lut_reg[13][15]  ( .D(n7113), .CK(Clk), .RN(n3890), .QN(n1800)
         );
  DFFR_X1 \pc_lut_reg[13][13]  ( .D(n7112), .CK(Clk), .RN(n3891), .QN(n1799)
         );
  DFFR_X1 \pc_lut_reg[13][11]  ( .D(n7111), .CK(Clk), .RN(n3891), .QN(n1798)
         );
  DFFR_X1 \pc_lut_reg[13][9]  ( .D(n7110), .CK(Clk), .RN(n3891), .QN(n1797) );
  DFFR_X1 \pc_lut_reg[13][7]  ( .D(n7109), .CK(Clk), .RN(n3891), .QN(n1796) );
  DFFR_X1 \pc_lut_reg[13][5]  ( .D(n7108), .CK(Clk), .RN(n3859), .QN(n1795) );
  DFFR_X1 \pc_lut_reg[13][3]  ( .D(n7107), .CK(Clk), .RN(n3891), .QN(n1794) );
  DFFR_X1 \pc_lut_reg[13][0]  ( .D(n7105), .CK(Clk), .RN(n3891), .QN(n1792) );
  DFFR_X1 \pc_lut_reg[13][2]  ( .D(n7104), .CK(Clk), .RN(n3891), .QN(n1791) );
  DFFR_X1 \pc_lut_reg[13][6]  ( .D(n7102), .CK(Clk), .RN(n3891), .QN(n1789) );
  DFFR_X1 \pc_lut_reg[13][8]  ( .D(n7101), .CK(Clk), .RN(n3891), .QN(n1788) );
  DFFR_X1 \pc_lut_reg[13][10]  ( .D(n7100), .CK(Clk), .RN(n3891), .QN(n1787)
         );
  DFFR_X1 \pc_lut_reg[13][12]  ( .D(n7099), .CK(Clk), .RN(n3891), .QN(n1786)
         );
  DFFR_X1 \pc_lut_reg[13][14]  ( .D(n7098), .CK(Clk), .RN(n3891), .QN(n1785)
         );
  DFFR_X1 \pc_lut_reg[13][16]  ( .D(n7097), .CK(Clk), .RN(n3891), .QN(n1784)
         );
  DFFR_X1 \pc_lut_reg[13][18]  ( .D(n7096), .CK(Clk), .RN(n3862), .QN(n1783)
         );
  DFFR_X1 \pc_lut_reg[13][20]  ( .D(n7095), .CK(Clk), .RN(n3891), .QN(n1782)
         );
  DFFR_X1 \pc_lut_reg[13][22]  ( .D(n7094), .CK(Clk), .RN(n3891), .QN(n1781)
         );
  DFFR_X1 \pc_lut_reg[13][24]  ( .D(n7093), .CK(Clk), .RN(n3892), .QN(n1780)
         );
  DFFR_X1 \pc_lut_reg[13][26]  ( .D(n7092), .CK(Clk), .RN(n3892), .QN(n1779)
         );
  DFFR_X1 \pc_lut_reg[13][28]  ( .D(n7091), .CK(Clk), .RN(n3892), .QN(n1778)
         );
  DFFR_X1 \pc_lut_reg[13][30]  ( .D(n7090), .CK(Clk), .RN(n3892), .QN(n1776)
         );
  DFFR_X1 \pc_lut_reg[14][31]  ( .D(n7089), .CK(Clk), .RN(n3892), .Q(
        \pc_lut[14][31] ), .QN(n1774) );
  DFFR_X1 \pc_lut_reg[14][29]  ( .D(n7088), .CK(Clk), .RN(n3892), .Q(
        \pc_lut[14][29] ), .QN(n1773) );
  DFFR_X1 \pc_lut_reg[14][27]  ( .D(n7087), .CK(Clk), .RN(n3892), .Q(
        \pc_lut[14][27] ), .QN(n1772) );
  DFFR_X1 \pc_lut_reg[14][25]  ( .D(n7086), .CK(Clk), .RN(n3892), .Q(
        \pc_lut[14][25] ), .QN(n1771) );
  DFFR_X1 \pc_lut_reg[14][23]  ( .D(n7085), .CK(Clk), .RN(n3892), .Q(
        \pc_lut[14][23] ), .QN(n1770) );
  DFFR_X1 \pc_lut_reg[14][21]  ( .D(n7084), .CK(Clk), .RN(n3892), .Q(
        \pc_lut[14][21] ), .QN(n1769) );
  DFFR_X1 \pc_lut_reg[14][19]  ( .D(n7083), .CK(Clk), .RN(n3892), .Q(
        \pc_lut[14][19] ), .QN(n1768) );
  DFFR_X1 \pc_lut_reg[14][17]  ( .D(n7082), .CK(Clk), .RN(n3892), .Q(
        \pc_lut[14][17] ), .QN(n1767) );
  DFFR_X1 \pc_lut_reg[14][15]  ( .D(n7081), .CK(Clk), .RN(n3892), .Q(
        \pc_lut[14][15] ), .QN(n1766) );
  DFFR_X1 \pc_lut_reg[14][13]  ( .D(n7080), .CK(Clk), .RN(n3892), .Q(
        \pc_lut[14][13] ), .QN(n1765) );
  DFFR_X1 \pc_lut_reg[14][11]  ( .D(n7079), .CK(Clk), .RN(n3893), .Q(
        \pc_lut[14][11] ), .QN(n1764) );
  DFFR_X1 \pc_lut_reg[14][9]  ( .D(n7078), .CK(Clk), .RN(n3893), .Q(
        \pc_lut[14][9] ), .QN(n1763) );
  DFFR_X1 \pc_lut_reg[14][7]  ( .D(n7077), .CK(Clk), .RN(n3893), .Q(
        \pc_lut[14][7] ), .QN(n1762) );
  DFFR_X1 \pc_lut_reg[14][5]  ( .D(n7076), .CK(Clk), .RN(n3859), .Q(
        \pc_lut[14][5] ), .QN(n1761) );
  DFFR_X1 \pc_lut_reg[14][6]  ( .D(n7070), .CK(Clk), .RN(n3893), .Q(
        \pc_lut[14][6] ), .QN(n1757) );
  DFFR_X1 \pc_lut_reg[14][8]  ( .D(n7069), .CK(Clk), .RN(n3893), .Q(
        \pc_lut[14][8] ), .QN(n1756) );
  DFFR_X1 \pc_lut_reg[14][10]  ( .D(n7068), .CK(Clk), .RN(n3893), .Q(
        \pc_lut[14][10] ), .QN(n1755) );
  DFFR_X1 \pc_lut_reg[14][12]  ( .D(n7067), .CK(Clk), .RN(n3893), .Q(
        \pc_lut[14][12] ), .QN(n1754) );
  DFFR_X1 \pc_lut_reg[14][14]  ( .D(n7066), .CK(Clk), .RN(n3893), .Q(
        \pc_lut[14][14] ), .QN(n1753) );
  DFFR_X1 \pc_lut_reg[14][16]  ( .D(n7065), .CK(Clk), .RN(n3893), .Q(
        \pc_lut[14][16] ), .QN(n1752) );
  DFFR_X1 \pc_lut_reg[14][18]  ( .D(n7064), .CK(Clk), .RN(n3862), .Q(
        \pc_lut[14][18] ), .QN(n1751) );
  DFFR_X1 \pc_lut_reg[14][20]  ( .D(n7063), .CK(Clk), .RN(n3893), .Q(
        \pc_lut[14][20] ), .QN(n1750) );
  DFFR_X1 \pc_lut_reg[14][22]  ( .D(n7062), .CK(Clk), .RN(n3893), .Q(
        \pc_lut[14][22] ), .QN(n1749) );
  DFFR_X1 \pc_lut_reg[14][24]  ( .D(n7061), .CK(Clk), .RN(n3893), .Q(
        \pc_lut[14][24] ), .QN(n1748) );
  DFFR_X1 \pc_lut_reg[14][26]  ( .D(n7060), .CK(Clk), .RN(n3893), .Q(
        \pc_lut[14][26] ), .QN(n1747) );
  DFFR_X1 \pc_lut_reg[14][28]  ( .D(n7059), .CK(Clk), .RN(n3893), .Q(
        \pc_lut[14][28] ), .QN(n1746) );
  DFFR_X1 \pc_lut_reg[14][30]  ( .D(n7058), .CK(Clk), .RN(n3893), .Q(
        \pc_lut[14][30] ), .QN(n1744) );
  DFFR_X1 \pc_lut_reg[15][31]  ( .D(n7057), .CK(Clk), .RN(n3894), .Q(
        \pc_lut[15][31] ), .QN(n1741) );
  DFFR_X1 \pc_lut_reg[15][29]  ( .D(n7056), .CK(Clk), .RN(n3894), .Q(
        \pc_lut[15][29] ), .QN(n1740) );
  DFFR_X1 \pc_lut_reg[15][27]  ( .D(n7055), .CK(Clk), .RN(n3894), .Q(
        \pc_lut[15][27] ), .QN(n1739) );
  DFFR_X1 \pc_lut_reg[15][25]  ( .D(n7054), .CK(Clk), .RN(n3894), .Q(
        \pc_lut[15][25] ), .QN(n1738) );
  DFFR_X1 \pc_lut_reg[15][23]  ( .D(n7053), .CK(Clk), .RN(n3894), .Q(
        \pc_lut[15][23] ), .QN(n1737) );
  DFFR_X1 \pc_lut_reg[15][21]  ( .D(n7052), .CK(Clk), .RN(n3894), .Q(
        \pc_lut[15][21] ), .QN(n1736) );
  DFFR_X1 \pc_lut_reg[15][19]  ( .D(n7051), .CK(Clk), .RN(n3894), .Q(
        \pc_lut[15][19] ), .QN(n1735) );
  DFFR_X1 \pc_lut_reg[15][17]  ( .D(n7050), .CK(Clk), .RN(n3894), .Q(
        \pc_lut[15][17] ), .QN(n1734) );
  DFFR_X1 \pc_lut_reg[15][15]  ( .D(n7049), .CK(Clk), .RN(n3894), .Q(
        \pc_lut[15][15] ), .QN(n1733) );
  DFFR_X1 \pc_lut_reg[15][13]  ( .D(n7048), .CK(Clk), .RN(n3894), .Q(
        \pc_lut[15][13] ), .QN(n1732) );
  DFFR_X1 \pc_lut_reg[15][11]  ( .D(n7047), .CK(Clk), .RN(n3894), .Q(
        \pc_lut[15][11] ), .QN(n1731) );
  DFFR_X1 \pc_lut_reg[15][9]  ( .D(n7046), .CK(Clk), .RN(n3894), .Q(
        \pc_lut[15][9] ), .QN(n1730) );
  DFFR_X1 \pc_lut_reg[15][7]  ( .D(n7045), .CK(Clk), .RN(n3894), .Q(
        \pc_lut[15][7] ), .QN(n1729) );
  DFFR_X1 \pc_lut_reg[15][5]  ( .D(n7044), .CK(Clk), .RN(n3859), .Q(
        \pc_lut[15][5] ), .QN(n1728) );
  DFFR_X1 \pc_lut_reg[15][6]  ( .D(n7038), .CK(Clk), .RN(n3947), .Q(
        \pc_lut[15][6] ), .QN(n1723) );
  DFFR_X1 \pc_lut_reg[15][8]  ( .D(n7037), .CK(Clk), .RN(n3947), .Q(
        \pc_lut[15][8] ), .QN(n1722) );
  DFFR_X1 \pc_lut_reg[15][10]  ( .D(n7036), .CK(Clk), .RN(n3947), .Q(
        \pc_lut[15][10] ), .QN(n1721) );
  DFFR_X1 \pc_lut_reg[15][12]  ( .D(n7035), .CK(Clk), .RN(n3947), .Q(
        \pc_lut[15][12] ), .QN(n1720) );
  DFFR_X1 \pc_lut_reg[15][14]  ( .D(n7034), .CK(Clk), .RN(n3947), .Q(
        \pc_lut[15][14] ), .QN(n1719) );
  DFFR_X1 \pc_lut_reg[15][16]  ( .D(n7033), .CK(Clk), .RN(n3948), .Q(
        \pc_lut[15][16] ), .QN(n1718) );
  DFFR_X1 \pc_lut_reg[15][18]  ( .D(n7032), .CK(Clk), .RN(n3863), .Q(
        \pc_lut[15][18] ), .QN(n1717) );
  DFFR_X1 \pc_lut_reg[15][20]  ( .D(n7031), .CK(Clk), .RN(n3948), .Q(
        \pc_lut[15][20] ), .QN(n1716) );
  DFFR_X1 \pc_lut_reg[15][22]  ( .D(n7030), .CK(Clk), .RN(n3948), .Q(
        \pc_lut[15][22] ), .QN(n1715) );
  DFFR_X1 \pc_lut_reg[15][24]  ( .D(n7029), .CK(Clk), .RN(n3948), .Q(
        \pc_lut[15][24] ), .QN(n1714) );
  DFFR_X1 \pc_lut_reg[15][26]  ( .D(n7028), .CK(Clk), .RN(n3948), .Q(
        \pc_lut[15][26] ), .QN(n1713) );
  DFFR_X1 \pc_lut_reg[15][28]  ( .D(n7027), .CK(Clk), .RN(n3948), .Q(
        \pc_lut[15][28] ), .QN(n1712) );
  DFFR_X1 \pc_lut_reg[15][30]  ( .D(n7026), .CK(Clk), .RN(n3949), .Q(
        \pc_lut[15][30] ), .QN(n1710) );
  DFFR_X1 \pc_lut_reg[16][31]  ( .D(n7025), .CK(Clk), .RN(n3948), .QN(n1707)
         );
  DFFR_X1 \pc_lut_reg[16][29]  ( .D(n7024), .CK(Clk), .RN(n3948), .QN(n1706)
         );
  DFFR_X1 \pc_lut_reg[16][27]  ( .D(n7023), .CK(Clk), .RN(n3948), .QN(n1705)
         );
  DFFR_X1 \pc_lut_reg[16][25]  ( .D(n7022), .CK(Clk), .RN(n3948), .QN(n1704)
         );
  DFFR_X1 \pc_lut_reg[16][23]  ( .D(n7021), .CK(Clk), .RN(n3948), .QN(n1703)
         );
  DFFR_X1 \pc_lut_reg[16][21]  ( .D(n7020), .CK(Clk), .RN(n3948), .QN(n1702)
         );
  DFFR_X1 \pc_lut_reg[16][19]  ( .D(n7019), .CK(Clk), .RN(n3948), .QN(n1701)
         );
  DFFR_X1 \pc_lut_reg[16][17]  ( .D(n7018), .CK(Clk), .RN(n3948), .QN(n1700)
         );
  DFFR_X1 \pc_lut_reg[16][15]  ( .D(n7017), .CK(Clk), .RN(n3948), .QN(n1699)
         );
  DFFR_X1 \pc_lut_reg[16][13]  ( .D(n7016), .CK(Clk), .RN(n3949), .QN(n1698)
         );
  DFFR_X1 \pc_lut_reg[16][11]  ( .D(n7015), .CK(Clk), .RN(n3949), .QN(n1697)
         );
  DFFR_X1 \pc_lut_reg[16][9]  ( .D(n7014), .CK(Clk), .RN(n3949), .QN(n1696) );
  DFFR_X1 \pc_lut_reg[16][7]  ( .D(n7013), .CK(Clk), .RN(n3949), .QN(n1695) );
  DFFR_X1 \pc_lut_reg[16][5]  ( .D(n7012), .CK(Clk), .RN(n3859), .QN(n1694) );
  DFFR_X1 \pc_lut_reg[16][4]  ( .D(n7007), .CK(Clk), .RN(n3949), .QN(n1689) );
  DFFR_X1 \pc_lut_reg[16][6]  ( .D(n7006), .CK(Clk), .RN(n3949), .QN(n1688) );
  DFFR_X1 \pc_lut_reg[16][8]  ( .D(n7005), .CK(Clk), .RN(n3949), .QN(n1687) );
  DFFR_X1 \pc_lut_reg[16][10]  ( .D(n7004), .CK(Clk), .RN(n3949), .QN(n1686)
         );
  DFFR_X1 \pc_lut_reg[16][12]  ( .D(n7003), .CK(Clk), .RN(n3949), .QN(n1685)
         );
  DFFR_X1 \pc_lut_reg[16][14]  ( .D(n7002), .CK(Clk), .RN(n3949), .QN(n1684)
         );
  DFFR_X1 \pc_lut_reg[16][16]  ( .D(n7001), .CK(Clk), .RN(n3949), .QN(n1683)
         );
  DFFR_X1 \pc_lut_reg[16][18]  ( .D(n7000), .CK(Clk), .RN(n3862), .QN(n1682)
         );
  DFFR_X1 \pc_lut_reg[16][20]  ( .D(n6999), .CK(Clk), .RN(n3949), .QN(n1681)
         );
  DFFR_X1 \pc_lut_reg[16][22]  ( .D(n6998), .CK(Clk), .RN(n3950), .QN(n1680)
         );
  DFFR_X1 \pc_lut_reg[16][24]  ( .D(n6997), .CK(Clk), .RN(n3950), .QN(n1679)
         );
  DFFR_X1 \pc_lut_reg[16][26]  ( .D(n6996), .CK(Clk), .RN(n3950), .QN(n1678)
         );
  DFFR_X1 \pc_lut_reg[16][28]  ( .D(n6995), .CK(Clk), .RN(n3950), .QN(n1677)
         );
  DFFR_X1 \pc_lut_reg[16][30]  ( .D(n6994), .CK(Clk), .RN(n3950), .QN(n1675)
         );
  DFFR_X1 \pc_lut_reg[17][31]  ( .D(n6993), .CK(Clk), .RN(n3950), .QN(n1673)
         );
  DFFR_X1 \pc_lut_reg[17][29]  ( .D(n6992), .CK(Clk), .RN(n3950), .QN(n1672)
         );
  DFFR_X1 \pc_lut_reg[17][27]  ( .D(n6991), .CK(Clk), .RN(n3950), .QN(n1671)
         );
  DFFR_X1 \pc_lut_reg[17][25]  ( .D(n6990), .CK(Clk), .RN(n3950), .QN(n1670)
         );
  DFFR_X1 \pc_lut_reg[17][23]  ( .D(n6989), .CK(Clk), .RN(n3950), .QN(n1669)
         );
  DFFR_X1 \pc_lut_reg[17][21]  ( .D(n6988), .CK(Clk), .RN(n3950), .QN(n1668)
         );
  DFFR_X1 \pc_lut_reg[17][19]  ( .D(n6987), .CK(Clk), .RN(n3950), .QN(n1667)
         );
  DFFR_X1 \pc_lut_reg[17][17]  ( .D(n6986), .CK(Clk), .RN(n3950), .QN(n1666)
         );
  DFFR_X1 \pc_lut_reg[17][15]  ( .D(n6985), .CK(Clk), .RN(n3950), .QN(n1665)
         );
  DFFR_X1 \pc_lut_reg[17][13]  ( .D(n6984), .CK(Clk), .RN(n3951), .QN(n1664)
         );
  DFFR_X1 \pc_lut_reg[17][11]  ( .D(n6983), .CK(Clk), .RN(n3951), .QN(n1663)
         );
  DFFR_X1 \pc_lut_reg[17][9]  ( .D(n6982), .CK(Clk), .RN(n3951), .QN(n1662) );
  DFFR_X1 \pc_lut_reg[17][7]  ( .D(n6981), .CK(Clk), .RN(n3950), .QN(n1661) );
  DFFR_X1 \pc_lut_reg[17][5]  ( .D(n6980), .CK(Clk), .RN(n3859), .QN(n1660) );
  DFFR_X1 \pc_lut_reg[17][0]  ( .D(n6977), .CK(Clk), .RN(n3951), .QN(n1657) );
  DFFR_X1 \pc_lut_reg[17][4]  ( .D(n6975), .CK(Clk), .RN(n3951), .QN(n1655) );
  DFFR_X1 \pc_lut_reg[17][6]  ( .D(n6974), .CK(Clk), .RN(n3951), .QN(n1654) );
  DFFR_X1 \pc_lut_reg[17][8]  ( .D(n6973), .CK(Clk), .RN(n3951), .QN(n1653) );
  DFFR_X1 \pc_lut_reg[17][10]  ( .D(n6972), .CK(Clk), .RN(n3951), .QN(n1652)
         );
  DFFR_X1 \pc_lut_reg[17][12]  ( .D(n6971), .CK(Clk), .RN(n3951), .QN(n1651)
         );
  DFFR_X1 \pc_lut_reg[17][14]  ( .D(n6970), .CK(Clk), .RN(n3949), .QN(n1650)
         );
  DFFR_X1 \pc_lut_reg[17][16]  ( .D(n6969), .CK(Clk), .RN(n3951), .QN(n1649)
         );
  DFFR_X1 \pc_lut_reg[17][18]  ( .D(n6968), .CK(Clk), .RN(n3862), .QN(n1648)
         );
  DFFR_X1 \pc_lut_reg[17][20]  ( .D(n6967), .CK(Clk), .RN(n3952), .QN(n1647)
         );
  DFFR_X1 \pc_lut_reg[17][22]  ( .D(n6966), .CK(Clk), .RN(n3952), .QN(n1646)
         );
  DFFR_X1 \pc_lut_reg[17][24]  ( .D(n6965), .CK(Clk), .RN(n3951), .QN(n1645)
         );
  DFFR_X1 \pc_lut_reg[17][26]  ( .D(n6964), .CK(Clk), .RN(n3952), .QN(n1644)
         );
  DFFR_X1 \pc_lut_reg[17][28]  ( .D(n6963), .CK(Clk), .RN(n3951), .QN(n1643)
         );
  DFFR_X1 \pc_lut_reg[17][30]  ( .D(n6962), .CK(Clk), .RN(n3952), .QN(n1641)
         );
  DFFR_X1 \pc_lut_reg[18][31]  ( .D(n6961), .CK(Clk), .RN(n3951), .Q(
        \pc_lut[18][31] ), .QN(n1639) );
  DFFR_X1 \pc_lut_reg[18][29]  ( .D(n6960), .CK(Clk), .RN(n3951), .Q(
        \pc_lut[18][29] ), .QN(n1638) );
  DFFR_X1 \pc_lut_reg[18][27]  ( .D(n6959), .CK(Clk), .RN(n3952), .Q(
        \pc_lut[18][27] ), .QN(n1637) );
  DFFR_X1 \pc_lut_reg[18][25]  ( .D(n6958), .CK(Clk), .RN(n3952), .Q(
        \pc_lut[18][25] ), .QN(n1636) );
  DFFR_X1 \pc_lut_reg[18][23]  ( .D(n6957), .CK(Clk), .RN(n3952), .Q(
        \pc_lut[18][23] ), .QN(n1635) );
  DFFR_X1 \pc_lut_reg[18][21]  ( .D(n6956), .CK(Clk), .RN(n3952), .Q(
        \pc_lut[18][21] ), .QN(n1634) );
  DFFR_X1 \pc_lut_reg[18][19]  ( .D(n6955), .CK(Clk), .RN(n3953), .Q(
        \pc_lut[18][19] ), .QN(n1633) );
  DFFR_X1 \pc_lut_reg[18][17]  ( .D(n6954), .CK(Clk), .RN(n3952), .Q(
        \pc_lut[18][17] ), .QN(n1632) );
  DFFR_X1 \pc_lut_reg[18][15]  ( .D(n6953), .CK(Clk), .RN(n3953), .Q(
        \pc_lut[18][15] ), .QN(n1631) );
  DFFR_X1 \pc_lut_reg[18][13]  ( .D(n6952), .CK(Clk), .RN(n3952), .Q(
        \pc_lut[18][13] ), .QN(n1630) );
  DFFR_X1 \pc_lut_reg[18][11]  ( .D(n6951), .CK(Clk), .RN(n3953), .Q(
        \pc_lut[18][11] ), .QN(n1629) );
  DFFR_X1 \pc_lut_reg[18][9]  ( .D(n6950), .CK(Clk), .RN(n3952), .Q(
        \pc_lut[18][9] ), .QN(n1628) );
  DFFR_X1 \pc_lut_reg[18][7]  ( .D(n6949), .CK(Clk), .RN(n3951), .Q(
        \pc_lut[18][7] ), .QN(n1627) );
  DFFR_X1 \pc_lut_reg[18][5]  ( .D(n6948), .CK(Clk), .RN(n3860), .Q(
        \pc_lut[18][5] ), .QN(n1626) );
  DFFR_X1 \pc_lut_reg[18][1]  ( .D(n6946), .CK(Clk), .RN(n3952), .Q(
        \pc_lut[18][1] ) );
  DFFR_X1 \pc_lut_reg[18][4]  ( .D(n6943), .CK(Clk), .RN(n3952), .Q(
        \pc_lut[18][4] ) );
  DFFR_X1 \pc_lut_reg[18][6]  ( .D(n6942), .CK(Clk), .RN(n3952), .Q(
        \pc_lut[18][6] ), .QN(n1623) );
  DFFR_X1 \pc_lut_reg[18][8]  ( .D(n6941), .CK(Clk), .RN(n3952), .Q(
        \pc_lut[18][8] ), .QN(n1622) );
  DFFR_X1 \pc_lut_reg[18][10]  ( .D(n6940), .CK(Clk), .RN(n3941), .Q(
        \pc_lut[18][10] ), .QN(n1621) );
  DFFR_X1 \pc_lut_reg[18][12]  ( .D(n6939), .CK(Clk), .RN(n3937), .Q(
        \pc_lut[18][12] ), .QN(n1620) );
  DFFR_X1 \pc_lut_reg[18][14]  ( .D(n6938), .CK(Clk), .RN(n3937), .Q(
        \pc_lut[18][14] ), .QN(n1619) );
  DFFR_X1 \pc_lut_reg[18][16]  ( .D(n6937), .CK(Clk), .RN(n3937), .Q(
        \pc_lut[18][16] ), .QN(n1618) );
  DFFR_X1 \pc_lut_reg[18][18]  ( .D(n6936), .CK(Clk), .RN(n3862), .Q(
        \pc_lut[18][18] ), .QN(n1617) );
  DFFR_X1 \pc_lut_reg[18][20]  ( .D(n6935), .CK(Clk), .RN(n3937), .Q(
        \pc_lut[18][20] ), .QN(n1616) );
  DFFR_X1 \pc_lut_reg[18][22]  ( .D(n6934), .CK(Clk), .RN(n3937), .Q(
        \pc_lut[18][22] ), .QN(n1615) );
  DFFR_X1 \pc_lut_reg[18][24]  ( .D(n6933), .CK(Clk), .RN(n3937), .Q(
        \pc_lut[18][24] ), .QN(n1614) );
  DFFR_X1 \pc_lut_reg[18][26]  ( .D(n6932), .CK(Clk), .RN(n3938), .Q(
        \pc_lut[18][26] ), .QN(n1613) );
  DFFR_X1 \pc_lut_reg[18][28]  ( .D(n6931), .CK(Clk), .RN(n3937), .Q(
        \pc_lut[18][28] ), .QN(n1612) );
  DFFR_X1 \pc_lut_reg[18][30]  ( .D(n6930), .CK(Clk), .RN(n3938), .Q(
        \pc_lut[18][30] ), .QN(n1610) );
  DFFR_X1 \pc_lut_reg[19][31]  ( .D(n6929), .CK(Clk), .RN(n3937), .Q(
        \pc_lut[19][31] ), .QN(n1607) );
  DFFR_X1 \pc_lut_reg[19][29]  ( .D(n6928), .CK(Clk), .RN(n3937), .Q(
        \pc_lut[19][29] ), .QN(n1606) );
  DFFR_X1 \pc_lut_reg[19][27]  ( .D(n6927), .CK(Clk), .RN(n3937), .Q(
        \pc_lut[19][27] ), .QN(n1605) );
  DFFR_X1 \pc_lut_reg[19][25]  ( .D(n6926), .CK(Clk), .RN(n3938), .Q(
        \pc_lut[19][25] ), .QN(n1604) );
  DFFR_X1 \pc_lut_reg[19][23]  ( .D(n6925), .CK(Clk), .RN(n3938), .Q(
        \pc_lut[19][23] ), .QN(n1603) );
  DFFR_X1 \pc_lut_reg[19][21]  ( .D(n6924), .CK(Clk), .RN(n3938), .Q(
        \pc_lut[19][21] ), .QN(n1602) );
  DFFR_X1 \pc_lut_reg[19][19]  ( .D(n6923), .CK(Clk), .RN(n3938), .Q(
        \pc_lut[19][19] ), .QN(n1601) );
  DFFR_X1 \pc_lut_reg[19][17]  ( .D(n6922), .CK(Clk), .RN(n3938), .Q(
        \pc_lut[19][17] ), .QN(n1600) );
  DFFR_X1 \pc_lut_reg[19][15]  ( .D(n6921), .CK(Clk), .RN(n3938), .Q(
        \pc_lut[19][15] ), .QN(n1599) );
  DFFR_X1 \pc_lut_reg[19][13]  ( .D(n6920), .CK(Clk), .RN(n3938), .Q(
        \pc_lut[19][13] ), .QN(n1598) );
  DFFR_X1 \pc_lut_reg[19][11]  ( .D(n6919), .CK(Clk), .RN(n3938), .Q(
        \pc_lut[19][11] ), .QN(n1597) );
  DFFR_X1 \pc_lut_reg[19][9]  ( .D(n6918), .CK(Clk), .RN(n3938), .Q(
        \pc_lut[19][9] ), .QN(n1596) );
  DFFR_X1 \pc_lut_reg[19][7]  ( .D(n6917), .CK(Clk), .RN(n3938), .Q(
        \pc_lut[19][7] ), .QN(n1595) );
  DFFR_X1 \pc_lut_reg[19][5]  ( .D(n6916), .CK(Clk), .RN(n3860), .Q(
        \pc_lut[19][5] ), .QN(n1594) );
  DFFR_X1 \pc_lut_reg[19][1]  ( .D(n6914), .CK(Clk), .RN(n3938), .Q(
        \pc_lut[19][1] ) );
  DFFR_X1 \pc_lut_reg[19][0]  ( .D(n6913), .CK(Clk), .RN(n3938), .Q(
        \pc_lut[19][0] ) );
  DFFR_X1 \pc_lut_reg[19][4]  ( .D(n6911), .CK(Clk), .RN(n3938), .Q(
        \pc_lut[19][4] ) );
  DFFR_X1 \pc_lut_reg[19][6]  ( .D(n6910), .CK(Clk), .RN(n3939), .Q(
        \pc_lut[19][6] ), .QN(n1590) );
  DFFR_X1 \pc_lut_reg[19][8]  ( .D(n6909), .CK(Clk), .RN(n3939), .Q(
        \pc_lut[19][8] ), .QN(n1589) );
  DFFR_X1 \pc_lut_reg[19][10]  ( .D(n6908), .CK(Clk), .RN(n3939), .Q(
        \pc_lut[19][10] ), .QN(n1588) );
  DFFR_X1 \pc_lut_reg[19][12]  ( .D(n6907), .CK(Clk), .RN(n3939), .Q(
        \pc_lut[19][12] ), .QN(n1587) );
  DFFR_X1 \pc_lut_reg[19][14]  ( .D(n6906), .CK(Clk), .RN(n3939), .Q(
        \pc_lut[19][14] ), .QN(n1586) );
  DFFR_X1 \pc_lut_reg[19][16]  ( .D(n6905), .CK(Clk), .RN(n3939), .Q(
        \pc_lut[19][16] ), .QN(n1585) );
  DFFR_X1 \pc_lut_reg[19][18]  ( .D(n6904), .CK(Clk), .RN(n3862), .Q(
        \pc_lut[19][18] ), .QN(n1584) );
  DFFR_X1 \pc_lut_reg[19][20]  ( .D(n6903), .CK(Clk), .RN(n3939), .Q(
        \pc_lut[19][20] ), .QN(n1583) );
  DFFR_X1 \pc_lut_reg[19][22]  ( .D(n6902), .CK(Clk), .RN(n3939), .Q(
        \pc_lut[19][22] ), .QN(n1582) );
  DFFR_X1 \pc_lut_reg[19][24]  ( .D(n6901), .CK(Clk), .RN(n3939), .Q(
        \pc_lut[19][24] ), .QN(n1581) );
  DFFR_X1 \pc_lut_reg[19][26]  ( .D(n6900), .CK(Clk), .RN(n3939), .Q(
        \pc_lut[19][26] ), .QN(n1580) );
  DFFR_X1 \pc_lut_reg[19][28]  ( .D(n6899), .CK(Clk), .RN(n3939), .Q(
        \pc_lut[19][28] ), .QN(n1579) );
  DFFR_X1 \pc_lut_reg[19][30]  ( .D(n6898), .CK(Clk), .RN(n3939), .Q(
        \pc_lut[19][30] ), .QN(n1577) );
  DFFR_X1 \pc_lut_reg[20][31]  ( .D(n6897), .CK(Clk), .RN(n3939), .Q(
        \pc_lut[20][31] ), .QN(n1575) );
  DFFR_X1 \pc_lut_reg[20][29]  ( .D(n6896), .CK(Clk), .RN(n3939), .Q(
        \pc_lut[20][29] ), .QN(n1574) );
  DFFR_X1 \pc_lut_reg[20][27]  ( .D(n6895), .CK(Clk), .RN(n3939), .Q(
        \pc_lut[20][27] ), .QN(n1573) );
  DFFR_X1 \pc_lut_reg[20][25]  ( .D(n6894), .CK(Clk), .RN(n3940), .Q(
        \pc_lut[20][25] ), .QN(n1572) );
  DFFR_X1 \pc_lut_reg[20][23]  ( .D(n6893), .CK(Clk), .RN(n3940), .Q(
        \pc_lut[20][23] ), .QN(n1571) );
  DFFR_X1 \pc_lut_reg[20][21]  ( .D(n6892), .CK(Clk), .RN(n3940), .Q(
        \pc_lut[20][21] ), .QN(n1570) );
  DFFR_X1 \pc_lut_reg[20][19]  ( .D(n6891), .CK(Clk), .RN(n3940), .Q(
        \pc_lut[20][19] ), .QN(n1569) );
  DFFR_X1 \pc_lut_reg[20][17]  ( .D(n6890), .CK(Clk), .RN(n3940), .Q(
        \pc_lut[20][17] ), .QN(n1568) );
  DFFR_X1 \pc_lut_reg[20][15]  ( .D(n6889), .CK(Clk), .RN(n3940), .Q(
        \pc_lut[20][15] ), .QN(n1567) );
  DFFR_X1 \pc_lut_reg[20][13]  ( .D(n6888), .CK(Clk), .RN(n3940), .Q(
        \pc_lut[20][13] ), .QN(n1566) );
  DFFR_X1 \pc_lut_reg[20][11]  ( .D(n6887), .CK(Clk), .RN(n3940), .Q(
        \pc_lut[20][11] ), .QN(n1565) );
  DFFR_X1 \pc_lut_reg[20][9]  ( .D(n6886), .CK(Clk), .RN(n3940), .Q(
        \pc_lut[20][9] ), .QN(n1564) );
  DFFR_X1 \pc_lut_reg[20][7]  ( .D(n6885), .CK(Clk), .RN(n3940), .Q(
        \pc_lut[20][7] ), .QN(n1563) );
  DFFR_X1 \pc_lut_reg[20][5]  ( .D(n6884), .CK(Clk), .RN(n3860), .Q(
        \pc_lut[20][5] ), .QN(n1562) );
  DFFR_X1 \pc_lut_reg[20][2]  ( .D(n6880), .CK(Clk), .RN(n3940), .Q(
        \pc_lut[20][2] ) );
  DFFR_X1 \pc_lut_reg[20][4]  ( .D(n6879), .CK(Clk), .RN(n3940), .Q(
        \pc_lut[20][4] ) );
  DFFR_X1 \pc_lut_reg[20][6]  ( .D(n6878), .CK(Clk), .RN(n3940), .Q(
        \pc_lut[20][6] ), .QN(n1559) );
  DFFR_X1 \pc_lut_reg[20][8]  ( .D(n6877), .CK(Clk), .RN(n3940), .Q(
        \pc_lut[20][8] ), .QN(n1558) );
  DFFR_X1 \pc_lut_reg[20][10]  ( .D(n6876), .CK(Clk), .RN(n3940), .Q(
        \pc_lut[20][10] ), .QN(n1557) );
  DFFR_X1 \pc_lut_reg[20][12]  ( .D(n6875), .CK(Clk), .RN(n3941), .Q(
        \pc_lut[20][12] ), .QN(n1556) );
  DFFR_X1 \pc_lut_reg[20][14]  ( .D(n6874), .CK(Clk), .RN(n3941), .Q(
        \pc_lut[20][14] ), .QN(n1555) );
  DFFR_X1 \pc_lut_reg[20][16]  ( .D(n6873), .CK(Clk), .RN(n3941), .Q(
        \pc_lut[20][16] ), .QN(n1554) );
  DFFR_X1 \pc_lut_reg[20][18]  ( .D(n6872), .CK(Clk), .RN(n3863), .Q(
        \pc_lut[20][18] ), .QN(n1553) );
  DFFR_X1 \pc_lut_reg[20][20]  ( .D(n6871), .CK(Clk), .RN(n3941), .Q(
        \pc_lut[20][20] ), .QN(n1552) );
  DFFR_X1 \pc_lut_reg[20][22]  ( .D(n6870), .CK(Clk), .RN(n3941), .Q(
        \pc_lut[20][22] ), .QN(n1551) );
  DFFR_X1 \pc_lut_reg[20][24]  ( .D(n6869), .CK(Clk), .RN(n3941), .Q(
        \pc_lut[20][24] ), .QN(n1550) );
  DFFR_X1 \pc_lut_reg[20][26]  ( .D(n6868), .CK(Clk), .RN(n3941), .Q(
        \pc_lut[20][26] ), .QN(n1549) );
  DFFR_X1 \pc_lut_reg[20][28]  ( .D(n6867), .CK(Clk), .RN(n3941), .Q(
        \pc_lut[20][28] ), .QN(n1548) );
  DFFR_X1 \pc_lut_reg[20][30]  ( .D(n6866), .CK(Clk), .RN(n3941), .Q(
        \pc_lut[20][30] ), .QN(n1546) );
  DFFR_X1 \pc_lut_reg[21][31]  ( .D(n6865), .CK(Clk), .RN(n3941), .Q(
        \pc_lut[21][31] ), .QN(n1544) );
  DFFR_X1 \pc_lut_reg[21][29]  ( .D(n6864), .CK(Clk), .RN(n3941), .Q(
        \pc_lut[21][29] ), .QN(n1543) );
  DFFR_X1 \pc_lut_reg[21][27]  ( .D(n6863), .CK(Clk), .RN(n3941), .Q(
        \pc_lut[21][27] ), .QN(n1542) );
  DFFR_X1 \pc_lut_reg[21][25]  ( .D(n6862), .CK(Clk), .RN(n3941), .Q(
        \pc_lut[21][25] ), .QN(n1541) );
  DFFR_X1 \pc_lut_reg[21][23]  ( .D(n6861), .CK(Clk), .RN(n3941), .Q(
        \pc_lut[21][23] ), .QN(n1540) );
  DFFR_X1 \pc_lut_reg[21][21]  ( .D(n6860), .CK(Clk), .RN(n3942), .Q(
        \pc_lut[21][21] ), .QN(n1539) );
  DFFR_X1 \pc_lut_reg[21][19]  ( .D(n6859), .CK(Clk), .RN(n3942), .Q(
        \pc_lut[21][19] ), .QN(n1538) );
  DFFR_X1 \pc_lut_reg[21][17]  ( .D(n6858), .CK(Clk), .RN(n3942), .Q(
        \pc_lut[21][17] ), .QN(n1537) );
  DFFR_X1 \pc_lut_reg[21][15]  ( .D(n6857), .CK(Clk), .RN(n3942), .Q(
        \pc_lut[21][15] ), .QN(n1536) );
  DFFR_X1 \pc_lut_reg[21][13]  ( .D(n6856), .CK(Clk), .RN(n3942), .Q(
        \pc_lut[21][13] ), .QN(n1535) );
  DFFR_X1 \pc_lut_reg[21][11]  ( .D(n6855), .CK(Clk), .RN(n3942), .Q(
        \pc_lut[21][11] ), .QN(n1534) );
  DFFR_X1 \pc_lut_reg[21][9]  ( .D(n6854), .CK(Clk), .RN(n3942), .Q(
        \pc_lut[21][9] ), .QN(n1533) );
  DFFR_X1 \pc_lut_reg[21][7]  ( .D(n6853), .CK(Clk), .RN(n3942), .Q(
        \pc_lut[21][7] ), .QN(n1532) );
  DFFR_X1 \pc_lut_reg[21][5]  ( .D(n6852), .CK(Clk), .RN(n3860), .Q(
        \pc_lut[21][5] ), .QN(n1531) );
  DFFR_X1 \pc_lut_reg[21][0]  ( .D(n6849), .CK(Clk), .RN(n3942), .Q(
        \pc_lut[21][0] ) );
  DFFR_X1 \pc_lut_reg[21][2]  ( .D(n6848), .CK(Clk), .RN(n3942), .Q(
        \pc_lut[21][2] ) );
  DFFR_X1 \pc_lut_reg[21][4]  ( .D(n6847), .CK(Clk), .RN(n3942), .Q(
        \pc_lut[21][4] ) );
  DFFR_X1 \pc_lut_reg[21][6]  ( .D(n6846), .CK(Clk), .RN(n3942), .Q(
        \pc_lut[21][6] ), .QN(n1527) );
  DFFR_X1 \pc_lut_reg[21][8]  ( .D(n6845), .CK(Clk), .RN(n3942), .Q(
        \pc_lut[21][8] ), .QN(n1526) );
  DFFR_X1 \pc_lut_reg[21][10]  ( .D(n6844), .CK(Clk), .RN(n3942), .Q(
        \pc_lut[21][10] ), .QN(n1525) );
  DFFR_X1 \pc_lut_reg[21][12]  ( .D(n6843), .CK(Clk), .RN(n3942), .Q(
        \pc_lut[21][12] ), .QN(n1524) );
  DFFR_X1 \pc_lut_reg[21][14]  ( .D(n6842), .CK(Clk), .RN(n3943), .Q(
        \pc_lut[21][14] ), .QN(n1523) );
  DFFR_X1 \pc_lut_reg[21][16]  ( .D(n6841), .CK(Clk), .RN(n3943), .Q(
        \pc_lut[21][16] ), .QN(n1522) );
  DFFR_X1 \pc_lut_reg[21][18]  ( .D(n6840), .CK(Clk), .RN(n3863), .Q(
        \pc_lut[21][18] ), .QN(n1521) );
  DFFR_X1 \pc_lut_reg[21][20]  ( .D(n6839), .CK(Clk), .RN(n3943), .Q(
        \pc_lut[21][20] ), .QN(n1520) );
  DFFR_X1 \pc_lut_reg[21][22]  ( .D(n6838), .CK(Clk), .RN(n3943), .Q(
        \pc_lut[21][22] ), .QN(n1519) );
  DFFR_X1 \pc_lut_reg[21][24]  ( .D(n6837), .CK(Clk), .RN(n3943), .Q(
        \pc_lut[21][24] ), .QN(n1518) );
  DFFR_X1 \pc_lut_reg[21][26]  ( .D(n6836), .CK(Clk), .RN(n3943), .Q(
        \pc_lut[21][26] ), .QN(n1517) );
  DFFR_X1 \pc_lut_reg[21][28]  ( .D(n6835), .CK(Clk), .RN(n3943), .Q(
        \pc_lut[21][28] ), .QN(n1516) );
  DFFR_X1 \pc_lut_reg[21][30]  ( .D(n6834), .CK(Clk), .RN(n3943), .Q(
        \pc_lut[21][30] ), .QN(n1514) );
  DFFR_X1 \pc_lut_reg[22][31]  ( .D(n6833), .CK(Clk), .RN(n3943), .QN(n1512)
         );
  DFFR_X1 \pc_lut_reg[22][29]  ( .D(n6832), .CK(Clk), .RN(n3943), .QN(n1511)
         );
  DFFR_X1 \pc_lut_reg[22][27]  ( .D(n6831), .CK(Clk), .RN(n3943), .QN(n1510)
         );
  DFFR_X1 \pc_lut_reg[22][25]  ( .D(n6830), .CK(Clk), .RN(n3943), .QN(n1509)
         );
  DFFR_X1 \pc_lut_reg[22][23]  ( .D(n6829), .CK(Clk), .RN(n3943), .QN(n1508)
         );
  DFFR_X1 \pc_lut_reg[22][21]  ( .D(n6828), .CK(Clk), .RN(n3943), .QN(n1507)
         );
  DFFR_X1 \pc_lut_reg[22][19]  ( .D(n6827), .CK(Clk), .RN(n3943), .QN(n1506)
         );
  DFFR_X1 \pc_lut_reg[22][17]  ( .D(n6826), .CK(Clk), .RN(n3944), .QN(n1505)
         );
  DFFR_X1 \pc_lut_reg[22][15]  ( .D(n6825), .CK(Clk), .RN(n3944), .QN(n1504)
         );
  DFFR_X1 \pc_lut_reg[22][13]  ( .D(n6824), .CK(Clk), .RN(n3944), .QN(n1503)
         );
  DFFR_X1 \pc_lut_reg[22][11]  ( .D(n6823), .CK(Clk), .RN(n3944), .QN(n1502)
         );
  DFFR_X1 \pc_lut_reg[22][9]  ( .D(n6822), .CK(Clk), .RN(n3944), .QN(n1501) );
  DFFR_X1 \pc_lut_reg[22][7]  ( .D(n6821), .CK(Clk), .RN(n3944), .QN(n1500) );
  DFFR_X1 \pc_lut_reg[22][5]  ( .D(n6820), .CK(Clk), .RN(n3860), .QN(n1499) );
  DFFR_X1 \pc_lut_reg[22][1]  ( .D(n6818), .CK(Clk), .RN(n3944), .QN(n1497) );
  DFFR_X1 \pc_lut_reg[22][2]  ( .D(n6816), .CK(Clk), .RN(n3944), .QN(n1495) );
  DFFR_X1 \pc_lut_reg[22][4]  ( .D(n6815), .CK(Clk), .RN(n3944), .QN(n1494) );
  DFFR_X1 \pc_lut_reg[22][6]  ( .D(n6814), .CK(Clk), .RN(n3944), .QN(n1493) );
  DFFR_X1 \pc_lut_reg[22][8]  ( .D(n6813), .CK(Clk), .RN(n3944), .QN(n1492) );
  DFFR_X1 \pc_lut_reg[22][10]  ( .D(n6812), .CK(Clk), .RN(n3944), .QN(n1491)
         );
  DFFR_X1 \pc_lut_reg[22][12]  ( .D(n6811), .CK(Clk), .RN(n3944), .QN(n1490)
         );
  DFFR_X1 \pc_lut_reg[22][14]  ( .D(n6810), .CK(Clk), .RN(n3944), .QN(n1489)
         );
  DFFR_X1 \pc_lut_reg[22][16]  ( .D(n6809), .CK(Clk), .RN(n3945), .QN(n1488)
         );
  DFFR_X1 \pc_lut_reg[22][18]  ( .D(n6808), .CK(Clk), .RN(n3863), .QN(n1487)
         );
  DFFR_X1 \pc_lut_reg[22][20]  ( .D(n6807), .CK(Clk), .RN(n3945), .QN(n1486)
         );
  DFFR_X1 \pc_lut_reg[22][22]  ( .D(n6806), .CK(Clk), .RN(n3944), .QN(n1485)
         );
  DFFR_X1 \pc_lut_reg[22][24]  ( .D(n6805), .CK(Clk), .RN(n3945), .QN(n1484)
         );
  DFFR_X1 \pc_lut_reg[22][26]  ( .D(n6804), .CK(Clk), .RN(n3945), .QN(n1483)
         );
  DFFR_X1 \pc_lut_reg[22][28]  ( .D(n6803), .CK(Clk), .RN(n3945), .QN(n1482)
         );
  DFFR_X1 \pc_lut_reg[22][30]  ( .D(n6802), .CK(Clk), .RN(n3945), .QN(n1480)
         );
  DFFR_X1 \pc_lut_reg[23][31]  ( .D(n6801), .CK(Clk), .RN(n3904), .QN(n1477)
         );
  DFFR_X1 \pc_lut_reg[23][29]  ( .D(n6800), .CK(Clk), .RN(n3900), .QN(n1476)
         );
  DFFR_X1 \pc_lut_reg[23][27]  ( .D(n6799), .CK(Clk), .RN(n3896), .QN(n1475)
         );
  DFFR_X1 \pc_lut_reg[23][25]  ( .D(n6798), .CK(Clk), .RN(n3896), .QN(n1474)
         );
  DFFR_X1 \pc_lut_reg[23][23]  ( .D(n6797), .CK(Clk), .RN(n3896), .QN(n1473)
         );
  DFFR_X1 \pc_lut_reg[23][21]  ( .D(n6796), .CK(Clk), .RN(n3896), .QN(n1472)
         );
  DFFR_X1 \pc_lut_reg[23][19]  ( .D(n6795), .CK(Clk), .RN(n3896), .QN(n1471)
         );
  DFFR_X1 \pc_lut_reg[23][17]  ( .D(n6794), .CK(Clk), .RN(n3896), .QN(n1470)
         );
  DFFR_X1 \pc_lut_reg[23][15]  ( .D(n6793), .CK(Clk), .RN(n3896), .QN(n1469)
         );
  DFFR_X1 \pc_lut_reg[23][13]  ( .D(n6792), .CK(Clk), .RN(n3896), .QN(n1468)
         );
  DFFR_X1 \pc_lut_reg[23][11]  ( .D(n6791), .CK(Clk), .RN(n3897), .QN(n1467)
         );
  DFFR_X1 \pc_lut_reg[23][9]  ( .D(n6790), .CK(Clk), .RN(n3897), .QN(n1466) );
  DFFR_X1 \pc_lut_reg[23][7]  ( .D(n6789), .CK(Clk), .RN(n3934), .QN(n1465) );
  DFFR_X1 \pc_lut_reg[23][5]  ( .D(n6788), .CK(Clk), .RN(n3860), .QN(n1464) );
  DFFR_X1 \pc_lut_reg[23][1]  ( .D(n6786), .CK(Clk), .RN(n3934), .QN(n1462) );
  DFFR_X1 \pc_lut_reg[23][0]  ( .D(n6785), .CK(Clk), .RN(n3934), .QN(n1461) );
  DFFR_X1 \pc_lut_reg[23][2]  ( .D(n6784), .CK(Clk), .RN(n3934), .QN(n1460) );
  DFFR_X1 \pc_lut_reg[23][4]  ( .D(n6783), .CK(Clk), .RN(n3934), .QN(n1459) );
  DFFR_X1 \pc_lut_reg[23][6]  ( .D(n6782), .CK(Clk), .RN(n3934), .QN(n1458) );
  DFFR_X1 \pc_lut_reg[23][8]  ( .D(n6781), .CK(Clk), .RN(n3934), .QN(n1457) );
  DFFR_X1 \pc_lut_reg[23][10]  ( .D(n6780), .CK(Clk), .RN(n3934), .QN(n1456)
         );
  DFFR_X1 \pc_lut_reg[23][12]  ( .D(n6779), .CK(Clk), .RN(n3934), .QN(n1455)
         );
  DFFR_X1 \pc_lut_reg[23][14]  ( .D(n6778), .CK(Clk), .RN(n3934), .QN(n1454)
         );
  DFFR_X1 \pc_lut_reg[23][16]  ( .D(n6777), .CK(Clk), .RN(n3934), .QN(n1453)
         );
  DFFR_X1 \pc_lut_reg[23][18]  ( .D(n6776), .CK(Clk), .RN(n3863), .QN(n1452)
         );
  DFFR_X1 \pc_lut_reg[23][20]  ( .D(n6775), .CK(Clk), .RN(n3934), .QN(n1451)
         );
  DFFR_X1 \pc_lut_reg[23][22]  ( .D(n6774), .CK(Clk), .RN(n3934), .QN(n1450)
         );
  DFFR_X1 \pc_lut_reg[23][24]  ( .D(n6773), .CK(Clk), .RN(n3934), .QN(n1449)
         );
  DFFR_X1 \pc_lut_reg[23][26]  ( .D(n6772), .CK(Clk), .RN(n3934), .QN(n1448)
         );
  DFFR_X1 \pc_lut_reg[23][28]  ( .D(n6771), .CK(Clk), .RN(n3935), .QN(n1447)
         );
  DFFR_X1 \pc_lut_reg[23][30]  ( .D(n6770), .CK(Clk), .RN(n3935), .QN(n1445)
         );
  DFFR_X1 \pc_lut_reg[24][31]  ( .D(n6769), .CK(Clk), .RN(n3935), .QN(n1443)
         );
  DFFR_X1 \pc_lut_reg[24][29]  ( .D(n6768), .CK(Clk), .RN(n3935), .QN(n1442)
         );
  DFFR_X1 \pc_lut_reg[24][27]  ( .D(n6767), .CK(Clk), .RN(n3935), .QN(n1441)
         );
  DFFR_X1 \pc_lut_reg[24][25]  ( .D(n6766), .CK(Clk), .RN(n3935), .QN(n1440)
         );
  DFFR_X1 \pc_lut_reg[24][23]  ( .D(n6765), .CK(Clk), .RN(n3935), .QN(n1439)
         );
  DFFR_X1 \pc_lut_reg[24][21]  ( .D(n6764), .CK(Clk), .RN(n3935), .QN(n1438)
         );
  DFFR_X1 \pc_lut_reg[24][19]  ( .D(n6763), .CK(Clk), .RN(n3935), .QN(n1437)
         );
  DFFR_X1 \pc_lut_reg[24][17]  ( .D(n6762), .CK(Clk), .RN(n3935), .QN(n1436)
         );
  DFFR_X1 \pc_lut_reg[24][15]  ( .D(n6761), .CK(Clk), .RN(n3935), .QN(n1435)
         );
  DFFR_X1 \pc_lut_reg[24][13]  ( .D(n6760), .CK(Clk), .RN(n3935), .QN(n1434)
         );
  DFFR_X1 \pc_lut_reg[24][11]  ( .D(n6759), .CK(Clk), .RN(n3935), .QN(n1433)
         );
  DFFR_X1 \pc_lut_reg[24][9]  ( .D(n6758), .CK(Clk), .RN(n3935), .QN(n1432) );
  DFFR_X1 \pc_lut_reg[24][7]  ( .D(n6757), .CK(Clk), .RN(n3935), .QN(n1431) );
  DFFR_X1 \pc_lut_reg[24][5]  ( .D(n6756), .CK(Clk), .RN(n3860), .QN(n1430) );
  DFFR_X1 \pc_lut_reg[24][3]  ( .D(n6755), .CK(Clk), .RN(n3936), .QN(n1429) );
  DFFR_X1 \pc_lut_reg[24][4]  ( .D(n6751), .CK(Clk), .RN(n3936), .QN(n1425) );
  DFFR_X1 \pc_lut_reg[24][6]  ( .D(n6750), .CK(Clk), .RN(n3936), .QN(n1424) );
  DFFR_X1 \pc_lut_reg[24][8]  ( .D(n6749), .CK(Clk), .RN(n3936), .QN(n1423) );
  DFFR_X1 \pc_lut_reg[24][10]  ( .D(n6748), .CK(Clk), .RN(n3936), .QN(n1422)
         );
  DFFR_X1 \pc_lut_reg[24][12]  ( .D(n6747), .CK(Clk), .RN(n3936), .QN(n1421)
         );
  DFFR_X1 \pc_lut_reg[24][14]  ( .D(n6746), .CK(Clk), .RN(n3936), .QN(n1420)
         );
  DFFR_X1 \pc_lut_reg[24][16]  ( .D(n6745), .CK(Clk), .RN(n3936), .QN(n1419)
         );
  DFFR_X1 \pc_lut_reg[24][18]  ( .D(n6744), .CK(Clk), .RN(n3863), .QN(n1418)
         );
  DFFR_X1 \pc_lut_reg[24][20]  ( .D(n6743), .CK(Clk), .RN(n3936), .QN(n1417)
         );
  DFFR_X1 \pc_lut_reg[24][22]  ( .D(n6742), .CK(Clk), .RN(n3936), .QN(n1416)
         );
  DFFR_X1 \pc_lut_reg[24][24]  ( .D(n6741), .CK(Clk), .RN(n3936), .QN(n1415)
         );
  DFFR_X1 \pc_lut_reg[24][26]  ( .D(n6740), .CK(Clk), .RN(n3936), .QN(n1414)
         );
  DFFR_X1 \pc_lut_reg[24][28]  ( .D(n6739), .CK(Clk), .RN(n3936), .QN(n1413)
         );
  DFFR_X1 \pc_lut_reg[24][30]  ( .D(n6738), .CK(Clk), .RN(n3936), .QN(n1411)
         );
  DFFR_X1 \pc_lut_reg[25][31]  ( .D(n6737), .CK(Clk), .RN(n3936), .QN(n1409)
         );
  DFFR_X1 \pc_lut_reg[25][29]  ( .D(n6736), .CK(Clk), .RN(n3937), .QN(n1408)
         );
  DFFR_X1 \pc_lut_reg[25][27]  ( .D(n6735), .CK(Clk), .RN(n3937), .QN(n1407)
         );
  DFFR_X1 \pc_lut_reg[25][25]  ( .D(n6734), .CK(Clk), .RN(n3937), .QN(n1406)
         );
  DFFR_X1 \pc_lut_reg[25][23]  ( .D(n6733), .CK(Clk), .RN(n3937), .QN(n1405)
         );
  DFFR_X1 \pc_lut_reg[25][21]  ( .D(n6732), .CK(Clk), .RN(n3925), .QN(n1404)
         );
  DFFR_X1 \pc_lut_reg[25][19]  ( .D(n6731), .CK(Clk), .RN(n3921), .QN(n1403)
         );
  DFFR_X1 \pc_lut_reg[25][17]  ( .D(n6730), .CK(Clk), .RN(n3921), .QN(n1402)
         );
  DFFR_X1 \pc_lut_reg[25][15]  ( .D(n6729), .CK(Clk), .RN(n3921), .QN(n1401)
         );
  DFFR_X1 \pc_lut_reg[25][13]  ( .D(n6728), .CK(Clk), .RN(n3921), .QN(n1400)
         );
  DFFR_X1 \pc_lut_reg[25][11]  ( .D(n6727), .CK(Clk), .RN(n3921), .QN(n1399)
         );
  DFFR_X1 \pc_lut_reg[25][9]  ( .D(n6726), .CK(Clk), .RN(n3921), .QN(n1398) );
  DFFR_X1 \pc_lut_reg[25][7]  ( .D(n6725), .CK(Clk), .RN(n3921), .QN(n1397) );
  DFFR_X1 \pc_lut_reg[25][5]  ( .D(n6724), .CK(Clk), .RN(n3860), .QN(n1396) );
  DFFR_X1 \pc_lut_reg[25][3]  ( .D(n6723), .CK(Clk), .RN(n3921), .QN(n1395) );
  DFFR_X1 \pc_lut_reg[25][0]  ( .D(n6721), .CK(Clk), .RN(n3921), .QN(n1393) );
  DFFR_X1 \pc_lut_reg[25][4]  ( .D(n6719), .CK(Clk), .RN(n3921), .QN(n1391) );
  DFFR_X1 \pc_lut_reg[25][6]  ( .D(n6718), .CK(Clk), .RN(n3921), .QN(n1390) );
  DFFR_X1 \pc_lut_reg[25][8]  ( .D(n6717), .CK(Clk), .RN(n3921), .QN(n1389) );
  DFFR_X1 \pc_lut_reg[25][10]  ( .D(n6716), .CK(Clk), .RN(n3921), .QN(n1388)
         );
  DFFR_X1 \pc_lut_reg[25][12]  ( .D(n6715), .CK(Clk), .RN(n3921), .QN(n1387)
         );
  DFFR_X1 \pc_lut_reg[25][14]  ( .D(n6714), .CK(Clk), .RN(n3922), .QN(n1386)
         );
  DFFR_X1 \pc_lut_reg[25][16]  ( .D(n6713), .CK(Clk), .RN(n3922), .QN(n1385)
         );
  DFFR_X1 \pc_lut_reg[25][18]  ( .D(n6712), .CK(Clk), .RN(n3863), .QN(n1384)
         );
  DFFR_X1 \pc_lut_reg[25][20]  ( .D(n6711), .CK(Clk), .RN(n3922), .QN(n1383)
         );
  DFFR_X1 \pc_lut_reg[25][22]  ( .D(n6710), .CK(Clk), .RN(n3922), .QN(n1382)
         );
  DFFR_X1 \pc_lut_reg[25][24]  ( .D(n6709), .CK(Clk), .RN(n3922), .QN(n1381)
         );
  DFFR_X1 \pc_lut_reg[25][26]  ( .D(n6708), .CK(Clk), .RN(n3922), .QN(n1380)
         );
  DFFR_X1 \pc_lut_reg[25][28]  ( .D(n6707), .CK(Clk), .RN(n3922), .QN(n1379)
         );
  DFFR_X1 \pc_lut_reg[25][30]  ( .D(n6706), .CK(Clk), .RN(n3922), .QN(n1377)
         );
  DFFR_X1 \pc_lut_reg[26][31]  ( .D(n6705), .CK(Clk), .RN(n3922), .Q(
        \pc_lut[26][31] ), .QN(n1375) );
  DFFR_X1 \pc_lut_reg[26][29]  ( .D(n6704), .CK(Clk), .RN(n3922), .Q(
        \pc_lut[26][29] ), .QN(n1374) );
  DFFR_X1 \pc_lut_reg[26][27]  ( .D(n6703), .CK(Clk), .RN(n3922), .Q(
        \pc_lut[26][27] ), .QN(n1373) );
  DFFR_X1 \pc_lut_reg[26][25]  ( .D(n6702), .CK(Clk), .RN(n3922), .Q(
        \pc_lut[26][25] ), .QN(n1372) );
  DFFR_X1 \pc_lut_reg[26][23]  ( .D(n6701), .CK(Clk), .RN(n3922), .Q(
        \pc_lut[26][23] ), .QN(n1371) );
  DFFR_X1 \pc_lut_reg[26][21]  ( .D(n6700), .CK(Clk), .RN(n3922), .Q(
        \pc_lut[26][21] ), .QN(n1370) );
  DFFR_X1 \pc_lut_reg[26][19]  ( .D(n6699), .CK(Clk), .RN(n3922), .Q(
        \pc_lut[26][19] ), .QN(n1369) );
  DFFR_X1 \pc_lut_reg[26][17]  ( .D(n6698), .CK(Clk), .RN(n3923), .Q(
        \pc_lut[26][17] ), .QN(n1368) );
  DFFR_X1 \pc_lut_reg[26][15]  ( .D(n6697), .CK(Clk), .RN(n3923), .Q(
        \pc_lut[26][15] ), .QN(n1367) );
  DFFR_X1 \pc_lut_reg[26][13]  ( .D(n6696), .CK(Clk), .RN(n3923), .Q(
        \pc_lut[26][13] ), .QN(n1366) );
  DFFR_X1 \pc_lut_reg[26][11]  ( .D(n6695), .CK(Clk), .RN(n3923), .Q(
        \pc_lut[26][11] ), .QN(n1365) );
  DFFR_X1 \pc_lut_reg[26][9]  ( .D(n6694), .CK(Clk), .RN(n3923), .Q(
        \pc_lut[26][9] ), .QN(n1364) );
  DFFR_X1 \pc_lut_reg[26][7]  ( .D(n6693), .CK(Clk), .RN(n3923), .Q(
        \pc_lut[26][7] ), .QN(n1363) );
  DFFR_X1 \pc_lut_reg[26][5]  ( .D(n6692), .CK(Clk), .RN(n3860), .Q(
        \pc_lut[26][5] ), .QN(n1362) );
  DFFR_X1 \pc_lut_reg[26][6]  ( .D(n6686), .CK(Clk), .RN(n3923), .Q(
        \pc_lut[26][6] ), .QN(n1358) );
  DFFR_X1 \pc_lut_reg[26][8]  ( .D(n6685), .CK(Clk), .RN(n3923), .Q(
        \pc_lut[26][8] ), .QN(n1357) );
  DFFR_X1 \pc_lut_reg[26][10]  ( .D(n6684), .CK(Clk), .RN(n3923), .Q(
        \pc_lut[26][10] ), .QN(n1356) );
  DFFR_X1 \pc_lut_reg[26][12]  ( .D(n6683), .CK(Clk), .RN(n3923), .Q(
        \pc_lut[26][12] ), .QN(n1355) );
  DFFR_X1 \pc_lut_reg[26][14]  ( .D(n6682), .CK(Clk), .RN(n3923), .Q(
        \pc_lut[26][14] ), .QN(n1354) );
  DFFR_X1 \pc_lut_reg[26][16]  ( .D(n6681), .CK(Clk), .RN(n3923), .Q(
        \pc_lut[26][16] ), .QN(n1353) );
  DFFR_X1 \pc_lut_reg[26][18]  ( .D(n6680), .CK(Clk), .RN(n3863), .Q(
        \pc_lut[26][18] ), .QN(n1352) );
  DFFR_X1 \pc_lut_reg[26][20]  ( .D(n6679), .CK(Clk), .RN(n3923), .Q(
        \pc_lut[26][20] ), .QN(n1351) );
  DFFR_X1 \pc_lut_reg[26][22]  ( .D(n6678), .CK(Clk), .RN(n3923), .Q(
        \pc_lut[26][22] ), .QN(n1350) );
  DFFR_X1 \pc_lut_reg[26][24]  ( .D(n6677), .CK(Clk), .RN(n3923), .Q(
        \pc_lut[26][24] ), .QN(n1349) );
  DFFR_X1 \pc_lut_reg[26][26]  ( .D(n6676), .CK(Clk), .RN(n3924), .Q(
        \pc_lut[26][26] ), .QN(n1348) );
  DFFR_X1 \pc_lut_reg[26][28]  ( .D(n6675), .CK(Clk), .RN(n3924), .Q(
        \pc_lut[26][28] ), .QN(n1347) );
  DFFR_X1 \pc_lut_reg[26][30]  ( .D(n6674), .CK(Clk), .RN(n3924), .Q(
        \pc_lut[26][30] ), .QN(n1345) );
  DFFR_X1 \pc_lut_reg[27][31]  ( .D(n6673), .CK(Clk), .RN(n3924), .Q(
        \pc_lut[27][31] ), .QN(n1342) );
  DFFR_X1 \pc_lut_reg[27][29]  ( .D(n6672), .CK(Clk), .RN(n3924), .Q(
        \pc_lut[27][29] ), .QN(n1341) );
  DFFR_X1 \pc_lut_reg[27][27]  ( .D(n6671), .CK(Clk), .RN(n3924), .Q(
        \pc_lut[27][27] ), .QN(n1340) );
  DFFR_X1 \pc_lut_reg[27][25]  ( .D(n6670), .CK(Clk), .RN(n3924), .Q(
        \pc_lut[27][25] ), .QN(n1339) );
  DFFR_X1 \pc_lut_reg[27][23]  ( .D(n6669), .CK(Clk), .RN(n3924), .Q(
        \pc_lut[27][23] ), .QN(n1338) );
  DFFR_X1 \pc_lut_reg[27][21]  ( .D(n6668), .CK(Clk), .RN(n3924), .Q(
        \pc_lut[27][21] ), .QN(n1337) );
  DFFR_X1 \pc_lut_reg[27][19]  ( .D(n6667), .CK(Clk), .RN(n3924), .Q(
        \pc_lut[27][19] ), .QN(n1336) );
  DFFR_X1 \pc_lut_reg[27][17]  ( .D(n6666), .CK(Clk), .RN(n3924), .Q(
        \pc_lut[27][17] ), .QN(n1335) );
  DFFR_X1 \pc_lut_reg[27][15]  ( .D(n6665), .CK(Clk), .RN(n3924), .Q(
        \pc_lut[27][15] ), .QN(n1334) );
  DFFR_X1 \pc_lut_reg[27][13]  ( .D(n6664), .CK(Clk), .RN(n3924), .Q(
        \pc_lut[27][13] ), .QN(n1333) );
  DFFR_X1 \pc_lut_reg[27][11]  ( .D(n6663), .CK(Clk), .RN(n3924), .Q(
        \pc_lut[27][11] ), .QN(n1332) );
  DFFR_X1 \pc_lut_reg[27][9]  ( .D(n6662), .CK(Clk), .RN(n3924), .Q(
        \pc_lut[27][9] ), .QN(n1331) );
  DFFR_X1 \pc_lut_reg[27][7]  ( .D(n6661), .CK(Clk), .RN(n3925), .Q(
        \pc_lut[27][7] ), .QN(n1330) );
  DFFR_X1 \pc_lut_reg[27][5]  ( .D(n6660), .CK(Clk), .RN(n3860), .Q(
        \pc_lut[27][5] ), .QN(n1329) );
  DFFR_X1 \pc_lut_reg[27][6]  ( .D(n6654), .CK(Clk), .RN(n3925), .Q(
        \pc_lut[27][6] ), .QN(n1324) );
  DFFR_X1 \pc_lut_reg[27][8]  ( .D(n6653), .CK(Clk), .RN(n3925), .Q(
        \pc_lut[27][8] ), .QN(n1323) );
  DFFR_X1 \pc_lut_reg[27][10]  ( .D(n6652), .CK(Clk), .RN(n3925), .Q(
        \pc_lut[27][10] ), .QN(n1322) );
  DFFR_X1 \pc_lut_reg[27][12]  ( .D(n6651), .CK(Clk), .RN(n3925), .Q(
        \pc_lut[27][12] ), .QN(n1321) );
  DFFR_X1 \pc_lut_reg[27][14]  ( .D(n6650), .CK(Clk), .RN(n3925), .Q(
        \pc_lut[27][14] ), .QN(n1320) );
  DFFR_X1 \pc_lut_reg[27][16]  ( .D(n6649), .CK(Clk), .RN(n3925), .Q(
        \pc_lut[27][16] ), .QN(n1319) );
  DFFR_X1 \pc_lut_reg[27][18]  ( .D(n6648), .CK(Clk), .RN(n3863), .Q(
        \pc_lut[27][18] ), .QN(n1318) );
  DFFR_X1 \pc_lut_reg[27][20]  ( .D(n6647), .CK(Clk), .RN(n3925), .Q(
        \pc_lut[27][20] ), .QN(n1317) );
  DFFR_X1 \pc_lut_reg[27][22]  ( .D(n6646), .CK(Clk), .RN(n3925), .Q(
        \pc_lut[27][22] ), .QN(n1316) );
  DFFR_X1 \pc_lut_reg[27][24]  ( .D(n6645), .CK(Clk), .RN(n3925), .Q(
        \pc_lut[27][24] ), .QN(n1315) );
  DFFR_X1 \pc_lut_reg[27][26]  ( .D(n6644), .CK(Clk), .RN(n3926), .Q(
        \pc_lut[27][26] ), .QN(n1314) );
  DFFR_X1 \pc_lut_reg[27][28]  ( .D(n6643), .CK(Clk), .RN(n3926), .Q(
        \pc_lut[27][28] ), .QN(n1313) );
  DFFR_X1 \pc_lut_reg[27][30]  ( .D(n6642), .CK(Clk), .RN(n3926), .Q(
        \pc_lut[27][30] ), .QN(n1311) );
  DFFR_X1 \pc_lut_reg[28][31]  ( .D(n6641), .CK(Clk), .RN(n3926), .QN(n1308)
         );
  DFFR_X1 \pc_lut_reg[28][29]  ( .D(n6640), .CK(Clk), .RN(n3926), .QN(n1307)
         );
  DFFR_X1 \pc_lut_reg[28][27]  ( .D(n6639), .CK(Clk), .RN(n3926), .QN(n1306)
         );
  DFFR_X1 \pc_lut_reg[28][25]  ( .D(n6638), .CK(Clk), .RN(n3926), .QN(n1305)
         );
  DFFR_X1 \pc_lut_reg[28][23]  ( .D(n6637), .CK(Clk), .RN(n3926), .QN(n1304)
         );
  DFFR_X1 \pc_lut_reg[28][21]  ( .D(n6636), .CK(Clk), .RN(n3926), .QN(n1303)
         );
  DFFR_X1 \pc_lut_reg[28][19]  ( .D(n6635), .CK(Clk), .RN(n3926), .QN(n1302)
         );
  DFFR_X1 \pc_lut_reg[28][17]  ( .D(n6634), .CK(Clk), .RN(n3926), .QN(n1301)
         );
  DFFR_X1 \pc_lut_reg[28][15]  ( .D(n6633), .CK(Clk), .RN(n3926), .QN(n1300)
         );
  DFFR_X1 \pc_lut_reg[28][13]  ( .D(n6632), .CK(Clk), .RN(n3926), .QN(n1299)
         );
  DFFR_X1 \pc_lut_reg[28][11]  ( .D(n6631), .CK(Clk), .RN(n3926), .QN(n1298)
         );
  DFFR_X1 \pc_lut_reg[28][9]  ( .D(n6630), .CK(Clk), .RN(n3926), .QN(n1297) );
  DFFR_X1 \pc_lut_reg[28][7]  ( .D(n6629), .CK(Clk), .RN(n3927), .QN(n1296) );
  DFFR_X1 \pc_lut_reg[28][5]  ( .D(n6628), .CK(Clk), .RN(n3860), .QN(n1295) );
  DFFR_X1 \pc_lut_reg[28][6]  ( .D(n6622), .CK(Clk), .RN(n3927), .QN(n1289) );
  DFFR_X1 \pc_lut_reg[28][8]  ( .D(n6621), .CK(Clk), .RN(n3927), .QN(n1288) );
  DFFR_X1 \pc_lut_reg[28][10]  ( .D(n6620), .CK(Clk), .RN(n3927), .QN(n1287)
         );
  DFFR_X1 \pc_lut_reg[28][12]  ( .D(n6619), .CK(Clk), .RN(n3927), .QN(n1286)
         );
  DFFR_X1 \pc_lut_reg[28][14]  ( .D(n6618), .CK(Clk), .RN(n3927), .QN(n1285)
         );
  DFFR_X1 \pc_lut_reg[28][16]  ( .D(n6617), .CK(Clk), .RN(n3927), .QN(n1284)
         );
  DFFR_X1 \pc_lut_reg[28][18]  ( .D(n6616), .CK(Clk), .RN(n3863), .QN(n1283)
         );
  DFFR_X1 \pc_lut_reg[28][20]  ( .D(n6615), .CK(Clk), .RN(n3927), .QN(n1282)
         );
  DFFR_X1 \pc_lut_reg[28][22]  ( .D(n6614), .CK(Clk), .RN(n3927), .QN(n1281)
         );
  DFFR_X1 \pc_lut_reg[28][24]  ( .D(n6613), .CK(Clk), .RN(n3927), .QN(n1280)
         );
  DFFR_X1 \pc_lut_reg[28][26]  ( .D(n6612), .CK(Clk), .RN(n3927), .QN(n1279)
         );
  DFFR_X1 \pc_lut_reg[28][28]  ( .D(n6611), .CK(Clk), .RN(n3927), .QN(n1278)
         );
  DFFR_X1 \pc_lut_reg[28][30]  ( .D(n6610), .CK(Clk), .RN(n3927), .QN(n1276)
         );
  DFFR_X1 \pc_lut_reg[29][31]  ( .D(n6609), .CK(Clk), .RN(n3927), .QN(n1274)
         );
  DFFR_X1 \pc_lut_reg[29][29]  ( .D(n6608), .CK(Clk), .RN(n3927), .QN(n1273)
         );
  DFFR_X1 \pc_lut_reg[29][27]  ( .D(n6607), .CK(Clk), .RN(n3928), .QN(n1272)
         );
  DFFR_X1 \pc_lut_reg[29][25]  ( .D(n6606), .CK(Clk), .RN(n3928), .QN(n1271)
         );
  DFFR_X1 \pc_lut_reg[29][23]  ( .D(n6605), .CK(Clk), .RN(n3928), .QN(n1270)
         );
  DFFR_X1 \pc_lut_reg[29][21]  ( .D(n6604), .CK(Clk), .RN(n3928), .QN(n1269)
         );
  DFFR_X1 \pc_lut_reg[29][19]  ( .D(n6603), .CK(Clk), .RN(n3928), .QN(n1268)
         );
  DFFR_X1 \pc_lut_reg[29][17]  ( .D(n6602), .CK(Clk), .RN(n3928), .QN(n1267)
         );
  DFFR_X1 \pc_lut_reg[29][15]  ( .D(n6601), .CK(Clk), .RN(n3928), .QN(n1266)
         );
  DFFR_X1 \pc_lut_reg[29][13]  ( .D(n6600), .CK(Clk), .RN(n3928), .QN(n1265)
         );
  DFFR_X1 \pc_lut_reg[29][11]  ( .D(n6599), .CK(Clk), .RN(n3928), .QN(n1264)
         );
  DFFR_X1 \pc_lut_reg[29][9]  ( .D(n6598), .CK(Clk), .RN(n3928), .QN(n1263) );
  DFFR_X1 \pc_lut_reg[29][7]  ( .D(n6597), .CK(Clk), .RN(n3928), .QN(n1262) );
  DFFR_X1 \pc_lut_reg[29][5]  ( .D(n6596), .CK(Clk), .RN(n3860), .QN(n1261) );
  DFFR_X1 \pc_lut_reg[29][6]  ( .D(n6590), .CK(Clk), .RN(n3928), .QN(n1254) );
  DFFR_X1 \pc_lut_reg[29][8]  ( .D(n6589), .CK(Clk), .RN(n3928), .QN(n1253) );
  DFFR_X1 \pc_lut_reg[29][10]  ( .D(n6588), .CK(Clk), .RN(n3928), .QN(n1252)
         );
  DFFR_X1 \pc_lut_reg[29][12]  ( .D(n6587), .CK(Clk), .RN(n3928), .QN(n1251)
         );
  DFFR_X1 \pc_lut_reg[29][14]  ( .D(n6586), .CK(Clk), .RN(n3929), .QN(n1250)
         );
  DFFR_X1 \pc_lut_reg[29][16]  ( .D(n6585), .CK(Clk), .RN(n3929), .QN(n1249)
         );
  DFFR_X1 \pc_lut_reg[29][18]  ( .D(n6584), .CK(Clk), .RN(n3884), .QN(n1248)
         );
  DFFR_X1 \pc_lut_reg[29][20]  ( .D(n6583), .CK(Clk), .RN(n3929), .QN(n1247)
         );
  DFFR_X1 \pc_lut_reg[29][22]  ( .D(n6582), .CK(Clk), .RN(n3949), .QN(n1246)
         );
  DFFR_X1 \pc_lut_reg[29][24]  ( .D(n6581), .CK(Clk), .RN(n3945), .QN(n1245)
         );
  DFFR_X1 \pc_lut_reg[29][26]  ( .D(n6580), .CK(Clk), .RN(n3945), .QN(n1244)
         );
  DFFR_X1 \pc_lut_reg[29][28]  ( .D(n6579), .CK(Clk), .RN(n3945), .QN(n1243)
         );
  DFFR_X1 \pc_lut_reg[29][30]  ( .D(n6578), .CK(Clk), .RN(n3945), .QN(n1241)
         );
  DFFR_X1 \pc_lut_reg[30][31]  ( .D(n6577), .CK(Clk), .RN(n3945), .Q(
        \pc_lut[30][31] ), .QN(n1239) );
  DFFR_X1 \pc_lut_reg[30][29]  ( .D(n6576), .CK(Clk), .RN(n3945), .Q(
        \pc_lut[30][29] ), .QN(n1238) );
  DFFR_X1 \pc_lut_reg[30][27]  ( .D(n6575), .CK(Clk), .RN(n3945), .Q(
        \pc_lut[30][27] ), .QN(n1237) );
  DFFR_X1 \pc_lut_reg[30][25]  ( .D(n6574), .CK(Clk), .RN(n3945), .Q(
        \pc_lut[30][25] ), .QN(n1236) );
  DFFR_X1 \pc_lut_reg[30][23]  ( .D(n6573), .CK(Clk), .RN(n3945), .Q(
        \pc_lut[30][23] ), .QN(n1235) );
  DFFR_X1 \pc_lut_reg[30][21]  ( .D(n6572), .CK(Clk), .RN(n3946), .Q(
        \pc_lut[30][21] ), .QN(n1234) );
  DFFR_X1 \pc_lut_reg[30][19]  ( .D(n6571), .CK(Clk), .RN(n3946), .Q(
        \pc_lut[30][19] ), .QN(n1233) );
  DFFR_X1 \pc_lut_reg[30][17]  ( .D(n6570), .CK(Clk), .RN(n3946), .Q(
        \pc_lut[30][17] ), .QN(n1232) );
  DFFR_X1 \pc_lut_reg[30][15]  ( .D(n6569), .CK(Clk), .RN(n3946), .Q(
        \pc_lut[30][15] ), .QN(n1231) );
  DFFR_X1 \pc_lut_reg[30][13]  ( .D(n6568), .CK(Clk), .RN(n3946), .Q(
        \pc_lut[30][13] ), .QN(n1230) );
  DFFR_X1 \pc_lut_reg[30][11]  ( .D(n6567), .CK(Clk), .RN(n3946), .Q(
        \pc_lut[30][11] ), .QN(n1229) );
  DFFR_X1 \pc_lut_reg[30][9]  ( .D(n6566), .CK(Clk), .RN(n3946), .Q(
        \pc_lut[30][9] ), .QN(n1228) );
  DFFR_X1 \pc_lut_reg[30][7]  ( .D(n6565), .CK(Clk), .RN(n3946), .Q(
        \pc_lut[30][7] ), .QN(n1227) );
  DFFR_X1 \pc_lut_reg[30][5]  ( .D(n6564), .CK(Clk), .RN(n3861), .Q(
        \pc_lut[30][5] ), .QN(n1226) );
  DFFR_X1 \pc_lut_reg[30][3]  ( .D(n6563), .CK(Clk), .RN(n3946), .Q(
        \pc_lut[30][3] ) );
  DFFR_X1 \pc_lut_reg[30][1]  ( .D(n6562), .CK(Clk), .RN(n3946), .Q(
        \pc_lut[30][1] ) );
  DFFR_X1 \pc_lut_reg[30][2]  ( .D(n6560), .CK(Clk), .RN(n3946), .Q(
        \pc_lut[30][2] ) );
  DFFR_X1 \pc_lut_reg[30][4]  ( .D(n6559), .CK(Clk), .RN(n3946), .Q(
        \pc_lut[30][4] ) );
  DFFR_X1 \pc_lut_reg[30][6]  ( .D(n6558), .CK(Clk), .RN(n3946), .Q(
        \pc_lut[30][6] ), .QN(n1221) );
  DFFR_X1 \pc_lut_reg[30][8]  ( .D(n6557), .CK(Clk), .RN(n3946), .Q(
        \pc_lut[30][8] ), .QN(n1220) );
  DFFR_X1 \pc_lut_reg[30][10]  ( .D(n6556), .CK(Clk), .RN(n3946), .Q(
        \pc_lut[30][10] ), .QN(n1219) );
  DFFR_X1 \pc_lut_reg[30][12]  ( .D(n6555), .CK(Clk), .RN(n3947), .Q(
        \pc_lut[30][12] ), .QN(n1218) );
  DFFR_X1 \pc_lut_reg[30][14]  ( .D(n6554), .CK(Clk), .RN(n3947), .Q(
        \pc_lut[30][14] ), .QN(n1217) );
  DFFR_X1 \pc_lut_reg[30][16]  ( .D(n6553), .CK(Clk), .RN(n3947), .Q(
        \pc_lut[30][16] ), .QN(n1216) );
  DFFR_X1 \pc_lut_reg[30][18]  ( .D(n6552), .CK(Clk), .RN(n3880), .Q(
        \pc_lut[30][18] ), .QN(n1215) );
  DFFR_X1 \pc_lut_reg[30][20]  ( .D(n6551), .CK(Clk), .RN(n3947), .Q(
        \pc_lut[30][20] ), .QN(n1214) );
  DFFR_X1 \pc_lut_reg[30][22]  ( .D(n6550), .CK(Clk), .RN(n3947), .Q(
        \pc_lut[30][22] ), .QN(n1213) );
  DFFR_X1 \pc_lut_reg[30][24]  ( .D(n6549), .CK(Clk), .RN(n3947), .Q(
        \pc_lut[30][24] ), .QN(n1212) );
  DFFR_X1 \pc_lut_reg[30][26]  ( .D(n6548), .CK(Clk), .RN(n3947), .Q(
        \pc_lut[30][26] ), .QN(n1211) );
  DFFR_X1 \pc_lut_reg[30][28]  ( .D(n6547), .CK(Clk), .RN(n3947), .Q(
        \pc_lut[30][28] ), .QN(n1210) );
  DFFR_X1 \pc_lut_reg[30][30]  ( .D(n6546), .CK(Clk), .RN(n3947), .Q(
        \pc_lut[30][30] ), .QN(n1208) );
  DFFR_X1 \pc_lut_reg[31][31]  ( .D(n6545), .CK(Clk), .RN(n3947), .Q(
        \pc_lut[31][31] ), .QN(n1204) );
  DFFR_X1 \pc_lut_reg[31][29]  ( .D(n6544), .CK(Clk), .RN(n3841), .Q(
        \pc_lut[31][29] ), .QN(n1202) );
  DFFR_X1 \pc_lut_reg[31][27]  ( .D(n6543), .CK(Clk), .RN(n3841), .Q(
        \pc_lut[31][27] ), .QN(n1200) );
  DFFR_X1 \pc_lut_reg[31][25]  ( .D(n6542), .CK(Clk), .RN(n3894), .Q(
        \pc_lut[31][25] ), .QN(n1198) );
  DFFR_X1 \pc_lut_reg[31][23]  ( .D(n6541), .CK(Clk), .RN(n3841), .Q(
        \pc_lut[31][23] ), .QN(n1196) );
  DFFR_X1 \pc_lut_reg[31][21]  ( .D(n6540), .CK(Clk), .RN(n3841), .Q(
        \pc_lut[31][21] ), .QN(n1194) );
  DFFR_X1 \pc_lut_reg[31][19]  ( .D(n6539), .CK(Clk), .RN(n3841), .Q(
        \pc_lut[31][19] ), .QN(n1192) );
  DFFR_X1 \pc_lut_reg[31][17]  ( .D(n6538), .CK(Clk), .RN(n3841), .Q(
        \pc_lut[31][17] ), .QN(n1190) );
  DFFR_X1 \pc_lut_reg[31][15]  ( .D(n6537), .CK(Clk), .RN(n3842), .Q(
        \pc_lut[31][15] ), .QN(n1188) );
  DFFR_X1 \pc_lut_reg[31][13]  ( .D(n6536), .CK(Clk), .RN(n3842), .Q(
        \pc_lut[31][13] ), .QN(n1186) );
  DFFR_X1 \pc_lut_reg[31][11]  ( .D(n6535), .CK(Clk), .RN(n3842), .Q(
        \pc_lut[31][11] ), .QN(n1184) );
  DFFR_X1 \pc_lut_reg[31][9]  ( .D(n6534), .CK(Clk), .RN(n3842), .Q(
        \pc_lut[31][9] ), .QN(n1182) );
  DFFR_X1 \pc_lut_reg[31][7]  ( .D(n6533), .CK(Clk), .RN(n3842), .Q(
        \pc_lut[31][7] ), .QN(n1180) );
  DFFR_X1 \pc_lut_reg[31][5]  ( .D(n6532), .CK(Clk), .RN(n3861), .Q(
        \pc_lut[31][5] ), .QN(n1178) );
  DFFR_X1 \pc_lut_reg[31][6]  ( .D(n6526), .CK(Clk), .RN(n3842), .Q(
        \pc_lut[31][6] ), .QN(n1171) );
  DFFR_X1 \pc_lut_reg[31][8]  ( .D(n6525), .CK(Clk), .RN(n3842), .Q(
        \pc_lut[31][8] ), .QN(n1169) );
  DFFR_X1 \pc_lut_reg[31][10]  ( .D(n6524), .CK(Clk), .RN(n3842), .Q(
        \pc_lut[31][10] ), .QN(n1167) );
  DFFR_X1 \pc_lut_reg[31][12]  ( .D(n6523), .CK(Clk), .RN(n3842), .Q(
        \pc_lut[31][12] ), .QN(n1165) );
  DFFR_X1 \pc_lut_reg[31][14]  ( .D(n6522), .CK(Clk), .RN(n3842), .Q(
        \pc_lut[31][14] ), .QN(n1163) );
  DFFR_X1 \pc_lut_reg[31][16]  ( .D(n6521), .CK(Clk), .RN(n3843), .Q(
        \pc_lut[31][16] ), .QN(n1161) );
  DFFR_X1 \pc_lut_reg[31][18]  ( .D(n6520), .CK(Clk), .RN(n3880), .Q(
        \pc_lut[31][18] ), .QN(n1159) );
  DFFR_X1 \pc_lut_reg[31][20]  ( .D(n6519), .CK(Clk), .RN(n3843), .Q(
        \pc_lut[31][20] ), .QN(n1157) );
  DFFR_X1 \pc_lut_reg[31][22]  ( .D(n6518), .CK(Clk), .RN(n3843), .Q(
        \pc_lut[31][22] ), .QN(n1155) );
  DFFR_X1 \pc_lut_reg[31][24]  ( .D(n6517), .CK(Clk), .RN(n3843), .Q(
        \pc_lut[31][24] ), .QN(n1153) );
  DFFR_X1 \pc_lut_reg[31][26]  ( .D(n6516), .CK(Clk), .RN(n3843), .Q(
        \pc_lut[31][26] ), .QN(n1151) );
  DFFR_X1 \pc_lut_reg[31][28]  ( .D(n6515), .CK(Clk), .RN(n3843), .Q(
        \pc_lut[31][28] ), .QN(n1149) );
  DFFR_X1 \pc_lut_reg[31][30]  ( .D(n6514), .CK(Clk), .RN(n3844), .Q(
        \pc_lut[31][30] ), .QN(n1146) );
  DLH_X1 OUTT_NTs_reg ( .G(Enable), .D(N220), .Q(OUTT_NT) );
  DFFR_X1 \pc_target_reg[0][31]  ( .D(n6513), .CK(Clk), .RN(n3864), .QN(n1142)
         );
  DFFR_X1 \pc_target_reg[0][29]  ( .D(n6512), .CK(Clk), .RN(n3843), .QN(n1141)
         );
  DFFR_X1 \pc_target_reg[0][27]  ( .D(n6511), .CK(Clk), .RN(n3843), .QN(n1140)
         );
  DFFR_X1 \pc_target_reg[0][25]  ( .D(n6510), .CK(Clk), .RN(n3843), .QN(n1139)
         );
  DFFR_X1 \pc_target_reg[0][23]  ( .D(n6509), .CK(Clk), .RN(n3843), .QN(n1138)
         );
  DFFR_X1 \pc_target_reg[0][21]  ( .D(n6508), .CK(Clk), .RN(n3843), .QN(n1137)
         );
  DFFR_X1 \pc_target_reg[0][19]  ( .D(n6507), .CK(Clk), .RN(n3843), .QN(n1136)
         );
  DFFR_X1 \pc_target_reg[0][17]  ( .D(n6506), .CK(Clk), .RN(n3843), .QN(n1135)
         );
  DFFR_X1 \pc_target_reg[0][15]  ( .D(n6505), .CK(Clk), .RN(n3843), .QN(n1134)
         );
  DFFR_X1 \pc_target_reg[0][13]  ( .D(n6504), .CK(Clk), .RN(n3844), .QN(n1133)
         );
  DFFR_X1 \pc_target_reg[0][11]  ( .D(n6503), .CK(Clk), .RN(n3844), .QN(n1132)
         );
  DFFR_X1 \pc_target_reg[0][9]  ( .D(n6502), .CK(Clk), .RN(n3844), .QN(n1131)
         );
  DFFR_X1 \pc_target_reg[0][7]  ( .D(n6501), .CK(Clk), .RN(n3844), .QN(n1130)
         );
  DFFR_X1 \pc_target_reg[0][5]  ( .D(n6500), .CK(Clk), .RN(n3844), .QN(n1129)
         );
  DFFR_X1 \pc_target_reg[0][3]  ( .D(n6499), .CK(Clk), .RN(n3844), .QN(n1128)
         );
  DFFR_X1 \pc_target_reg[0][1]  ( .D(n6498), .CK(Clk), .RN(n3844), .QN(n1127)
         );
  DFFR_X1 \pc_target_reg[0][0]  ( .D(n6497), .CK(Clk), .RN(n3844), .QN(n1126)
         );
  DFFR_X1 \pc_target_reg[0][2]  ( .D(n6496), .CK(Clk), .RN(n3844), .QN(n1125)
         );
  DFFR_X1 \pc_target_reg[0][4]  ( .D(n6495), .CK(Clk), .RN(n3844), .QN(n1124)
         );
  DFFR_X1 \pc_target_reg[0][6]  ( .D(n6494), .CK(Clk), .RN(n3844), .QN(n1123)
         );
  DFFR_X1 \pc_target_reg[0][8]  ( .D(n6493), .CK(Clk), .RN(n3844), .QN(n1122)
         );
  DFFR_X1 \pc_target_reg[0][10]  ( .D(n6492), .CK(Clk), .RN(n3844), .QN(n1121)
         );
  DFFR_X1 \pc_target_reg[0][12]  ( .D(n6491), .CK(Clk), .RN(n3844), .QN(n1120)
         );
  DFFR_X1 \pc_target_reg[0][14]  ( .D(n6490), .CK(Clk), .RN(n3845), .QN(n1119)
         );
  DFFR_X1 \pc_target_reg[0][16]  ( .D(n6489), .CK(Clk), .RN(n3845), .QN(n1118)
         );
  DFFR_X1 \pc_target_reg[0][18]  ( .D(n6488), .CK(Clk), .RN(n3845), .QN(n1117)
         );
  DFFR_X1 \pc_target_reg[0][20]  ( .D(n6487), .CK(Clk), .RN(n3845), .QN(n1116)
         );
  DFFR_X1 \pc_target_reg[0][22]  ( .D(n6486), .CK(Clk), .RN(n3845), .QN(n1115)
         );
  DFFR_X1 \pc_target_reg[0][24]  ( .D(n6485), .CK(Clk), .RN(n3845), .QN(n1114)
         );
  DFFR_X1 \pc_target_reg[0][26]  ( .D(n6484), .CK(Clk), .RN(n3845), .QN(n1113)
         );
  DFFR_X1 \pc_target_reg[0][28]  ( .D(n6483), .CK(Clk), .RN(n3845), .QN(n1112)
         );
  DFFR_X1 \pc_target_reg[1][31]  ( .D(n6481), .CK(Clk), .RN(n3865), .QN(n1108)
         );
  DFFR_X1 \pc_target_reg[1][29]  ( .D(n6480), .CK(Clk), .RN(n3845), .QN(n1107)
         );
  DFFR_X1 \pc_target_reg[1][27]  ( .D(n6479), .CK(Clk), .RN(n3845), .QN(n1106)
         );
  DFFR_X1 \pc_target_reg[1][25]  ( .D(n6478), .CK(Clk), .RN(n3845), .QN(n1105)
         );
  DFFR_X1 \pc_target_reg[1][23]  ( .D(n6477), .CK(Clk), .RN(n3845), .QN(n1104)
         );
  DFFR_X1 \pc_target_reg[1][21]  ( .D(n6476), .CK(Clk), .RN(n3845), .QN(n1103)
         );
  DFFR_X1 \pc_target_reg[1][19]  ( .D(n6475), .CK(Clk), .RN(n3845), .QN(n1102)
         );
  DFFR_X1 \pc_target_reg[1][17]  ( .D(n6474), .CK(Clk), .RN(n3845), .QN(n1101)
         );
  DFFR_X1 \pc_target_reg[1][15]  ( .D(n6473), .CK(Clk), .RN(n3846), .QN(n1100)
         );
  DFFR_X1 \pc_target_reg[1][13]  ( .D(n6472), .CK(Clk), .RN(n3846), .QN(n1099)
         );
  DFFR_X1 \pc_target_reg[1][11]  ( .D(n6471), .CK(Clk), .RN(n3846), .QN(n1098)
         );
  DFFR_X1 \pc_target_reg[1][9]  ( .D(n6470), .CK(Clk), .RN(n3846), .QN(n1097)
         );
  DFFR_X1 \pc_target_reg[1][7]  ( .D(n6469), .CK(Clk), .RN(n3846), .QN(n1096)
         );
  DFFR_X1 \pc_target_reg[1][5]  ( .D(n6468), .CK(Clk), .RN(n3846), .QN(n1095)
         );
  DFFR_X1 \pc_target_reg[1][3]  ( .D(n6467), .CK(Clk), .RN(n3846), .QN(n1094)
         );
  DFFR_X1 \pc_target_reg[1][1]  ( .D(n6466), .CK(Clk), .RN(n3846), .QN(n1093)
         );
  DFFR_X1 \pc_target_reg[1][0]  ( .D(n6465), .CK(Clk), .RN(n3847), .QN(n1092)
         );
  DFFR_X1 \pc_target_reg[1][2]  ( .D(n6464), .CK(Clk), .RN(n3846), .QN(n1091)
         );
  DFFR_X1 \pc_target_reg[1][4]  ( .D(n6463), .CK(Clk), .RN(n3846), .QN(n1090)
         );
  DFFR_X1 \pc_target_reg[1][6]  ( .D(n6462), .CK(Clk), .RN(n3846), .QN(n1089)
         );
  DFFR_X1 \pc_target_reg[1][8]  ( .D(n6461), .CK(Clk), .RN(n3846), .QN(n1088)
         );
  DFFR_X1 \pc_target_reg[1][10]  ( .D(n6460), .CK(Clk), .RN(n3846), .QN(n1087)
         );
  DFFR_X1 \pc_target_reg[1][12]  ( .D(n6459), .CK(Clk), .RN(n3846), .QN(n1086)
         );
  DFFR_X1 \pc_target_reg[1][14]  ( .D(n6458), .CK(Clk), .RN(n3846), .QN(n1085)
         );
  DFFR_X1 \pc_target_reg[1][16]  ( .D(n6457), .CK(Clk), .RN(n3847), .QN(n1084)
         );
  DFFR_X1 \pc_target_reg[1][18]  ( .D(n6456), .CK(Clk), .RN(n3847), .QN(n1083)
         );
  DFFR_X1 \pc_target_reg[1][20]  ( .D(n6455), .CK(Clk), .RN(n3847), .QN(n1082)
         );
  DFFR_X1 \pc_target_reg[1][22]  ( .D(n6454), .CK(Clk), .RN(n3847), .QN(n1081)
         );
  DFFR_X1 \pc_target_reg[1][24]  ( .D(n6453), .CK(Clk), .RN(n3847), .QN(n1080)
         );
  DFFR_X1 \pc_target_reg[1][26]  ( .D(n6452), .CK(Clk), .RN(n3847), .QN(n1079)
         );
  DFFR_X1 \pc_target_reg[1][28]  ( .D(n6451), .CK(Clk), .RN(n3847), .QN(n1078)
         );
  DFFR_X1 \pc_target_reg[3][31]  ( .D(n6417), .CK(Clk), .RN(n3864), .Q(
        \pc_target[3][31] ) );
  DFFR_X1 \pc_target_reg[3][29]  ( .D(n6416), .CK(Clk), .RN(n3847), .Q(
        \pc_target[3][29] ) );
  DFFR_X1 \pc_target_reg[3][27]  ( .D(n6415), .CK(Clk), .RN(n3847), .Q(
        \pc_target[3][27] ) );
  DFFR_X1 \pc_target_reg[3][25]  ( .D(n6414), .CK(Clk), .RN(n3847), .Q(
        \pc_target[3][25] ) );
  DFFR_X1 \pc_target_reg[3][23]  ( .D(n6413), .CK(Clk), .RN(n3847), .Q(
        \pc_target[3][23] ) );
  DFFR_X1 \pc_target_reg[3][21]  ( .D(n6412), .CK(Clk), .RN(n3847), .Q(
        \pc_target[3][21] ) );
  DFFR_X1 \pc_target_reg[3][19]  ( .D(n6411), .CK(Clk), .RN(n3855), .Q(
        \pc_target[3][19] ) );
  DFFR_X1 \pc_target_reg[3][17]  ( .D(n6410), .CK(Clk), .RN(n3937), .Q(
        \pc_target[3][17] ) );
  DFFR_X1 \pc_target_reg[3][15]  ( .D(n6409), .CK(Clk), .RN(n3933), .Q(
        \pc_target[3][15] ) );
  DFFR_X1 \pc_target_reg[3][13]  ( .D(n6408), .CK(Clk), .RN(n3929), .Q(
        \pc_target[3][13] ) );
  DFFR_X1 \pc_target_reg[3][11]  ( .D(n6407), .CK(Clk), .RN(n3929), .Q(
        \pc_target[3][11] ) );
  DFFR_X1 \pc_target_reg[3][7]  ( .D(n6405), .CK(Clk), .RN(n3929), .Q(
        \pc_target[3][7] ) );
  DFFR_X1 \pc_target_reg[3][12]  ( .D(n6395), .CK(Clk), .RN(n3929), .Q(
        \pc_target[3][12] ) );
  DFFR_X1 \pc_target_reg[3][14]  ( .D(n6394), .CK(Clk), .RN(n3929), .Q(
        \pc_target[3][14] ) );
  DFFR_X1 \pc_target_reg[3][16]  ( .D(n6393), .CK(Clk), .RN(n3929), .Q(
        \pc_target[3][16] ) );
  DFFR_X1 \pc_target_reg[3][18]  ( .D(n6392), .CK(Clk), .RN(n3929), .Q(
        \pc_target[3][18] ) );
  DFFR_X1 \pc_target_reg[3][20]  ( .D(n6391), .CK(Clk), .RN(n3929), .Q(
        \pc_target[3][20] ) );
  DFFR_X1 \pc_target_reg[3][22]  ( .D(n6390), .CK(Clk), .RN(n3930), .Q(
        \pc_target[3][22] ) );
  DFFR_X1 \pc_target_reg[3][24]  ( .D(n6389), .CK(Clk), .RN(n3930), .Q(
        \pc_target[3][24] ) );
  DFFR_X1 \pc_target_reg[3][26]  ( .D(n6388), .CK(Clk), .RN(n3930), .Q(
        \pc_target[3][26] ) );
  DFFR_X1 \pc_target_reg[3][28]  ( .D(n6387), .CK(Clk), .RN(n3930), .Q(
        \pc_target[3][28] ) );
  DFFR_X1 \pc_target_reg[3][30]  ( .D(n6386), .CK(Clk), .RN(n3930), .Q(
        \pc_target[3][30] ) );
  DFFR_X1 \pc_target_reg[4][31]  ( .D(n6385), .CK(Clk), .RN(n3864), .QN(n1005)
         );
  DFFR_X1 \pc_target_reg[4][29]  ( .D(n6384), .CK(Clk), .RN(n3929), .QN(n1004)
         );
  DFFR_X1 \pc_target_reg[4][27]  ( .D(n6383), .CK(Clk), .RN(n3929), .QN(n1003)
         );
  DFFR_X1 \pc_target_reg[4][25]  ( .D(n6382), .CK(Clk), .RN(n3929), .QN(n1002)
         );
  DFFR_X1 \pc_target_reg[4][23]  ( .D(n6381), .CK(Clk), .RN(n3929), .QN(n1001)
         );
  DFFR_X1 \pc_target_reg[4][21]  ( .D(n6380), .CK(Clk), .RN(n3930), .QN(n1000)
         );
  DFFR_X1 \pc_target_reg[4][19]  ( .D(n6379), .CK(Clk), .RN(n3930), .QN(n999)
         );
  DFFR_X1 \pc_target_reg[4][17]  ( .D(n6378), .CK(Clk), .RN(n3930), .QN(n998)
         );
  DFFR_X1 \pc_target_reg[4][15]  ( .D(n6377), .CK(Clk), .RN(n3930), .QN(n997)
         );
  DFFR_X1 \pc_target_reg[4][13]  ( .D(n6376), .CK(Clk), .RN(n3930), .QN(n996)
         );
  DFFR_X1 \pc_target_reg[4][11]  ( .D(n6375), .CK(Clk), .RN(n3930), .QN(n995)
         );
  DFFR_X1 \pc_target_reg[4][9]  ( .D(n6374), .CK(Clk), .RN(n3930), .QN(n994)
         );
  DFFR_X1 \pc_target_reg[4][7]  ( .D(n6373), .CK(Clk), .RN(n3930), .QN(n993)
         );
  DFFR_X1 \pc_target_reg[4][3]  ( .D(n6371), .CK(Clk), .RN(n3930), .QN(n991)
         );
  DFFR_X1 \pc_target_reg[4][1]  ( .D(n6370), .CK(Clk), .RN(n3930), .QN(n990)
         );
  DFFR_X1 \pc_target_reg[4][0]  ( .D(n6369), .CK(Clk), .RN(n3931), .QN(n989)
         );
  DFFR_X1 \pc_target_reg[4][2]  ( .D(n6368), .CK(Clk), .RN(n3931), .QN(n988)
         );
  DFFR_X1 \pc_target_reg[4][6]  ( .D(n6366), .CK(Clk), .RN(n3931), .QN(n986)
         );
  DFFR_X1 \pc_target_reg[4][8]  ( .D(n6365), .CK(Clk), .RN(n3931), .QN(n985)
         );
  DFFR_X1 \pc_target_reg[4][10]  ( .D(n6364), .CK(Clk), .RN(n3931), .QN(n984)
         );
  DFFR_X1 \pc_target_reg[4][12]  ( .D(n6363), .CK(Clk), .RN(n3931), .QN(n983)
         );
  DFFR_X1 \pc_target_reg[4][14]  ( .D(n6362), .CK(Clk), .RN(n3931), .QN(n982)
         );
  DFFR_X1 \pc_target_reg[4][16]  ( .D(n6361), .CK(Clk), .RN(n3931), .QN(n981)
         );
  DFFR_X1 \pc_target_reg[4][18]  ( .D(n6360), .CK(Clk), .RN(n3931), .QN(n980)
         );
  DFFR_X1 \pc_target_reg[4][20]  ( .D(n6359), .CK(Clk), .RN(n3931), .QN(n979)
         );
  DFFR_X1 \pc_target_reg[4][22]  ( .D(n6358), .CK(Clk), .RN(n3931), .QN(n978)
         );
  DFFR_X1 \pc_target_reg[4][24]  ( .D(n6357), .CK(Clk), .RN(n3931), .QN(n977)
         );
  DFFR_X1 \pc_target_reg[4][26]  ( .D(n6356), .CK(Clk), .RN(n3932), .QN(n976)
         );
  DFFR_X1 \pc_target_reg[4][28]  ( .D(n6355), .CK(Clk), .RN(n3932), .QN(n975)
         );
  DFFR_X1 \pc_target_reg[5][31]  ( .D(n6353), .CK(Clk), .RN(n3864), .QN(n971)
         );
  DFFR_X1 \pc_target_reg[5][29]  ( .D(n6352), .CK(Clk), .RN(n3931), .QN(n970)
         );
  DFFR_X1 \pc_target_reg[5][27]  ( .D(n6351), .CK(Clk), .RN(n3931), .QN(n969)
         );
  DFFR_X1 \pc_target_reg[5][25]  ( .D(n6350), .CK(Clk), .RN(n3931), .QN(n968)
         );
  DFFR_X1 \pc_target_reg[5][23]  ( .D(n6349), .CK(Clk), .RN(n3932), .QN(n967)
         );
  DFFR_X1 \pc_target_reg[5][21]  ( .D(n6348), .CK(Clk), .RN(n3932), .QN(n966)
         );
  DFFR_X1 \pc_target_reg[5][19]  ( .D(n6347), .CK(Clk), .RN(n3932), .QN(n965)
         );
  DFFR_X1 \pc_target_reg[5][17]  ( .D(n6346), .CK(Clk), .RN(n3932), .QN(n964)
         );
  DFFR_X1 \pc_target_reg[5][15]  ( .D(n6345), .CK(Clk), .RN(n3932), .QN(n963)
         );
  DFFR_X1 \pc_target_reg[5][13]  ( .D(n6344), .CK(Clk), .RN(n3932), .QN(n962)
         );
  DFFR_X1 \pc_target_reg[5][11]  ( .D(n6343), .CK(Clk), .RN(n3932), .QN(n961)
         );
  DFFR_X1 \pc_target_reg[5][9]  ( .D(n6342), .CK(Clk), .RN(n3932), .QN(n960)
         );
  DFFR_X1 \pc_target_reg[5][7]  ( .D(n6341), .CK(Clk), .RN(n3932), .QN(n959)
         );
  DFFR_X1 \pc_target_reg[5][5]  ( .D(n6340), .CK(Clk), .RN(n3932), .QN(n958)
         );
  DFFR_X1 \pc_target_reg[5][3]  ( .D(n6339), .CK(Clk), .RN(n3932), .QN(n957)
         );
  DFFR_X1 \pc_target_reg[5][1]  ( .D(n6338), .CK(Clk), .RN(n3932), .QN(n956)
         );
  DFFR_X1 \pc_target_reg[5][0]  ( .D(n6337), .CK(Clk), .RN(n3933), .QN(n955)
         );
  DFFR_X1 \pc_target_reg[5][2]  ( .D(n6336), .CK(Clk), .RN(n3932), .QN(n954)
         );
  DFFR_X1 \pc_target_reg[5][4]  ( .D(n6335), .CK(Clk), .RN(n3933), .QN(n953)
         );
  DFFR_X1 \pc_target_reg[5][6]  ( .D(n6334), .CK(Clk), .RN(n3933), .QN(n952)
         );
  DFFR_X1 \pc_target_reg[5][8]  ( .D(n6333), .CK(Clk), .RN(n3933), .QN(n951)
         );
  DFFR_X1 \pc_target_reg[5][10]  ( .D(n6332), .CK(Clk), .RN(n3933), .QN(n950)
         );
  DFFR_X1 \pc_target_reg[5][12]  ( .D(n6331), .CK(Clk), .RN(n3933), .QN(n949)
         );
  DFFR_X1 \pc_target_reg[5][14]  ( .D(n6330), .CK(Clk), .RN(n3933), .QN(n948)
         );
  DFFR_X1 \pc_target_reg[5][16]  ( .D(n6329), .CK(Clk), .RN(n3933), .QN(n947)
         );
  DFFR_X1 \pc_target_reg[5][18]  ( .D(n6328), .CK(Clk), .RN(n3933), .QN(n946)
         );
  DFFR_X1 \pc_target_reg[5][20]  ( .D(n6327), .CK(Clk), .RN(n3933), .QN(n945)
         );
  DFFR_X1 \pc_target_reg[5][22]  ( .D(n6326), .CK(Clk), .RN(n3933), .QN(n944)
         );
  DFFR_X1 \pc_target_reg[5][24]  ( .D(n6325), .CK(Clk), .RN(n3933), .QN(n943)
         );
  DFFR_X1 \pc_target_reg[5][26]  ( .D(n6324), .CK(Clk), .RN(n3933), .QN(n942)
         );
  DFFR_X1 \pc_target_reg[5][28]  ( .D(n6323), .CK(Clk), .RN(n3933), .QN(n941)
         );
  DFFR_X1 \pc_target_reg[7][5]  ( .D(n6276), .CK(Clk), .RN(n3830), .Q(
        \pc_target[7][5] ) );
  DFFR_X1 \pc_target_reg[7][3]  ( .D(n6275), .CK(Clk), .RN(n3830), .Q(
        \pc_target[7][3] ) );
  DFFR_X1 \pc_target_reg[7][1]  ( .D(n6274), .CK(Clk), .RN(n3830), .Q(
        \pc_target[7][1] ) );
  DFFR_X1 \pc_target_reg[7][0]  ( .D(n6273), .CK(Clk), .RN(n3831), .Q(
        \pc_target[7][0] ) );
  DFFR_X1 \pc_target_reg[7][2]  ( .D(n6272), .CK(Clk), .RN(n3830), .Q(
        \pc_target[7][2] ) );
  DFFR_X1 \pc_target_reg[7][4]  ( .D(n6271), .CK(Clk), .RN(n3830), .Q(
        \pc_target[7][4] ) );
  DFFR_X1 \pc_target_reg[7][6]  ( .D(n6270), .CK(Clk), .RN(n3830), .Q(
        \pc_target[7][6] ) );
  DFFR_X1 \pc_target_reg[8][31]  ( .D(n6257), .CK(Clk), .RN(n3865), .QN(n868)
         );
  DFFR_X1 \pc_target_reg[8][29]  ( .D(n6256), .CK(Clk), .RN(n3831), .QN(n867)
         );
  DFFR_X1 \pc_target_reg[8][27]  ( .D(n6255), .CK(Clk), .RN(n3831), .QN(n866)
         );
  DFFR_X1 \pc_target_reg[8][25]  ( .D(n6254), .CK(Clk), .RN(n3832), .QN(n865)
         );
  DFFR_X1 \pc_target_reg[8][23]  ( .D(n6253), .CK(Clk), .RN(n3832), .QN(n864)
         );
  DFFR_X1 \pc_target_reg[8][21]  ( .D(n6252), .CK(Clk), .RN(n3832), .QN(n863)
         );
  DFFR_X1 \pc_target_reg[8][19]  ( .D(n6251), .CK(Clk), .RN(n3832), .QN(n862)
         );
  DFFR_X1 \pc_target_reg[8][17]  ( .D(n6250), .CK(Clk), .RN(n3832), .QN(n861)
         );
  DFFR_X1 \pc_target_reg[8][15]  ( .D(n6249), .CK(Clk), .RN(n3832), .QN(n860)
         );
  DFFR_X1 \pc_target_reg[8][13]  ( .D(n6248), .CK(Clk), .RN(n3851), .QN(n859)
         );
  DFFR_X1 \pc_target_reg[8][11]  ( .D(n6247), .CK(Clk), .RN(n3847), .QN(n858)
         );
  DFFR_X1 \pc_target_reg[8][9]  ( .D(n6246), .CK(Clk), .RN(n3847), .QN(n857)
         );
  DFFR_X1 \pc_target_reg[8][7]  ( .D(n6245), .CK(Clk), .RN(n3848), .QN(n856)
         );
  DFFR_X1 \pc_target_reg[8][5]  ( .D(n6244), .CK(Clk), .RN(n3848), .QN(n855)
         );
  DFFR_X1 \pc_target_reg[8][3]  ( .D(n6243), .CK(Clk), .RN(n3848), .QN(n854)
         );
  DFFR_X1 \pc_target_reg[8][1]  ( .D(n6242), .CK(Clk), .RN(n3848), .QN(n853)
         );
  DFFR_X1 \pc_target_reg[8][0]  ( .D(n6241), .CK(Clk), .RN(n3848), .QN(n852)
         );
  DFFR_X1 \pc_target_reg[8][2]  ( .D(n6240), .CK(Clk), .RN(n3848), .QN(n851)
         );
  DFFR_X1 \pc_target_reg[8][4]  ( .D(n6239), .CK(Clk), .RN(n3848), .QN(n850)
         );
  DFFR_X1 \pc_target_reg[8][6]  ( .D(n6238), .CK(Clk), .RN(n3848), .QN(n849)
         );
  DFFR_X1 \pc_target_reg[8][8]  ( .D(n6237), .CK(Clk), .RN(n3848), .QN(n848)
         );
  DFFR_X1 \pc_target_reg[8][10]  ( .D(n6236), .CK(Clk), .RN(n3848), .QN(n847)
         );
  DFFR_X1 \pc_target_reg[8][12]  ( .D(n6235), .CK(Clk), .RN(n3848), .QN(n846)
         );
  DFFR_X1 \pc_target_reg[8][14]  ( .D(n6234), .CK(Clk), .RN(n3848), .QN(n845)
         );
  DFFR_X1 \pc_target_reg[8][16]  ( .D(n6233), .CK(Clk), .RN(n3848), .QN(n844)
         );
  DFFR_X1 \pc_target_reg[8][18]  ( .D(n6232), .CK(Clk), .RN(n3848), .QN(n843)
         );
  DFFR_X1 \pc_target_reg[8][20]  ( .D(n6231), .CK(Clk), .RN(n3848), .QN(n842)
         );
  DFFR_X1 \pc_target_reg[8][22]  ( .D(n6230), .CK(Clk), .RN(n3849), .QN(n841)
         );
  DFFR_X1 \pc_target_reg[8][24]  ( .D(n6229), .CK(Clk), .RN(n3849), .QN(n840)
         );
  DFFR_X1 \pc_target_reg[8][26]  ( .D(n6228), .CK(Clk), .RN(n3849), .QN(n839)
         );
  DFFR_X1 \pc_target_reg[8][28]  ( .D(n6227), .CK(Clk), .RN(n3849), .QN(n838)
         );
  DFFR_X1 \pc_target_reg[9][31]  ( .D(n6225), .CK(Clk), .RN(n3865), .QN(n834)
         );
  DFFR_X1 \pc_target_reg[9][29]  ( .D(n6224), .CK(Clk), .RN(n3849), .QN(n833)
         );
  DFFR_X1 \pc_target_reg[9][27]  ( .D(n6223), .CK(Clk), .RN(n3849), .QN(n832)
         );
  DFFR_X1 \pc_target_reg[9][25]  ( .D(n6222), .CK(Clk), .RN(n3849), .QN(n831)
         );
  DFFR_X1 \pc_target_reg[9][23]  ( .D(n6221), .CK(Clk), .RN(n3849), .QN(n830)
         );
  DFFR_X1 \pc_target_reg[9][21]  ( .D(n6220), .CK(Clk), .RN(n3849), .QN(n829)
         );
  DFFR_X1 \pc_target_reg[9][19]  ( .D(n6219), .CK(Clk), .RN(n3849), .QN(n828)
         );
  DFFR_X1 \pc_target_reg[9][17]  ( .D(n6218), .CK(Clk), .RN(n3849), .QN(n827)
         );
  DFFR_X1 \pc_target_reg[9][15]  ( .D(n6217), .CK(Clk), .RN(n3849), .QN(n826)
         );
  DFFR_X1 \pc_target_reg[9][13]  ( .D(n6216), .CK(Clk), .RN(n3849), .QN(n825)
         );
  DFFR_X1 \pc_target_reg[9][11]  ( .D(n6215), .CK(Clk), .RN(n3849), .QN(n824)
         );
  DFFR_X1 \pc_target_reg[9][9]  ( .D(n6214), .CK(Clk), .RN(n3849), .QN(n823)
         );
  DFFR_X1 \pc_target_reg[9][7]  ( .D(n6213), .CK(Clk), .RN(n3850), .QN(n822)
         );
  DFFR_X1 \pc_target_reg[9][3]  ( .D(n6211), .CK(Clk), .RN(n3850), .QN(n820)
         );
  DFFR_X1 \pc_target_reg[9][1]  ( .D(n6210), .CK(Clk), .RN(n3850), .QN(n819)
         );
  DFFR_X1 \pc_target_reg[9][0]  ( .D(n6209), .CK(Clk), .RN(n3850), .QN(n818)
         );
  DFFR_X1 \pc_target_reg[9][2]  ( .D(n6208), .CK(Clk), .RN(n3850), .QN(n817)
         );
  DFFR_X1 \pc_target_reg[9][6]  ( .D(n6206), .CK(Clk), .RN(n3850), .QN(n815)
         );
  DFFR_X1 \pc_target_reg[9][8]  ( .D(n6205), .CK(Clk), .RN(n3850), .QN(n814)
         );
  DFFR_X1 \pc_target_reg[9][10]  ( .D(n6204), .CK(Clk), .RN(n3850), .QN(n813)
         );
  DFFR_X1 \pc_target_reg[9][12]  ( .D(n6203), .CK(Clk), .RN(n3850), .QN(n812)
         );
  DFFR_X1 \pc_target_reg[9][14]  ( .D(n6202), .CK(Clk), .RN(n3850), .QN(n811)
         );
  DFFR_X1 \pc_target_reg[9][16]  ( .D(n6201), .CK(Clk), .RN(n3850), .QN(n810)
         );
  DFFR_X1 \pc_target_reg[9][18]  ( .D(n6200), .CK(Clk), .RN(n3850), .QN(n809)
         );
  DFFR_X1 \pc_target_reg[9][20]  ( .D(n6199), .CK(Clk), .RN(n3850), .QN(n808)
         );
  DFFR_X1 \pc_target_reg[9][22]  ( .D(n6198), .CK(Clk), .RN(n3850), .QN(n807)
         );
  DFFR_X1 \pc_target_reg[9][24]  ( .D(n6197), .CK(Clk), .RN(n3850), .QN(n806)
         );
  DFFR_X1 \pc_target_reg[9][26]  ( .D(n6196), .CK(Clk), .RN(n3851), .QN(n805)
         );
  DFFR_X1 \pc_target_reg[9][28]  ( .D(n6195), .CK(Clk), .RN(n3851), .QN(n804)
         );
  DFFR_X1 \pc_target_reg[10][31]  ( .D(n6193), .CK(Clk), .RN(n3864), .Q(
        \pc_target[10][31] ) );
  DFFR_X1 \pc_target_reg[10][29]  ( .D(n6192), .CK(Clk), .RN(n3851), .Q(
        \pc_target[10][29] ) );
  DFFR_X1 \pc_target_reg[10][27]  ( .D(n6191), .CK(Clk), .RN(n3851), .Q(
        \pc_target[10][27] ) );
  DFFR_X1 \pc_target_reg[10][25]  ( .D(n6190), .CK(Clk), .RN(n3851), .Q(
        \pc_target[10][25] ) );
  DFFR_X1 \pc_target_reg[10][23]  ( .D(n6189), .CK(Clk), .RN(n3851), .Q(
        \pc_target[10][23] ) );
  DFFR_X1 \pc_target_reg[10][21]  ( .D(n6188), .CK(Clk), .RN(n3851), .Q(
        \pc_target[10][21] ) );
  DFFR_X1 \pc_target_reg[10][19]  ( .D(n6187), .CK(Clk), .RN(n3851), .Q(
        \pc_target[10][19] ) );
  DFFR_X1 \pc_target_reg[10][17]  ( .D(n6186), .CK(Clk), .RN(n3851), .Q(
        \pc_target[10][17] ) );
  DFFR_X1 \pc_target_reg[10][15]  ( .D(n6185), .CK(Clk), .RN(n3851), .Q(
        \pc_target[10][15] ) );
  DFFR_X1 \pc_target_reg[10][13]  ( .D(n6184), .CK(Clk), .RN(n3851), .Q(
        \pc_target[10][13] ) );
  DFFR_X1 \pc_target_reg[10][11]  ( .D(n6183), .CK(Clk), .RN(n3851), .Q(
        \pc_target[10][11] ) );
  DFFR_X1 \pc_target_reg[10][7]  ( .D(n6181), .CK(Clk), .RN(n3851), .Q(
        \pc_target[10][7] ) );
  DFFR_X1 \pc_target_reg[10][5]  ( .D(n6180), .CK(Clk), .RN(n3851), .Q(
        \pc_target[10][5] ) );
  DFFR_X1 \pc_target_reg[10][1]  ( .D(n6178), .CK(Clk), .RN(n3852), .Q(
        \pc_target[10][1] ) );
  DFFR_X1 \pc_target_reg[10][0]  ( .D(n6177), .CK(Clk), .RN(n3852), .Q(
        \pc_target[10][0] ) );
  DFFR_X1 \pc_target_reg[10][2]  ( .D(n6176), .CK(Clk), .RN(n3852), .Q(
        \pc_target[10][2] ) );
  DFFR_X1 \pc_target_reg[10][4]  ( .D(n6175), .CK(Clk), .RN(n3852), .Q(
        \pc_target[10][4] ) );
  DFFR_X1 \pc_target_reg[10][6]  ( .D(n6174), .CK(Clk), .RN(n3852), .Q(
        \pc_target[10][6] ) );
  DFFR_X1 \pc_target_reg[10][12]  ( .D(n6171), .CK(Clk), .RN(n3852), .Q(
        \pc_target[10][12] ) );
  DFFR_X1 \pc_target_reg[10][14]  ( .D(n6170), .CK(Clk), .RN(n3852), .Q(
        \pc_target[10][14] ) );
  DFFR_X1 \pc_target_reg[10][16]  ( .D(n6169), .CK(Clk), .RN(n3852), .Q(
        \pc_target[10][16] ) );
  DFFR_X1 \pc_target_reg[10][18]  ( .D(n6168), .CK(Clk), .RN(n3852), .Q(
        \pc_target[10][18] ) );
  DFFR_X1 \pc_target_reg[10][20]  ( .D(n6167), .CK(Clk), .RN(n3852), .Q(
        \pc_target[10][20] ) );
  DFFR_X1 \pc_target_reg[10][22]  ( .D(n6166), .CK(Clk), .RN(n3852), .Q(
        \pc_target[10][22] ) );
  DFFR_X1 \pc_target_reg[10][24]  ( .D(n6165), .CK(Clk), .RN(n3853), .Q(
        \pc_target[10][24] ) );
  DFFR_X1 \pc_target_reg[10][26]  ( .D(n6164), .CK(Clk), .RN(n3853), .Q(
        \pc_target[10][26] ) );
  DFFR_X1 \pc_target_reg[10][28]  ( .D(n6163), .CK(Clk), .RN(n3853), .Q(
        \pc_target[10][28] ) );
  DFFR_X1 \pc_target_reg[10][30]  ( .D(n6162), .CK(Clk), .RN(n3852), .Q(
        \pc_target[10][30] ) );
  DFFR_X1 \pc_target_reg[11][31]  ( .D(n6161), .CK(Clk), .RN(n3864), .Q(
        \pc_target[11][31] ) );
  DFFR_X1 \pc_target_reg[11][29]  ( .D(n6160), .CK(Clk), .RN(n3852), .Q(
        \pc_target[11][29] ) );
  DFFR_X1 \pc_target_reg[11][27]  ( .D(n6159), .CK(Clk), .RN(n3852), .Q(
        \pc_target[11][27] ) );
  DFFR_X1 \pc_target_reg[11][25]  ( .D(n6158), .CK(Clk), .RN(n3852), .Q(
        \pc_target[11][25] ) );
  DFFR_X1 \pc_target_reg[11][23]  ( .D(n6157), .CK(Clk), .RN(n3853), .Q(
        \pc_target[11][23] ) );
  DFFR_X1 \pc_target_reg[11][21]  ( .D(n6156), .CK(Clk), .RN(n3853), .Q(
        \pc_target[11][21] ) );
  DFFR_X1 \pc_target_reg[11][19]  ( .D(n6155), .CK(Clk), .RN(n3853), .Q(
        \pc_target[11][19] ) );
  DFFR_X1 \pc_target_reg[11][17]  ( .D(n6154), .CK(Clk), .RN(n3853), .Q(
        \pc_target[11][17] ) );
  DFFR_X1 \pc_target_reg[11][15]  ( .D(n6153), .CK(Clk), .RN(n3853), .Q(
        \pc_target[11][15] ) );
  DFFR_X1 \pc_target_reg[11][13]  ( .D(n6152), .CK(Clk), .RN(n3853), .Q(
        \pc_target[11][13] ) );
  DFFR_X1 \pc_target_reg[11][11]  ( .D(n6151), .CK(Clk), .RN(n3853), .Q(
        \pc_target[11][11] ) );
  DFFR_X1 \pc_target_reg[11][9]  ( .D(n6150), .CK(Clk), .RN(n3853), .Q(
        \pc_target[11][9] ) );
  DFFR_X1 \pc_target_reg[11][7]  ( .D(n6149), .CK(Clk), .RN(n3853), .Q(
        \pc_target[11][7] ) );
  DFFR_X1 \pc_target_reg[11][5]  ( .D(n6148), .CK(Clk), .RN(n3853), .Q(
        \pc_target[11][5] ) );
  DFFR_X1 \pc_target_reg[11][3]  ( .D(n6147), .CK(Clk), .RN(n3853), .Q(
        \pc_target[11][3] ) );
  DFFR_X1 \pc_target_reg[11][1]  ( .D(n6146), .CK(Clk), .RN(n3853), .Q(
        \pc_target[11][1] ) );
  DFFR_X1 \pc_target_reg[11][0]  ( .D(n6145), .CK(Clk), .RN(n3854), .Q(
        \pc_target[11][0] ) );
  DFFR_X1 \pc_target_reg[11][2]  ( .D(n6144), .CK(Clk), .RN(n3854), .Q(
        \pc_target[11][2] ) );
  DFFR_X1 \pc_target_reg[11][4]  ( .D(n6143), .CK(Clk), .RN(n3854), .Q(
        \pc_target[11][4] ) );
  DFFR_X1 \pc_target_reg[11][6]  ( .D(n6142), .CK(Clk), .RN(n3854), .Q(
        \pc_target[11][6] ) );
  DFFR_X1 \pc_target_reg[11][8]  ( .D(n6141), .CK(Clk), .RN(n3854), .Q(
        \pc_target[11][8] ) );
  DFFR_X1 \pc_target_reg[11][10]  ( .D(n6140), .CK(Clk), .RN(n3854), .Q(
        \pc_target[11][10] ) );
  DFFR_X1 \pc_target_reg[11][12]  ( .D(n6139), .CK(Clk), .RN(n3854), .Q(
        \pc_target[11][12] ) );
  DFFR_X1 \pc_target_reg[11][14]  ( .D(n6138), .CK(Clk), .RN(n3854), .Q(
        \pc_target[11][14] ) );
  DFFR_X1 \pc_target_reg[11][16]  ( .D(n6137), .CK(Clk), .RN(n3854), .Q(
        \pc_target[11][16] ) );
  DFFR_X1 \pc_target_reg[11][18]  ( .D(n6136), .CK(Clk), .RN(n3854), .Q(
        \pc_target[11][18] ) );
  DFFR_X1 \pc_target_reg[11][20]  ( .D(n6135), .CK(Clk), .RN(n3854), .Q(
        \pc_target[11][20] ) );
  DFFR_X1 \pc_target_reg[11][22]  ( .D(n6134), .CK(Clk), .RN(n3854), .Q(
        \pc_target[11][22] ) );
  DFFR_X1 \pc_target_reg[11][24]  ( .D(n6133), .CK(Clk), .RN(n3854), .Q(
        \pc_target[11][24] ) );
  DFFR_X1 \pc_target_reg[11][26]  ( .D(n6132), .CK(Clk), .RN(n3854), .Q(
        \pc_target[11][26] ) );
  DFFR_X1 \pc_target_reg[11][28]  ( .D(n6131), .CK(Clk), .RN(n3854), .Q(
        \pc_target[11][28] ) );
  DFFR_X1 \pc_target_reg[11][30]  ( .D(n6130), .CK(Clk), .RN(n3855), .Q(
        \pc_target[11][30] ) );
  DFFR_X1 \pc_target_reg[12][31]  ( .D(n6129), .CK(Clk), .RN(n3865), .QN(n730)
         );
  DFFR_X1 \pc_target_reg[12][29]  ( .D(n6128), .CK(Clk), .RN(n3855), .QN(n729)
         );
  DFFR_X1 \pc_target_reg[12][27]  ( .D(n6127), .CK(Clk), .RN(n3855), .QN(n728)
         );
  DFFR_X1 \pc_target_reg[12][25]  ( .D(n6126), .CK(Clk), .RN(n3855), .QN(n727)
         );
  DFFR_X1 \pc_target_reg[12][23]  ( .D(n6125), .CK(Clk), .RN(n3855), .QN(n726)
         );
  DFFR_X1 \pc_target_reg[12][21]  ( .D(n6124), .CK(Clk), .RN(n3855), .QN(n725)
         );
  DFFR_X1 \pc_target_reg[12][19]  ( .D(n6123), .CK(Clk), .RN(n3855), .QN(n724)
         );
  DFFR_X1 \pc_target_reg[12][17]  ( .D(n6122), .CK(Clk), .RN(n3855), .QN(n723)
         );
  DFFR_X1 \pc_target_reg[12][15]  ( .D(n6121), .CK(Clk), .RN(n3855), .QN(n722)
         );
  DFFR_X1 \pc_target_reg[12][13]  ( .D(n6120), .CK(Clk), .RN(n3843), .QN(n721)
         );
  DFFR_X1 \pc_target_reg[12][11]  ( .D(n6119), .CK(Clk), .RN(n3840), .QN(n720)
         );
  DFFR_X1 \pc_target_reg[12][9]  ( .D(n6118), .CK(Clk), .RN(n3840), .QN(n719)
         );
  DFFR_X1 \pc_target_reg[12][7]  ( .D(n6117), .CK(Clk), .RN(n3840), .QN(n718)
         );
  DFFR_X1 \pc_target_reg[12][5]  ( .D(n6116), .CK(Clk), .RN(n3840), .QN(n717)
         );
  DFFR_X1 \pc_target_reg[12][3]  ( .D(n6115), .CK(Clk), .RN(n3840), .QN(n716)
         );
  DFFR_X1 \pc_target_reg[12][1]  ( .D(n6114), .CK(Clk), .RN(n3840), .QN(n715)
         );
  DFFR_X1 \pc_target_reg[12][0]  ( .D(n6113), .CK(Clk), .RN(n3840), .QN(n714)
         );
  DFFR_X1 \pc_target_reg[12][2]  ( .D(n6112), .CK(Clk), .RN(n3840), .QN(n713)
         );
  DFFR_X1 \pc_target_reg[12][4]  ( .D(n6111), .CK(Clk), .RN(n3840), .QN(n712)
         );
  DFFR_X1 \pc_target_reg[12][6]  ( .D(n6110), .CK(Clk), .RN(n3840), .QN(n711)
         );
  DFFR_X1 \pc_target_reg[12][8]  ( .D(n6109), .CK(Clk), .RN(n3840), .QN(n710)
         );
  DFFR_X1 \pc_target_reg[12][10]  ( .D(n6108), .CK(Clk), .RN(n3840), .QN(n709)
         );
  DFFR_X1 \pc_target_reg[12][12]  ( .D(n6107), .CK(Clk), .RN(n3840), .QN(n708)
         );
  DFFR_X1 \pc_target_reg[12][14]  ( .D(n6106), .CK(Clk), .RN(n3841), .QN(n707)
         );
  DFFR_X1 \pc_target_reg[12][16]  ( .D(n6105), .CK(Clk), .RN(n3841), .QN(n706)
         );
  DFFR_X1 \pc_target_reg[12][18]  ( .D(n6104), .CK(Clk), .RN(n3841), .QN(n705)
         );
  DFFR_X1 \pc_target_reg[12][20]  ( .D(n6103), .CK(Clk), .RN(n3841), .QN(n704)
         );
  DFFR_X1 \pc_target_reg[12][22]  ( .D(n6102), .CK(Clk), .RN(n3841), .QN(n703)
         );
  DFFR_X1 \pc_target_reg[12][24]  ( .D(n6101), .CK(Clk), .RN(n3841), .QN(n702)
         );
  DFFR_X1 \pc_target_reg[12][26]  ( .D(n6100), .CK(Clk), .RN(n3841), .QN(n701)
         );
  DFFR_X1 \pc_target_reg[12][28]  ( .D(n6099), .CK(Clk), .RN(n3841), .QN(n700)
         );
  DFFR_X1 \pc_target_reg[13][31]  ( .D(n6097), .CK(Clk), .RN(n3865), .QN(n696)
         );
  DFFR_X1 \pc_target_reg[13][29]  ( .D(n6096), .CK(Clk), .RN(n3841), .QN(n695)
         );
  DFFR_X1 \pc_target_reg[13][27]  ( .D(n6095), .CK(Clk), .RN(n3877), .QN(n694)
         );
  DFFR_X1 \pc_target_reg[13][25]  ( .D(n6094), .CK(Clk), .RN(n3877), .QN(n693)
         );
  DFFR_X1 \pc_target_reg[13][23]  ( .D(n6093), .CK(Clk), .RN(n3877), .QN(n692)
         );
  DFFR_X1 \pc_target_reg[13][21]  ( .D(n6092), .CK(Clk), .RN(n3877), .QN(n691)
         );
  DFFR_X1 \pc_target_reg[13][19]  ( .D(n6091), .CK(Clk), .RN(n3877), .QN(n690)
         );
  DFFR_X1 \pc_target_reg[13][17]  ( .D(n6090), .CK(Clk), .RN(n3877), .QN(n689)
         );
  DFFR_X1 \pc_target_reg[13][15]  ( .D(n6089), .CK(Clk), .RN(n3878), .QN(n688)
         );
  DFFR_X1 \pc_target_reg[13][13]  ( .D(n6088), .CK(Clk), .RN(n3878), .QN(n687)
         );
  DFFR_X1 \pc_target_reg[13][11]  ( .D(n6087), .CK(Clk), .RN(n3878), .QN(n686)
         );
  DFFR_X1 \pc_target_reg[13][9]  ( .D(n6086), .CK(Clk), .RN(n3878), .QN(n685)
         );
  DFFR_X1 \pc_target_reg[13][7]  ( .D(n6085), .CK(Clk), .RN(n3878), .QN(n684)
         );
  DFFR_X1 \pc_target_reg[13][5]  ( .D(n6084), .CK(Clk), .RN(n3878), .QN(n683)
         );
  DFFR_X1 \pc_target_reg[13][3]  ( .D(n6083), .CK(Clk), .RN(n3878), .QN(n682)
         );
  DFFR_X1 \pc_target_reg[13][1]  ( .D(n6082), .CK(Clk), .RN(n3878), .QN(n681)
         );
  DFFR_X1 \pc_target_reg[13][0]  ( .D(n6081), .CK(Clk), .RN(n3879), .QN(n680)
         );
  DFFR_X1 \pc_target_reg[13][2]  ( .D(n6080), .CK(Clk), .RN(n3878), .QN(n679)
         );
  DFFR_X1 \pc_target_reg[13][4]  ( .D(n6079), .CK(Clk), .RN(n3878), .QN(n678)
         );
  DFFR_X1 \pc_target_reg[13][6]  ( .D(n6078), .CK(Clk), .RN(n3878), .QN(n677)
         );
  DFFR_X1 \pc_target_reg[13][8]  ( .D(n6077), .CK(Clk), .RN(n3878), .QN(n676)
         );
  DFFR_X1 \pc_target_reg[13][10]  ( .D(n6076), .CK(Clk), .RN(n3878), .QN(n675)
         );
  DFFR_X1 \pc_target_reg[13][12]  ( .D(n6075), .CK(Clk), .RN(n3878), .QN(n674)
         );
  DFFR_X1 \pc_target_reg[13][14]  ( .D(n6074), .CK(Clk), .RN(n3878), .QN(n673)
         );
  DFFR_X1 \pc_target_reg[13][16]  ( .D(n6073), .CK(Clk), .RN(n3879), .QN(n672)
         );
  DFFR_X1 \pc_target_reg[13][18]  ( .D(n6072), .CK(Clk), .RN(n3879), .QN(n671)
         );
  DFFR_X1 \pc_target_reg[13][20]  ( .D(n6071), .CK(Clk), .RN(n3879), .QN(n670)
         );
  DFFR_X1 \pc_target_reg[13][22]  ( .D(n6070), .CK(Clk), .RN(n3879), .QN(n669)
         );
  DFFR_X1 \pc_target_reg[13][24]  ( .D(n6069), .CK(Clk), .RN(n3879), .QN(n668)
         );
  DFFR_X1 \pc_target_reg[13][26]  ( .D(n6068), .CK(Clk), .RN(n3879), .QN(n667)
         );
  DFFR_X1 \pc_target_reg[13][28]  ( .D(n6067), .CK(Clk), .RN(n3879), .QN(n666)
         );
  DFFR_X1 \pc_target_reg[14][31]  ( .D(n6065), .CK(Clk), .RN(n3864), .Q(
        \pc_target[14][31] ) );
  DFFR_X1 \pc_target_reg[14][29]  ( .D(n6064), .CK(Clk), .RN(n3879), .Q(
        \pc_target[14][29] ) );
  DFFR_X1 \pc_target_reg[14][27]  ( .D(n6063), .CK(Clk), .RN(n3879), .Q(
        \pc_target[14][27] ) );
  DFFR_X1 \pc_target_reg[14][25]  ( .D(n6062), .CK(Clk), .RN(n3879), .Q(
        \pc_target[14][25] ) );
  DFFR_X1 \pc_target_reg[14][23]  ( .D(n6061), .CK(Clk), .RN(n3879), .Q(
        \pc_target[14][23] ) );
  DFFR_X1 \pc_target_reg[14][21]  ( .D(n6060), .CK(Clk), .RN(n3879), .Q(
        \pc_target[14][21] ) );
  DFFR_X1 \pc_target_reg[14][19]  ( .D(n6059), .CK(Clk), .RN(n3879), .Q(
        \pc_target[14][19] ) );
  DFFR_X1 \pc_target_reg[14][17]  ( .D(n6058), .CK(Clk), .RN(n3879), .Q(
        \pc_target[14][17] ) );
  DFFR_X1 \pc_target_reg[14][15]  ( .D(n6057), .CK(Clk), .RN(n3880), .Q(
        \pc_target[14][15] ) );
  DFFR_X1 \pc_target_reg[14][13]  ( .D(n6056), .CK(Clk), .RN(n3840), .Q(
        \pc_target[14][13] ) );
  DFFR_X1 \pc_target_reg[14][11]  ( .D(n6055), .CK(Clk), .RN(n3836), .Q(
        \pc_target[14][11] ) );
  DFFR_X1 \pc_target_reg[14][9]  ( .D(n6054), .CK(Clk), .RN(n3832), .Q(
        \pc_target[14][9] ) );
  DFFR_X1 \pc_target_reg[14][7]  ( .D(n6053), .CK(Clk), .RN(n3832), .Q(
        \pc_target[14][7] ) );
  DFFR_X1 \pc_target_reg[14][5]  ( .D(n6052), .CK(Clk), .RN(n3832), .Q(
        \pc_target[14][5] ) );
  DFFR_X1 \pc_target_reg[14][3]  ( .D(n6051), .CK(Clk), .RN(n3832), .Q(
        \pc_target[14][3] ) );
  DFFR_X1 \pc_target_reg[14][1]  ( .D(n6050), .CK(Clk), .RN(n3832), .Q(
        \pc_target[14][1] ) );
  DFFR_X1 \pc_target_reg[14][0]  ( .D(n6049), .CK(Clk), .RN(n3832), .Q(
        \pc_target[14][0] ) );
  DFFR_X1 \pc_target_reg[14][2]  ( .D(n6048), .CK(Clk), .RN(n3832), .Q(
        \pc_target[14][2] ) );
  DFFR_X1 \pc_target_reg[14][4]  ( .D(n6047), .CK(Clk), .RN(n3832), .Q(
        \pc_target[14][4] ) );
  DFFR_X1 \pc_target_reg[14][6]  ( .D(n6046), .CK(Clk), .RN(n3832), .Q(
        \pc_target[14][6] ) );
  DFFR_X1 \pc_target_reg[14][8]  ( .D(n6045), .CK(Clk), .RN(n3833), .Q(
        \pc_target[14][8] ) );
  DFFR_X1 \pc_target_reg[14][10]  ( .D(n6044), .CK(Clk), .RN(n3833), .Q(
        \pc_target[14][10] ) );
  DFFR_X1 \pc_target_reg[14][12]  ( .D(n6043), .CK(Clk), .RN(n3833), .Q(
        \pc_target[14][12] ) );
  DFFR_X1 \pc_target_reg[14][14]  ( .D(n6042), .CK(Clk), .RN(n3833), .Q(
        \pc_target[14][14] ) );
  DFFR_X1 \pc_target_reg[14][16]  ( .D(n6041), .CK(Clk), .RN(n3833), .Q(
        \pc_target[14][16] ) );
  DFFR_X1 \pc_target_reg[14][18]  ( .D(n6040), .CK(Clk), .RN(n3833), .Q(
        \pc_target[14][18] ) );
  DFFR_X1 \pc_target_reg[14][20]  ( .D(n6039), .CK(Clk), .RN(n3833), .Q(
        \pc_target[14][20] ) );
  DFFR_X1 \pc_target_reg[14][22]  ( .D(n6038), .CK(Clk), .RN(n3833), .Q(
        \pc_target[14][22] ) );
  DFFR_X1 \pc_target_reg[14][24]  ( .D(n6037), .CK(Clk), .RN(n3833), .Q(
        \pc_target[14][24] ) );
  DFFR_X1 \pc_target_reg[14][26]  ( .D(n6036), .CK(Clk), .RN(n3833), .Q(
        \pc_target[14][26] ) );
  DFFR_X1 \pc_target_reg[14][28]  ( .D(n6035), .CK(Clk), .RN(n3833), .Q(
        \pc_target[14][28] ) );
  DFFR_X1 \pc_target_reg[14][30]  ( .D(n6034), .CK(Clk), .RN(n3834), .Q(
        \pc_target[14][30] ) );
  DFFR_X1 \pc_target_reg[15][31]  ( .D(n6033), .CK(Clk), .RN(n3864), .Q(
        \pc_target[15][31] ) );
  DFFR_X1 \pc_target_reg[15][29]  ( .D(n6032), .CK(Clk), .RN(n3833), .Q(
        \pc_target[15][29] ) );
  DFFR_X1 \pc_target_reg[15][27]  ( .D(n6031), .CK(Clk), .RN(n3833), .Q(
        \pc_target[15][27] ) );
  DFFR_X1 \pc_target_reg[15][25]  ( .D(n6030), .CK(Clk), .RN(n3833), .Q(
        \pc_target[15][25] ) );
  DFFR_X1 \pc_target_reg[15][23]  ( .D(n6029), .CK(Clk), .RN(n3833), .Q(
        \pc_target[15][23] ) );
  DFFR_X1 \pc_target_reg[15][21]  ( .D(n6028), .CK(Clk), .RN(n3834), .Q(
        \pc_target[15][21] ) );
  DFFR_X1 \pc_target_reg[15][19]  ( .D(n6027), .CK(Clk), .RN(n3834), .Q(
        \pc_target[15][19] ) );
  DFFR_X1 \pc_target_reg[15][17]  ( .D(n6026), .CK(Clk), .RN(n3834), .Q(
        \pc_target[15][17] ) );
  DFFR_X1 \pc_target_reg[15][15]  ( .D(n6025), .CK(Clk), .RN(n3834), .Q(
        \pc_target[15][15] ) );
  DFFR_X1 \pc_target_reg[15][13]  ( .D(n6024), .CK(Clk), .RN(n3834), .Q(
        \pc_target[15][13] ) );
  DFFR_X1 \pc_target_reg[15][11]  ( .D(n6023), .CK(Clk), .RN(n3834), .Q(
        \pc_target[15][11] ) );
  DFFR_X1 \pc_target_reg[15][7]  ( .D(n6021), .CK(Clk), .RN(n3838), .Q(
        \pc_target[15][7] ) );
  DFFR_X1 \pc_target_reg[15][12]  ( .D(n6011), .CK(Clk), .RN(n3838), .Q(
        \pc_target[15][12] ) );
  DFFR_X1 \pc_target_reg[15][14]  ( .D(n6010), .CK(Clk), .RN(n3838), .Q(
        \pc_target[15][14] ) );
  DFFR_X1 \pc_target_reg[15][16]  ( .D(n6009), .CK(Clk), .RN(n3834), .Q(
        \pc_target[15][16] ) );
  DFFR_X1 \pc_target_reg[15][18]  ( .D(n6008), .CK(Clk), .RN(n3834), .Q(
        \pc_target[15][18] ) );
  DFFR_X1 \pc_target_reg[15][20]  ( .D(n6007), .CK(Clk), .RN(n3834), .Q(
        \pc_target[15][20] ) );
  DFFR_X1 \pc_target_reg[15][22]  ( .D(n6006), .CK(Clk), .RN(n3834), .Q(
        \pc_target[15][22] ) );
  DFFR_X1 \pc_target_reg[15][24]  ( .D(n6005), .CK(Clk), .RN(n3834), .Q(
        \pc_target[15][24] ) );
  DFFR_X1 \pc_target_reg[15][26]  ( .D(n6004), .CK(Clk), .RN(n3834), .Q(
        \pc_target[15][26] ) );
  DFFR_X1 \pc_target_reg[15][28]  ( .D(n6003), .CK(Clk), .RN(n3834), .Q(
        \pc_target[15][28] ) );
  DFFR_X1 \pc_target_reg[15][30]  ( .D(n6002), .CK(Clk), .RN(n3834), .Q(
        \pc_target[15][30] ) );
  DFFR_X1 \pc_target_reg[16][31]  ( .D(n6001), .CK(Clk), .RN(n3865), .QN(n591)
         );
  DFFR_X1 \pc_target_reg[16][29]  ( .D(n6000), .CK(Clk), .RN(n3835), .QN(n590)
         );
  DFFR_X1 \pc_target_reg[16][27]  ( .D(n5999), .CK(Clk), .RN(n3835), .QN(n589)
         );
  DFFR_X1 \pc_target_reg[16][25]  ( .D(n5998), .CK(Clk), .RN(n3835), .QN(n588)
         );
  DFFR_X1 \pc_target_reg[16][23]  ( .D(n5997), .CK(Clk), .RN(n3835), .QN(n587)
         );
  DFFR_X1 \pc_target_reg[16][21]  ( .D(n5996), .CK(Clk), .RN(n3835), .QN(n586)
         );
  DFFR_X1 \pc_target_reg[16][19]  ( .D(n5995), .CK(Clk), .RN(n3835), .QN(n585)
         );
  DFFR_X1 \pc_target_reg[16][17]  ( .D(n5994), .CK(Clk), .RN(n3835), .QN(n584)
         );
  DFFR_X1 \pc_target_reg[16][15]  ( .D(n5993), .CK(Clk), .RN(n3835), .QN(n583)
         );
  DFFR_X1 \pc_target_reg[16][13]  ( .D(n5992), .CK(Clk), .RN(n3835), .QN(n582)
         );
  DFFR_X1 \pc_target_reg[16][11]  ( .D(n5991), .CK(Clk), .RN(n3835), .QN(n581)
         );
  DFFR_X1 \pc_target_reg[16][9]  ( .D(n5990), .CK(Clk), .RN(n3835), .QN(n580)
         );
  DFFR_X1 \pc_target_reg[16][7]  ( .D(n5989), .CK(Clk), .RN(n3835), .QN(n579)
         );
  DFFR_X1 \pc_target_reg[16][5]  ( .D(n5988), .CK(Clk), .RN(n3835), .QN(n578)
         );
  DFFR_X1 \pc_target_reg[16][3]  ( .D(n5987), .CK(Clk), .RN(n3835), .QN(n577)
         );
  DFFR_X1 \pc_target_reg[16][1]  ( .D(n5986), .CK(Clk), .RN(n3835), .QN(n576)
         );
  DFFR_X1 \pc_target_reg[16][0]  ( .D(n5985), .CK(Clk), .RN(n3836), .QN(n575)
         );
  DFFR_X1 \pc_target_reg[16][2]  ( .D(n5984), .CK(Clk), .RN(n3836), .QN(n574)
         );
  DFFR_X1 \pc_target_reg[16][4]  ( .D(n5983), .CK(Clk), .RN(n3836), .QN(n573)
         );
  DFFR_X1 \pc_target_reg[16][6]  ( .D(n5982), .CK(Clk), .RN(n3836), .QN(n572)
         );
  DFFR_X1 \pc_target_reg[16][8]  ( .D(n5981), .CK(Clk), .RN(n3836), .QN(n571)
         );
  DFFR_X1 \pc_target_reg[16][10]  ( .D(n5980), .CK(Clk), .RN(n3836), .QN(n570)
         );
  DFFR_X1 \pc_target_reg[16][12]  ( .D(n5979), .CK(Clk), .RN(n3836), .QN(n569)
         );
  DFFR_X1 \pc_target_reg[16][14]  ( .D(n5978), .CK(Clk), .RN(n3836), .QN(n568)
         );
  DFFR_X1 \pc_target_reg[16][16]  ( .D(n5977), .CK(Clk), .RN(n3836), .QN(n567)
         );
  DFFR_X1 \pc_target_reg[16][18]  ( .D(n5976), .CK(Clk), .RN(n3836), .QN(n566)
         );
  DFFR_X1 \pc_target_reg[16][20]  ( .D(n5975), .CK(Clk), .RN(n3836), .QN(n565)
         );
  DFFR_X1 \pc_target_reg[16][24]  ( .D(n5973), .CK(Clk), .RN(n3836), .QN(n563)
         );
  DFFR_X1 \pc_target_reg[16][26]  ( .D(n5972), .CK(Clk), .RN(n3836), .QN(n562)
         );
  DFFR_X1 \pc_target_reg[16][28]  ( .D(n5971), .CK(Clk), .RN(n3837), .QN(n561)
         );
  DFFR_X1 \pc_target_reg[17][31]  ( .D(n5969), .CK(Clk), .RN(n3865), .QN(n557)
         );
  DFFR_X1 \pc_target_reg[17][29]  ( .D(n5968), .CK(Clk), .RN(n3837), .QN(n556)
         );
  DFFR_X1 \pc_target_reg[17][27]  ( .D(n5967), .CK(Clk), .RN(n3837), .QN(n555)
         );
  DFFR_X1 \pc_target_reg[17][25]  ( .D(n5966), .CK(Clk), .RN(n3837), .QN(n554)
         );
  DFFR_X1 \pc_target_reg[17][23]  ( .D(n5965), .CK(Clk), .RN(n3837), .QN(n553)
         );
  DFFR_X1 \pc_target_reg[17][21]  ( .D(n5964), .CK(Clk), .RN(n3837), .QN(n552)
         );
  DFFR_X1 \pc_target_reg[17][19]  ( .D(n5963), .CK(Clk), .RN(n3837), .QN(n551)
         );
  DFFR_X1 \pc_target_reg[17][17]  ( .D(n5962), .CK(Clk), .RN(n3837), .QN(n550)
         );
  DFFR_X1 \pc_target_reg[17][15]  ( .D(n5961), .CK(Clk), .RN(n3837), .QN(n549)
         );
  DFFR_X1 \pc_target_reg[17][13]  ( .D(n5960), .CK(Clk), .RN(n3837), .QN(n548)
         );
  DFFR_X1 \pc_target_reg[17][11]  ( .D(n5959), .CK(Clk), .RN(n3837), .QN(n547)
         );
  DFFR_X1 \pc_target_reg[17][9]  ( .D(n5958), .CK(Clk), .RN(n3837), .QN(n546)
         );
  DFFR_X1 \pc_target_reg[17][7]  ( .D(n5957), .CK(Clk), .RN(n3837), .QN(n545)
         );
  DFFR_X1 \pc_target_reg[17][3]  ( .D(n5955), .CK(Clk), .RN(n3837), .QN(n543)
         );
  DFFR_X1 \pc_target_reg[17][1]  ( .D(n5954), .CK(Clk), .RN(n3837), .QN(n542)
         );
  DFFR_X1 \pc_target_reg[17][0]  ( .D(n5953), .CK(Clk), .RN(n3838), .QN(n541)
         );
  DFFR_X1 \pc_target_reg[17][2]  ( .D(n5952), .CK(Clk), .RN(n3838), .QN(n540)
         );
  DFFR_X1 \pc_target_reg[17][6]  ( .D(n5950), .CK(Clk), .RN(n3838), .QN(n538)
         );
  DFFR_X1 \pc_target_reg[17][8]  ( .D(n5949), .CK(Clk), .RN(n3838), .QN(n537)
         );
  DFFR_X1 \pc_target_reg[17][10]  ( .D(n5948), .CK(Clk), .RN(n3838), .QN(n536)
         );
  DFFR_X1 \pc_target_reg[17][12]  ( .D(n5947), .CK(Clk), .RN(n3838), .QN(n535)
         );
  DFFR_X1 \pc_target_reg[17][14]  ( .D(n5946), .CK(Clk), .RN(n3838), .QN(n534)
         );
  DFFR_X1 \pc_target_reg[17][16]  ( .D(n5945), .CK(Clk), .RN(n3838), .QN(n533)
         );
  DFFR_X1 \pc_target_reg[17][18]  ( .D(n5944), .CK(Clk), .RN(n3838), .QN(n532)
         );
  DFFR_X1 \pc_target_reg[17][20]  ( .D(n5943), .CK(Clk), .RN(n3838), .QN(n531)
         );
  DFFR_X1 \pc_target_reg[17][22]  ( .D(n5942), .CK(Clk), .RN(n3838), .QN(n530)
         );
  DFFR_X1 \pc_target_reg[17][24]  ( .D(n5941), .CK(Clk), .RN(n3838), .QN(n529)
         );
  DFFR_X1 \pc_target_reg[17][26]  ( .D(n5940), .CK(Clk), .RN(n3839), .QN(n528)
         );
  DFFR_X1 \pc_target_reg[17][28]  ( .D(n5939), .CK(Clk), .RN(n3839), .QN(n527)
         );
  DFFR_X1 \pc_target_reg[18][31]  ( .D(n5937), .CK(Clk), .RN(n3864), .Q(
        \pc_target[18][31] ) );
  DFFR_X1 \pc_target_reg[18][29]  ( .D(n5936), .CK(Clk), .RN(n3839), .Q(
        \pc_target[18][29] ) );
  DFFR_X1 \pc_target_reg[18][27]  ( .D(n5935), .CK(Clk), .RN(n3839), .Q(
        \pc_target[18][27] ) );
  DFFR_X1 \pc_target_reg[18][25]  ( .D(n5934), .CK(Clk), .RN(n3839), .Q(
        \pc_target[18][25] ) );
  DFFR_X1 \pc_target_reg[18][23]  ( .D(n5933), .CK(Clk), .RN(n3839), .Q(
        \pc_target[18][23] ) );
  DFFR_X1 \pc_target_reg[18][21]  ( .D(n5932), .CK(Clk), .RN(n3839), .Q(
        \pc_target[18][21] ) );
  DFFR_X1 \pc_target_reg[18][19]  ( .D(n5931), .CK(Clk), .RN(n3839), .Q(
        \pc_target[18][19] ) );
  DFFR_X1 \pc_target_reg[18][17]  ( .D(n5930), .CK(Clk), .RN(n3839), .Q(
        \pc_target[18][17] ) );
  DFFR_X1 \pc_target_reg[18][15]  ( .D(n5929), .CK(Clk), .RN(n3839), .Q(
        \pc_target[18][15] ) );
  DFFR_X1 \pc_target_reg[18][13]  ( .D(n5928), .CK(Clk), .RN(n3839), .Q(
        \pc_target[18][13] ) );
  DFFR_X1 \pc_target_reg[18][11]  ( .D(n5927), .CK(Clk), .RN(n3839), .Q(
        \pc_target[18][11] ) );
  DFFR_X1 \pc_target_reg[18][9]  ( .D(n5926), .CK(Clk), .RN(n3839), .Q(
        \pc_target[18][9] ) );
  DFFR_X1 \pc_target_reg[18][7]  ( .D(n5925), .CK(Clk), .RN(n3839), .Q(
        \pc_target[18][7] ) );
  DFFR_X1 \pc_target_reg[18][5]  ( .D(n5924), .CK(Clk), .RN(n3839), .Q(
        \pc_target[18][5] ) );
  DFFR_X1 \pc_target_reg[18][3]  ( .D(n5923), .CK(Clk), .RN(n3840), .Q(
        \pc_target[18][3] ) );
  DFFR_X1 \pc_target_reg[18][1]  ( .D(n5922), .CK(Clk), .RN(n3829), .Q(
        \pc_target[18][1] ) );
  DFFR_X1 \pc_target_reg[18][0]  ( .D(n5921), .CK(Clk), .RN(n3826), .Q(
        \pc_target[18][0] ) );
  DFFR_X1 \pc_target_reg[18][2]  ( .D(n5920), .CK(Clk), .RN(n3828), .Q(
        \pc_target[18][2] ) );
  DFFR_X1 \pc_target_reg[18][4]  ( .D(n5919), .CK(Clk), .RN(n3826), .Q(
        \pc_target[18][4] ) );
  DFFR_X1 \pc_target_reg[18][6]  ( .D(n5918), .CK(Clk), .RN(n3826), .Q(
        \pc_target[18][6] ) );
  DFFR_X1 \pc_target_reg[18][8]  ( .D(n5917), .CK(Clk), .RN(n3826), .Q(
        \pc_target[18][8] ) );
  DFFR_X1 \pc_target_reg[18][10]  ( .D(n5916), .CK(Clk), .RN(n3827), .Q(
        \pc_target[18][10] ) );
  DFFR_X1 \pc_target_reg[18][12]  ( .D(n5915), .CK(Clk), .RN(n3826), .Q(
        \pc_target[18][12] ) );
  DFFR_X1 \pc_target_reg[18][14]  ( .D(n5914), .CK(Clk), .RN(n3828), .Q(
        \pc_target[18][14] ) );
  DFFR_X1 \pc_target_reg[18][16]  ( .D(n5913), .CK(Clk), .RN(n3826), .Q(
        \pc_target[18][16] ) );
  DFFR_X1 \pc_target_reg[18][18]  ( .D(n5912), .CK(Clk), .RN(n3828), .Q(
        \pc_target[18][18] ) );
  DFFR_X1 \pc_target_reg[18][20]  ( .D(n5911), .CK(Clk), .RN(n3828), .Q(
        \pc_target[18][20] ) );
  DFFR_X1 \pc_target_reg[18][22]  ( .D(n5910), .CK(Clk), .RN(n3828), .Q(
        \pc_target[18][22] ) );
  DFFR_X1 \pc_target_reg[18][24]  ( .D(n5909), .CK(Clk), .RN(n3827), .Q(
        \pc_target[18][24] ) );
  DFFR_X1 \pc_target_reg[18][26]  ( .D(n5908), .CK(Clk), .RN(n3827), .Q(
        \pc_target[18][26] ) );
  DFFR_X1 \pc_target_reg[18][28]  ( .D(n5907), .CK(Clk), .RN(n3828), .Q(
        \pc_target[18][28] ) );
  DFFR_X1 \pc_target_reg[18][30]  ( .D(n5906), .CK(Clk), .RN(n3827), .Q(
        \pc_target[18][30] ) );
  DFFR_X1 \pc_target_reg[19][31]  ( .D(n5905), .CK(Clk), .RN(n3864), .Q(
        \pc_target[19][31] ) );
  DFFR_X1 \pc_target_reg[19][29]  ( .D(n5904), .CK(Clk), .RN(n3826), .Q(
        \pc_target[19][29] ) );
  DFFR_X1 \pc_target_reg[19][27]  ( .D(n5903), .CK(Clk), .RN(n3828), .Q(
        \pc_target[19][27] ) );
  DFFR_X1 \pc_target_reg[19][25]  ( .D(n5902), .CK(Clk), .RN(n3827), .Q(
        \pc_target[19][25] ) );
  DFFR_X1 \pc_target_reg[19][23]  ( .D(n5901), .CK(Clk), .RN(n3827), .Q(
        \pc_target[19][23] ) );
  DFFR_X1 \pc_target_reg[19][21]  ( .D(n5900), .CK(Clk), .RN(n3827), .Q(
        \pc_target[19][21] ) );
  DFFR_X1 \pc_target_reg[19][19]  ( .D(n5899), .CK(Clk), .RN(n3829), .Q(
        \pc_target[19][19] ) );
  DFFR_X1 \pc_target_reg[19][17]  ( .D(n5898), .CK(Clk), .RN(n3827), .Q(
        \pc_target[19][17] ) );
  DFFR_X1 \pc_target_reg[19][15]  ( .D(n5897), .CK(Clk), .RN(n3827), .Q(
        \pc_target[19][15] ) );
  DFFR_X1 \pc_target_reg[19][13]  ( .D(n5896), .CK(Clk), .RN(n3828), .Q(
        \pc_target[19][13] ) );
  DFFR_X1 \pc_target_reg[19][11]  ( .D(n5895), .CK(Clk), .RN(n3827), .Q(
        \pc_target[19][11] ) );
  DFFR_X1 \pc_target_reg[19][9]  ( .D(n5894), .CK(Clk), .RN(n3827), .Q(
        \pc_target[19][9] ) );
  DFFR_X1 \pc_target_reg[19][7]  ( .D(n5893), .CK(Clk), .RN(n3828), .Q(
        \pc_target[19][7] ) );
  DFFR_X1 \pc_target_reg[19][5]  ( .D(n5892), .CK(Clk), .RN(n3827), .Q(
        \pc_target[19][5] ) );
  DFFR_X1 \pc_target_reg[19][3]  ( .D(n5891), .CK(Clk), .RN(n3827), .Q(
        \pc_target[19][3] ) );
  DFFR_X1 \pc_target_reg[19][1]  ( .D(n5890), .CK(Clk), .RN(n3828), .Q(
        \pc_target[19][1] ) );
  DFFR_X1 \pc_target_reg[19][0]  ( .D(n5889), .CK(Clk), .RN(n3828), .Q(
        \pc_target[19][0] ) );
  DFFR_X1 \pc_target_reg[19][2]  ( .D(n5888), .CK(Clk), .RN(n3827), .Q(
        \pc_target[19][2] ) );
  DFFR_X1 \pc_target_reg[19][4]  ( .D(n5887), .CK(Clk), .RN(n3829), .Q(
        \pc_target[19][4] ) );
  DFFR_X1 \pc_target_reg[19][6]  ( .D(n5886), .CK(Clk), .RN(n3828), .Q(
        \pc_target[19][6] ) );
  DFFR_X1 \pc_target_reg[19][8]  ( .D(n5885), .CK(Clk), .RN(n3828), .Q(
        \pc_target[19][8] ) );
  DFFR_X1 \pc_target_reg[19][10]  ( .D(n5884), .CK(Clk), .RN(n3828), .Q(
        \pc_target[19][10] ) );
  DFFR_X1 \pc_target_reg[19][12]  ( .D(n5883), .CK(Clk), .RN(n3828), .Q(
        \pc_target[19][12] ) );
  DFFR_X1 \pc_target_reg[19][14]  ( .D(n5882), .CK(Clk), .RN(n3829), .Q(
        \pc_target[19][14] ) );
  DFFR_X1 \pc_target_reg[19][16]  ( .D(n5881), .CK(Clk), .RN(n3829), .Q(
        \pc_target[19][16] ) );
  DFFR_X1 \pc_target_reg[19][18]  ( .D(n5880), .CK(Clk), .RN(n3829), .Q(
        \pc_target[19][18] ) );
  DFFR_X1 \pc_target_reg[19][20]  ( .D(n5879), .CK(Clk), .RN(n3829), .Q(
        \pc_target[19][20] ) );
  DFFR_X1 \pc_target_reg[19][22]  ( .D(n5878), .CK(Clk), .RN(n3829), .Q(
        \pc_target[19][22] ) );
  DFFR_X1 \pc_target_reg[19][24]  ( .D(n5877), .CK(Clk), .RN(n3829), .Q(
        \pc_target[19][24] ) );
  DFFR_X1 \pc_target_reg[19][26]  ( .D(n5876), .CK(Clk), .RN(n3829), .Q(
        \pc_target[19][26] ) );
  DFFR_X1 \pc_target_reg[19][28]  ( .D(n5875), .CK(Clk), .RN(n3829), .Q(
        \pc_target[19][28] ) );
  DFFR_X1 \pc_target_reg[19][30]  ( .D(n5874), .CK(Clk), .RN(n3829), .Q(
        \pc_target[19][30] ) );
  DFFR_X1 \pc_target_reg[20][31]  ( .D(n5873), .CK(Clk), .RN(n3864), .Q(
        \pc_target[20][31] ) );
  DFFR_X1 \pc_target_reg[20][29]  ( .D(n5872), .CK(Clk), .RN(n3880), .Q(
        \pc_target[20][29] ) );
  DFFR_X1 \pc_target_reg[20][27]  ( .D(n5871), .CK(Clk), .RN(n3880), .Q(
        \pc_target[20][27] ) );
  DFFR_X1 \pc_target_reg[20][25]  ( .D(n5870), .CK(Clk), .RN(n3880), .Q(
        \pc_target[20][25] ) );
  DFFR_X1 \pc_target_reg[20][23]  ( .D(n5869), .CK(Clk), .RN(n3880), .Q(
        \pc_target[20][23] ) );
  DFFR_X1 \pc_target_reg[20][21]  ( .D(n5868), .CK(Clk), .RN(n3880), .Q(
        \pc_target[20][21] ) );
  DFFR_X1 \pc_target_reg[20][19]  ( .D(n5867), .CK(Clk), .RN(n3880), .Q(
        \pc_target[20][19] ) );
  DFFR_X1 \pc_target_reg[20][17]  ( .D(n5866), .CK(Clk), .RN(n3880), .Q(
        \pc_target[20][17] ) );
  DFFR_X1 \pc_target_reg[20][15]  ( .D(n5865), .CK(Clk), .RN(n3880), .Q(
        \pc_target[20][15] ) );
  DFFR_X1 \pc_target_reg[20][13]  ( .D(n5864), .CK(Clk), .RN(n3880), .Q(
        \pc_target[20][13] ) );
  DFFR_X1 \pc_target_reg[20][11]  ( .D(n5863), .CK(Clk), .RN(n3880), .Q(
        \pc_target[20][11] ) );
  DFFR_X1 \pc_target_reg[20][9]  ( .D(n5862), .CK(Clk), .RN(n3880), .Q(
        \pc_target[20][9] ) );
  DFFR_X1 \pc_target_reg[20][7]  ( .D(n5861), .CK(Clk), .RN(n3880), .Q(
        \pc_target[20][7] ) );
  DFFR_X1 \pc_target_reg[20][5]  ( .D(n5860), .CK(Clk), .RN(n3881), .Q(
        \pc_target[20][5] ) );
  DFFR_X1 \pc_target_reg[20][3]  ( .D(n5859), .CK(Clk), .RN(n3881), .Q(
        \pc_target[20][3] ) );
  DFFR_X1 \pc_target_reg[20][1]  ( .D(n5858), .CK(Clk), .RN(n3881), .Q(
        \pc_target[20][1] ) );
  DFFR_X1 \pc_target_reg[20][0]  ( .D(n5857), .CK(Clk), .RN(n3881), .Q(
        \pc_target[20][0] ) );
  DFFR_X1 \pc_target_reg[20][2]  ( .D(n5856), .CK(Clk), .RN(n3881), .Q(
        \pc_target[20][2] ) );
  DFFR_X1 \pc_target_reg[20][4]  ( .D(n5855), .CK(Clk), .RN(n3881), .Q(
        \pc_target[20][4] ) );
  DFFR_X1 \pc_target_reg[20][6]  ( .D(n5854), .CK(Clk), .RN(n3881), .Q(
        \pc_target[20][6] ) );
  DFFR_X1 \pc_target_reg[20][8]  ( .D(n5853), .CK(Clk), .RN(n3881), .Q(
        \pc_target[20][8] ) );
  DFFR_X1 \pc_target_reg[20][10]  ( .D(n5852), .CK(Clk), .RN(n3881), .Q(
        \pc_target[20][10] ) );
  DFFR_X1 \pc_target_reg[20][12]  ( .D(n5851), .CK(Clk), .RN(n3881), .Q(
        \pc_target[20][12] ) );
  DFFR_X1 \pc_target_reg[20][14]  ( .D(n5850), .CK(Clk), .RN(n3881), .Q(
        \pc_target[20][14] ) );
  DFFR_X1 \pc_target_reg[20][16]  ( .D(n5849), .CK(Clk), .RN(n3881), .Q(
        \pc_target[20][16] ) );
  DFFR_X1 \pc_target_reg[20][18]  ( .D(n5848), .CK(Clk), .RN(n3881), .Q(
        \pc_target[20][18] ) );
  DFFR_X1 \pc_target_reg[20][20]  ( .D(n5847), .CK(Clk), .RN(n3881), .Q(
        \pc_target[20][20] ) );
  DFFR_X1 \pc_target_reg[20][22]  ( .D(n5846), .CK(Clk), .RN(n3881), .Q(
        \pc_target[20][22] ) );
  DFFR_X1 \pc_target_reg[20][24]  ( .D(n5845), .CK(Clk), .RN(n3882), .Q(
        \pc_target[20][24] ) );
  DFFR_X1 \pc_target_reg[20][26]  ( .D(n5844), .CK(Clk), .RN(n3882), .Q(
        \pc_target[20][26] ) );
  DFFR_X1 \pc_target_reg[20][28]  ( .D(n5843), .CK(Clk), .RN(n3882), .Q(
        \pc_target[20][28] ) );
  DFFR_X1 \pc_target_reg[20][30]  ( .D(n5842), .CK(Clk), .RN(n3882), .Q(
        \pc_target[20][30] ) );
  DFFR_X1 \pc_target_reg[21][31]  ( .D(n5841), .CK(Clk), .RN(n3864), .Q(
        \pc_target[21][31] ) );
  DFFR_X1 \pc_target_reg[21][29]  ( .D(n5840), .CK(Clk), .RN(n3882), .Q(
        \pc_target[21][29] ) );
  DFFR_X1 \pc_target_reg[21][27]  ( .D(n5839), .CK(Clk), .RN(n3882), .Q(
        \pc_target[21][27] ) );
  DFFR_X1 \pc_target_reg[21][25]  ( .D(n5838), .CK(Clk), .RN(n3882), .Q(
        \pc_target[21][25] ) );
  DFFR_X1 \pc_target_reg[21][23]  ( .D(n5837), .CK(Clk), .RN(n3882), .Q(
        \pc_target[21][23] ) );
  DFFR_X1 \pc_target_reg[21][21]  ( .D(n5836), .CK(Clk), .RN(n3882), .Q(
        \pc_target[21][21] ) );
  DFFR_X1 \pc_target_reg[21][19]  ( .D(n5835), .CK(Clk), .RN(n3882), .Q(
        \pc_target[21][19] ) );
  DFFR_X1 \pc_target_reg[21][17]  ( .D(n5834), .CK(Clk), .RN(n3882), .Q(
        \pc_target[21][17] ) );
  DFFR_X1 \pc_target_reg[21][15]  ( .D(n5833), .CK(Clk), .RN(n3882), .Q(
        \pc_target[21][15] ) );
  DFFR_X1 \pc_target_reg[21][13]  ( .D(n5832), .CK(Clk), .RN(n3882), .Q(
        \pc_target[21][13] ) );
  DFFR_X1 \pc_target_reg[21][11]  ( .D(n5831), .CK(Clk), .RN(n3882), .Q(
        \pc_target[21][11] ) );
  DFFR_X1 \pc_target_reg[21][7]  ( .D(n5829), .CK(Clk), .RN(n3882), .Q(
        \pc_target[21][7] ) );
  DFFR_X1 \pc_target_reg[21][3]  ( .D(n5827), .CK(Clk), .RN(n3883), .Q(
        \pc_target[21][3] ) );
  DFFR_X1 \pc_target_reg[21][1]  ( .D(n5826), .CK(Clk), .RN(n3883), .Q(
        \pc_target[21][1] ) );
  DFFR_X1 \pc_target_reg[21][0]  ( .D(n5825), .CK(Clk), .RN(n3883), .Q(
        \pc_target[21][0] ) );
  DFFR_X1 \pc_target_reg[21][2]  ( .D(n5824), .CK(Clk), .RN(n3883), .Q(
        \pc_target[21][2] ) );
  DFFR_X1 \pc_target_reg[21][12]  ( .D(n5819), .CK(Clk), .RN(n3883), .Q(
        \pc_target[21][12] ) );
  DFFR_X1 \pc_target_reg[21][14]  ( .D(n5818), .CK(Clk), .RN(n3883), .Q(
        \pc_target[21][14] ) );
  DFFR_X1 \pc_target_reg[21][16]  ( .D(n5817), .CK(Clk), .RN(n3883), .Q(
        \pc_target[21][16] ) );
  DFFR_X1 \pc_target_reg[21][18]  ( .D(n5816), .CK(Clk), .RN(n3883), .Q(
        \pc_target[21][18] ) );
  DFFR_X1 \pc_target_reg[21][20]  ( .D(n5815), .CK(Clk), .RN(n3883), .Q(
        \pc_target[21][20] ) );
  DFFR_X1 \pc_target_reg[21][22]  ( .D(n5814), .CK(Clk), .RN(n3883), .Q(
        \pc_target[21][22] ) );
  DFFR_X1 \pc_target_reg[21][24]  ( .D(n5813), .CK(Clk), .RN(n3883), .Q(
        \pc_target[21][24] ) );
  DFFR_X1 \pc_target_reg[21][26]  ( .D(n5812), .CK(Clk), .RN(n3883), .Q(
        \pc_target[21][26] ) );
  DFFR_X1 \pc_target_reg[21][28]  ( .D(n5811), .CK(Clk), .RN(n3883), .Q(
        \pc_target[21][28] ) );
  DFFR_X1 \pc_target_reg[21][30]  ( .D(n5810), .CK(Clk), .RN(n3883), .Q(
        \pc_target[21][30] ) );
  DFFR_X1 \pc_target_reg[22][31]  ( .D(n5809), .CK(Clk), .RN(n3865), .QN(n385)
         );
  DFFR_X1 \pc_target_reg[22][29]  ( .D(n5808), .CK(Clk), .RN(n3883), .QN(n384)
         );
  DFFR_X1 \pc_target_reg[22][27]  ( .D(n5807), .CK(Clk), .RN(n3884), .QN(n383)
         );
  DFFR_X1 \pc_target_reg[22][25]  ( .D(n5806), .CK(Clk), .RN(n3884), .QN(n382)
         );
  DFFR_X1 \pc_target_reg[22][23]  ( .D(n5805), .CK(Clk), .RN(n3884), .QN(n381)
         );
  DFFR_X1 \pc_target_reg[22][21]  ( .D(n5804), .CK(Clk), .RN(n3884), .QN(n380)
         );
  DFFR_X1 \pc_target_reg[22][19]  ( .D(n5803), .CK(Clk), .RN(n3884), .QN(n379)
         );
  DFFR_X1 \pc_target_reg[22][17]  ( .D(n5802), .CK(Clk), .RN(n3884), .QN(n378)
         );
  DFFR_X1 \pc_target_reg[22][15]  ( .D(n5801), .CK(Clk), .RN(n3884), .QN(n377)
         );
  DFFR_X1 \pc_target_reg[22][13]  ( .D(n5800), .CK(Clk), .RN(n3884), .QN(n376)
         );
  DFFR_X1 \pc_target_reg[22][11]  ( .D(n5799), .CK(Clk), .RN(n3884), .QN(n375)
         );
  DFFR_X1 \pc_target_reg[22][9]  ( .D(n5798), .CK(Clk), .RN(n3884), .QN(n374)
         );
  DFFR_X1 \pc_target_reg[22][7]  ( .D(n5797), .CK(Clk), .RN(n3884), .QN(n373)
         );
  DFFR_X1 \pc_target_reg[22][5]  ( .D(n5796), .CK(Clk), .RN(n3884), .QN(n372)
         );
  DFFR_X1 \pc_target_reg[22][3]  ( .D(n5795), .CK(Clk), .RN(n3884), .QN(n371)
         );
  DFFR_X1 \pc_target_reg[22][1]  ( .D(n5794), .CK(Clk), .RN(n3884), .QN(n370)
         );
  DFFR_X1 \pc_target_reg[22][0]  ( .D(n5793), .CK(Clk), .RN(n3885), .QN(n369)
         );
  DFFR_X1 \pc_target_reg[22][2]  ( .D(n5792), .CK(Clk), .RN(n3885), .QN(n368)
         );
  DFFR_X1 \pc_target_reg[22][4]  ( .D(n5791), .CK(Clk), .RN(n3885), .QN(n367)
         );
  DFFR_X1 \pc_target_reg[22][6]  ( .D(n5790), .CK(Clk), .RN(n3885), .QN(n366)
         );
  DFFR_X1 \pc_target_reg[22][8]  ( .D(n5789), .CK(Clk), .RN(n3885), .QN(n365)
         );
  DFFR_X1 \pc_target_reg[22][10]  ( .D(n5788), .CK(Clk), .RN(n3885), .QN(n364)
         );
  DFFR_X1 \pc_target_reg[22][12]  ( .D(n5787), .CK(Clk), .RN(n3885), .QN(n363)
         );
  DFFR_X1 \pc_target_reg[22][14]  ( .D(n5786), .CK(Clk), .RN(n3885), .QN(n362)
         );
  DFFR_X1 \pc_target_reg[22][16]  ( .D(n5785), .CK(Clk), .RN(n3885), .QN(n361)
         );
  DFFR_X1 \pc_target_reg[22][18]  ( .D(n5784), .CK(Clk), .RN(n3885), .QN(n360)
         );
  DFFR_X1 \pc_target_reg[22][20]  ( .D(n5783), .CK(Clk), .RN(n3885), .QN(n359)
         );
  DFFR_X1 \pc_target_reg[22][22]  ( .D(n5782), .CK(Clk), .RN(n3885), .QN(n358)
         );
  DFFR_X1 \pc_target_reg[22][24]  ( .D(n5781), .CK(Clk), .RN(n3886), .QN(n357)
         );
  DFFR_X1 \pc_target_reg[22][26]  ( .D(n5780), .CK(Clk), .RN(n3886), .QN(n356)
         );
  DFFR_X1 \pc_target_reg[22][28]  ( .D(n5779), .CK(Clk), .RN(n3886), .QN(n355)
         );
  DFFR_X1 \pc_target_reg[23][31]  ( .D(n5777), .CK(Clk), .RN(n3865), .QN(n350)
         );
  DFFR_X1 \pc_target_reg[23][29]  ( .D(n5776), .CK(Clk), .RN(n3885), .QN(n349)
         );
  DFFR_X1 \pc_target_reg[23][27]  ( .D(n5775), .CK(Clk), .RN(n3885), .QN(n348)
         );
  DFFR_X1 \pc_target_reg[23][25]  ( .D(n5774), .CK(Clk), .RN(n3885), .QN(n347)
         );
  DFFR_X1 \pc_target_reg[23][23]  ( .D(n5773), .CK(Clk), .RN(n3886), .QN(n346)
         );
  DFFR_X1 \pc_target_reg[23][21]  ( .D(n5772), .CK(Clk), .RN(n3886), .QN(n345)
         );
  DFFR_X1 \pc_target_reg[23][19]  ( .D(n5771), .CK(Clk), .RN(n3886), .QN(n344)
         );
  DFFR_X1 \pc_target_reg[23][17]  ( .D(n5770), .CK(Clk), .RN(n3886), .QN(n343)
         );
  DFFR_X1 \pc_target_reg[23][15]  ( .D(n5769), .CK(Clk), .RN(n3886), .QN(n342)
         );
  DFFR_X1 \pc_target_reg[23][13]  ( .D(n5768), .CK(Clk), .RN(n3886), .QN(n341)
         );
  DFFR_X1 \pc_target_reg[23][11]  ( .D(n5767), .CK(Clk), .RN(n3886), .QN(n340)
         );
  DFFR_X1 \pc_target_reg[23][9]  ( .D(n5766), .CK(Clk), .RN(n3886), .QN(n339)
         );
  DFFR_X1 \pc_target_reg[23][7]  ( .D(n5765), .CK(Clk), .RN(n3886), .QN(n338)
         );
  DFFR_X1 \pc_target_reg[23][5]  ( .D(n5764), .CK(Clk), .RN(n3886), .QN(n337)
         );
  DFFR_X1 \pc_target_reg[23][3]  ( .D(n5763), .CK(Clk), .RN(n3886), .QN(n336)
         );
  DFFR_X1 \pc_target_reg[23][1]  ( .D(n5762), .CK(Clk), .RN(n3886), .QN(n335)
         );
  DFFR_X1 \pc_target_reg[23][0]  ( .D(n5761), .CK(Clk), .RN(n3887), .QN(n334)
         );
  DFFR_X1 \pc_target_reg[23][2]  ( .D(n5760), .CK(Clk), .RN(n3887), .QN(n333)
         );
  DFFR_X1 \pc_target_reg[23][4]  ( .D(n5759), .CK(Clk), .RN(n3887), .QN(n332)
         );
  DFFR_X1 \pc_target_reg[23][6]  ( .D(n5758), .CK(Clk), .RN(n3887), .QN(n331)
         );
  DFFR_X1 \pc_target_reg[23][8]  ( .D(n5757), .CK(Clk), .RN(n3887), .QN(n330)
         );
  DFFR_X1 \pc_target_reg[23][10]  ( .D(n5756), .CK(Clk), .RN(n3887), .QN(n329)
         );
  DFFR_X1 \pc_target_reg[23][12]  ( .D(n5755), .CK(Clk), .RN(n3887), .QN(n328)
         );
  DFFR_X1 \pc_target_reg[23][14]  ( .D(n5754), .CK(Clk), .RN(n3887), .QN(n327)
         );
  DFFR_X1 \pc_target_reg[23][16]  ( .D(n5753), .CK(Clk), .RN(n3887), .QN(n326)
         );
  DFFR_X1 \pc_target_reg[23][18]  ( .D(n5752), .CK(Clk), .RN(n3887), .QN(n325)
         );
  DFFR_X1 \pc_target_reg[23][20]  ( .D(n5751), .CK(Clk), .RN(n3887), .QN(n324)
         );
  DFFR_X1 \pc_target_reg[23][22]  ( .D(n5750), .CK(Clk), .RN(n3887), .QN(n323)
         );
  DFFR_X1 \pc_target_reg[23][24]  ( .D(n5749), .CK(Clk), .RN(n3872), .QN(n322)
         );
  DFFR_X1 \pc_target_reg[23][26]  ( .D(n5748), .CK(Clk), .RN(n3872), .QN(n321)
         );
  DFFR_X1 \pc_target_reg[23][28]  ( .D(n5747), .CK(Clk), .RN(n3872), .QN(n320)
         );
  DFFR_X1 \pc_target_reg[24][31]  ( .D(n5745), .CK(Clk), .RN(n3865), .QN(n315)
         );
  DFFR_X1 \pc_target_reg[24][29]  ( .D(n5744), .CK(Clk), .RN(n3887), .QN(n314)
         );
  DFFR_X1 \pc_target_reg[24][27]  ( .D(n5743), .CK(Clk), .RN(n3887), .QN(n313)
         );
  DFFR_X1 \pc_target_reg[24][25]  ( .D(n5742), .CK(Clk), .RN(n3887), .QN(n312)
         );
  DFFR_X1 \pc_target_reg[24][23]  ( .D(n5741), .CK(Clk), .RN(n3888), .QN(n311)
         );
  DFFR_X1 \pc_target_reg[24][21]  ( .D(n5740), .CK(Clk), .RN(n3888), .QN(n310)
         );
  DFFR_X1 \pc_target_reg[24][19]  ( .D(n5739), .CK(Clk), .RN(n3888), .QN(n309)
         );
  DFFR_X1 \pc_target_reg[24][17]  ( .D(n5738), .CK(Clk), .RN(n3875), .QN(n308)
         );
  DFFR_X1 \pc_target_reg[24][15]  ( .D(n5737), .CK(Clk), .RN(n3871), .QN(n307)
         );
  DFFR_X1 \pc_target_reg[24][13]  ( .D(n5736), .CK(Clk), .RN(n3872), .QN(n306)
         );
  DFFR_X1 \pc_target_reg[24][11]  ( .D(n5735), .CK(Clk), .RN(n3872), .QN(n305)
         );
  DFFR_X1 \pc_target_reg[24][9]  ( .D(n5734), .CK(Clk), .RN(n3872), .QN(n304)
         );
  DFFR_X1 \pc_target_reg[24][7]  ( .D(n5733), .CK(Clk), .RN(n3872), .QN(n303)
         );
  DFFR_X1 \pc_target_reg[24][3]  ( .D(n5731), .CK(Clk), .RN(n3872), .QN(n301)
         );
  DFFR_X1 \pc_target_reg[24][1]  ( .D(n5730), .CK(Clk), .RN(n3872), .QN(n300)
         );
  DFFR_X1 \pc_target_reg[24][0]  ( .D(n5729), .CK(Clk), .RN(n3872), .QN(n299)
         );
  DFFR_X1 \pc_target_reg[24][2]  ( .D(n5728), .CK(Clk), .RN(n3872), .QN(n298)
         );
  DFFR_X1 \pc_target_reg[24][6]  ( .D(n5726), .CK(Clk), .RN(n3872), .QN(n296)
         );
  DFFR_X1 \pc_target_reg[24][8]  ( .D(n5725), .CK(Clk), .RN(n3872), .QN(n295)
         );
  DFFR_X1 \pc_target_reg[24][10]  ( .D(n5724), .CK(Clk), .RN(n3872), .QN(n294)
         );
  DFFR_X1 \pc_target_reg[24][12]  ( .D(n5723), .CK(Clk), .RN(n3873), .QN(n293)
         );
  DFFR_X1 \pc_target_reg[24][14]  ( .D(n5722), .CK(Clk), .RN(n3873), .QN(n292)
         );
  DFFR_X1 \pc_target_reg[24][16]  ( .D(n5721), .CK(Clk), .RN(n3873), .QN(n291)
         );
  DFFR_X1 \pc_target_reg[24][18]  ( .D(n5720), .CK(Clk), .RN(n3873), .QN(n290)
         );
  DFFR_X1 \pc_target_reg[24][20]  ( .D(n5719), .CK(Clk), .RN(n3873), .QN(n289)
         );
  DFFR_X1 \pc_target_reg[24][22]  ( .D(n5718), .CK(Clk), .RN(n3873), .QN(n288)
         );
  DFFR_X1 \pc_target_reg[24][24]  ( .D(n5717), .CK(Clk), .RN(n3873), .QN(n287)
         );
  DFFR_X1 \pc_target_reg[24][26]  ( .D(n5716), .CK(Clk), .RN(n3873), .QN(n286)
         );
  DFFR_X1 \pc_target_reg[24][28]  ( .D(n5715), .CK(Clk), .RN(n3873), .QN(n285)
         );
  DFFR_X1 \pc_target_reg[25][31]  ( .D(n5713), .CK(Clk), .RN(n3865), .QN(n281)
         );
  DFFR_X1 \pc_target_reg[25][29]  ( .D(n5712), .CK(Clk), .RN(n3872), .QN(n280)
         );
  DFFR_X1 \pc_target_reg[25][27]  ( .D(n5711), .CK(Clk), .RN(n3873), .QN(n279)
         );
  DFFR_X1 \pc_target_reg[25][25]  ( .D(n5710), .CK(Clk), .RN(n3873), .QN(n278)
         );
  DFFR_X1 \pc_target_reg[25][23]  ( .D(n5709), .CK(Clk), .RN(n3873), .QN(n277)
         );
  DFFR_X1 \pc_target_reg[25][21]  ( .D(n5708), .CK(Clk), .RN(n3873), .QN(n276)
         );
  DFFR_X1 \pc_target_reg[25][19]  ( .D(n5707), .CK(Clk), .RN(n3873), .QN(n275)
         );
  DFFR_X1 \pc_target_reg[25][17]  ( .D(n5706), .CK(Clk), .RN(n3873), .QN(n274)
         );
  DFFR_X1 \pc_target_reg[25][15]  ( .D(n5705), .CK(Clk), .RN(n3874), .QN(n273)
         );
  DFFR_X1 \pc_target_reg[25][13]  ( .D(n5704), .CK(Clk), .RN(n3874), .QN(n272)
         );
  DFFR_X1 \pc_target_reg[25][11]  ( .D(n5703), .CK(Clk), .RN(n3874), .QN(n271)
         );
  DFFR_X1 \pc_target_reg[25][9]  ( .D(n5702), .CK(Clk), .RN(n3874), .QN(n270)
         );
  DFFR_X1 \pc_target_reg[25][7]  ( .D(n5701), .CK(Clk), .RN(n3874), .QN(n269)
         );
  DFFR_X1 \pc_target_reg[25][5]  ( .D(n5700), .CK(Clk), .RN(n3874), .QN(n268)
         );
  DFFR_X1 \pc_target_reg[25][3]  ( .D(n5699), .CK(Clk), .RN(n3874), .QN(n267)
         );
  DFFR_X1 \pc_target_reg[25][1]  ( .D(n5698), .CK(Clk), .RN(n3874), .QN(n266)
         );
  DFFR_X1 \pc_target_reg[25][0]  ( .D(n5697), .CK(Clk), .RN(n3875), .QN(n265)
         );
  DFFR_X1 \pc_target_reg[25][2]  ( .D(n5696), .CK(Clk), .RN(n3874), .QN(n264)
         );
  DFFR_X1 \pc_target_reg[25][4]  ( .D(n5695), .CK(Clk), .RN(n3874), .QN(n263)
         );
  DFFR_X1 \pc_target_reg[25][6]  ( .D(n5694), .CK(Clk), .RN(n3874), .QN(n262)
         );
  DFFR_X1 \pc_target_reg[25][8]  ( .D(n5693), .CK(Clk), .RN(n3874), .QN(n261)
         );
  DFFR_X1 \pc_target_reg[25][10]  ( .D(n5692), .CK(Clk), .RN(n3874), .QN(n260)
         );
  DFFR_X1 \pc_target_reg[25][12]  ( .D(n5691), .CK(Clk), .RN(n3874), .QN(n259)
         );
  DFFR_X1 \pc_target_reg[25][14]  ( .D(n5690), .CK(Clk), .RN(n3874), .QN(n258)
         );
  DFFR_X1 \pc_target_reg[25][16]  ( .D(n5689), .CK(Clk), .RN(n3875), .QN(n257)
         );
  DFFR_X1 \pc_target_reg[25][18]  ( .D(n5688), .CK(Clk), .RN(n3875), .QN(n256)
         );
  DFFR_X1 \pc_target_reg[25][20]  ( .D(n5687), .CK(Clk), .RN(n3875), .QN(n255)
         );
  DFFR_X1 \pc_target_reg[25][22]  ( .D(n5686), .CK(Clk), .RN(n3875), .QN(n254)
         );
  DFFR_X1 \pc_target_reg[25][24]  ( .D(n5685), .CK(Clk), .RN(n3875), .QN(n253)
         );
  DFFR_X1 \pc_target_reg[25][26]  ( .D(n5684), .CK(Clk), .RN(n3875), .QN(n252)
         );
  DFFR_X1 \pc_target_reg[25][28]  ( .D(n5683), .CK(Clk), .RN(n3875), .QN(n251)
         );
  DFFR_X1 \pc_target_reg[26][31]  ( .D(n5681), .CK(Clk), .RN(n3871), .Q(
        \pc_target[26][31] ) );
  DFFR_X1 \pc_target_reg[26][29]  ( .D(n5680), .CK(Clk), .RN(n3875), .Q(
        \pc_target[26][29] ) );
  DFFR_X1 \pc_target_reg[26][27]  ( .D(n5679), .CK(Clk), .RN(n3875), .Q(
        \pc_target[26][27] ) );
  DFFR_X1 \pc_target_reg[26][25]  ( .D(n5678), .CK(Clk), .RN(n3875), .Q(
        \pc_target[26][25] ) );
  DFFR_X1 \pc_target_reg[26][23]  ( .D(n5677), .CK(Clk), .RN(n3875), .Q(
        \pc_target[26][23] ) );
  DFFR_X1 \pc_target_reg[26][21]  ( .D(n5676), .CK(Clk), .RN(n3875), .Q(
        \pc_target[26][21] ) );
  DFFR_X1 \pc_target_reg[26][19]  ( .D(n5675), .CK(Clk), .RN(n3875), .Q(
        \pc_target[26][19] ) );
  DFFR_X1 \pc_target_reg[26][17]  ( .D(n5674), .CK(Clk), .RN(n3876), .Q(
        \pc_target[26][17] ) );
  DFFR_X1 \pc_target_reg[26][15]  ( .D(n5673), .CK(Clk), .RN(n3876), .Q(
        \pc_target[26][15] ) );
  DFFR_X1 \pc_target_reg[26][13]  ( .D(n5672), .CK(Clk), .RN(n3876), .Q(
        \pc_target[26][13] ) );
  DFFR_X1 \pc_target_reg[26][11]  ( .D(n5671), .CK(Clk), .RN(n3876), .Q(
        \pc_target[26][11] ) );
  DFFR_X1 \pc_target_reg[26][9]  ( .D(n5670), .CK(Clk), .RN(n3876), .Q(
        \pc_target[26][9] ) );
  DFFR_X1 \pc_target_reg[26][7]  ( .D(n5669), .CK(Clk), .RN(n3876), .Q(
        \pc_target[26][7] ) );
  DFFR_X1 \pc_target_reg[26][5]  ( .D(n5668), .CK(Clk), .RN(n3876), .Q(
        \pc_target[26][5] ) );
  DFFR_X1 \pc_target_reg[26][3]  ( .D(n5667), .CK(Clk), .RN(n3876), .Q(
        \pc_target[26][3] ) );
  DFFR_X1 \pc_target_reg[26][1]  ( .D(n5666), .CK(Clk), .RN(n3876), .Q(
        \pc_target[26][1] ) );
  DFFR_X1 \pc_target_reg[26][0]  ( .D(n5665), .CK(Clk), .RN(n3876), .Q(
        \pc_target[26][0] ) );
  DFFR_X1 \pc_target_reg[26][2]  ( .D(n5664), .CK(Clk), .RN(n3876), .Q(
        \pc_target[26][2] ) );
  DFFR_X1 \pc_target_reg[26][4]  ( .D(n5663), .CK(Clk), .RN(n3876), .Q(
        \pc_target[26][4] ) );
  DFFR_X1 \pc_target_reg[26][6]  ( .D(n5662), .CK(Clk), .RN(n3876), .Q(
        \pc_target[26][6] ) );
  DFFR_X1 \pc_target_reg[26][8]  ( .D(n5661), .CK(Clk), .RN(n3876), .Q(
        \pc_target[26][8] ) );
  DFFR_X1 \pc_target_reg[26][10]  ( .D(n5660), .CK(Clk), .RN(n3876), .Q(
        \pc_target[26][10] ) );
  DFFR_X1 \pc_target_reg[26][12]  ( .D(n5659), .CK(Clk), .RN(n3877), .Q(
        \pc_target[26][12] ) );
  DFFR_X1 \pc_target_reg[26][14]  ( .D(n5658), .CK(Clk), .RN(n3877), .Q(
        \pc_target[26][14] ) );
  DFFR_X1 \pc_target_reg[26][16]  ( .D(n5657), .CK(Clk), .RN(n3877), .Q(
        \pc_target[26][16] ) );
  DFFR_X1 \pc_target_reg[26][18]  ( .D(n5656), .CK(Clk), .RN(n3877), .Q(
        \pc_target[26][18] ) );
  DFFR_X1 \pc_target_reg[26][20]  ( .D(n5655), .CK(Clk), .RN(n3877), .Q(
        \pc_target[26][20] ) );
  DFFR_X1 \pc_target_reg[26][22]  ( .D(n5654), .CK(Clk), .RN(n3877), .Q(
        \pc_target[26][22] ) );
  DFFR_X1 \pc_target_reg[26][24]  ( .D(n5653), .CK(Clk), .RN(n3877), .Q(
        \pc_target[26][24] ) );
  DFFR_X1 \pc_target_reg[26][26]  ( .D(n5652), .CK(Clk), .RN(n3877), .Q(
        \pc_target[26][26] ) );
  DFFR_X1 \pc_target_reg[26][28]  ( .D(n5651), .CK(Clk), .RN(n3877), .Q(
        \pc_target[26][28] ) );
  DFFR_X1 \pc_target_reg[26][30]  ( .D(n5650), .CK(Clk), .RN(n3866), .Q(
        \pc_target[26][30] ) );
  DFFR_X1 \pc_target_reg[27][31]  ( .D(n5649), .CK(Clk), .RN(n3888), .Q(
        \pc_target[27][31] ) );
  DFFR_X1 \pc_target_reg[27][29]  ( .D(n5648), .CK(Clk), .RN(n3865), .Q(
        \pc_target[27][29] ) );
  DFFR_X1 \pc_target_reg[27][27]  ( .D(n5647), .CK(Clk), .RN(n3865), .Q(
        \pc_target[27][27] ) );
  DFFR_X1 \pc_target_reg[27][25]  ( .D(n5646), .CK(Clk), .RN(n3866), .Q(
        \pc_target[27][25] ) );
  DFFR_X1 \pc_target_reg[27][23]  ( .D(n5645), .CK(Clk), .RN(n3866), .Q(
        \pc_target[27][23] ) );
  DFFR_X1 \pc_target_reg[27][21]  ( .D(n5644), .CK(Clk), .RN(n3866), .Q(
        \pc_target[27][21] ) );
  DFFR_X1 \pc_target_reg[27][19]  ( .D(n5643), .CK(Clk), .RN(n3866), .Q(
        \pc_target[27][19] ) );
  DFFR_X1 \pc_target_reg[27][17]  ( .D(n5642), .CK(Clk), .RN(n3866), .Q(
        \pc_target[27][17] ) );
  DFFR_X1 \pc_target_reg[27][15]  ( .D(n5641), .CK(Clk), .RN(n3866), .Q(
        \pc_target[27][15] ) );
  DFFR_X1 \pc_target_reg[27][13]  ( .D(n5640), .CK(Clk), .RN(n3866), .Q(
        \pc_target[27][13] ) );
  DFFR_X1 \pc_target_reg[27][11]  ( .D(n5639), .CK(Clk), .RN(n3866), .Q(
        \pc_target[27][11] ) );
  DFFR_X1 \pc_target_reg[27][9]  ( .D(n5638), .CK(Clk), .RN(n3866), .Q(
        \pc_target[27][9] ) );
  DFFR_X1 \pc_target_reg[27][7]  ( .D(n5637), .CK(Clk), .RN(n3866), .Q(
        \pc_target[27][7] ) );
  DFFR_X1 \pc_target_reg[27][5]  ( .D(n5636), .CK(Clk), .RN(n3866), .Q(
        \pc_target[27][5] ) );
  DFFR_X1 \pc_target_reg[27][3]  ( .D(n5635), .CK(Clk), .RN(n3866), .Q(
        \pc_target[27][3] ) );
  DFFR_X1 \pc_target_reg[27][1]  ( .D(n5634), .CK(Clk), .RN(n3866), .Q(
        \pc_target[27][1] ) );
  DFFR_X1 \pc_target_reg[27][0]  ( .D(n5633), .CK(Clk), .RN(n3867), .Q(
        \pc_target[27][0] ) );
  DFFR_X1 \pc_target_reg[27][2]  ( .D(n5632), .CK(Clk), .RN(n3866), .Q(
        \pc_target[27][2] ) );
  DFFR_X1 \pc_target_reg[27][4]  ( .D(n5631), .CK(Clk), .RN(n3867), .Q(
        \pc_target[27][4] ) );
  DFFR_X1 \pc_target_reg[27][6]  ( .D(n5630), .CK(Clk), .RN(n3867), .Q(
        \pc_target[27][6] ) );
  DFFR_X1 \pc_target_reg[27][8]  ( .D(n5629), .CK(Clk), .RN(n3867), .Q(
        \pc_target[27][8] ) );
  DFFR_X1 \pc_target_reg[27][10]  ( .D(n5628), .CK(Clk), .RN(n3867), .Q(
        \pc_target[27][10] ) );
  DFFR_X1 \pc_target_reg[27][12]  ( .D(n5627), .CK(Clk), .RN(n3867), .Q(
        \pc_target[27][12] ) );
  DFFR_X1 \pc_target_reg[27][14]  ( .D(n5626), .CK(Clk), .RN(n3867), .Q(
        \pc_target[27][14] ) );
  DFFR_X1 \pc_target_reg[27][16]  ( .D(n5625), .CK(Clk), .RN(n3867), .Q(
        \pc_target[27][16] ) );
  DFFR_X1 \pc_target_reg[27][18]  ( .D(n5624), .CK(Clk), .RN(n3867), .Q(
        \pc_target[27][18] ) );
  DFFR_X1 \pc_target_reg[27][20]  ( .D(n5623), .CK(Clk), .RN(n3867), .Q(
        \pc_target[27][20] ) );
  DFFR_X1 \pc_target_reg[27][22]  ( .D(n5622), .CK(Clk), .RN(n3867), .Q(
        \pc_target[27][22] ) );
  DFFR_X1 \pc_target_reg[27][24]  ( .D(n5621), .CK(Clk), .RN(n3867), .Q(
        \pc_target[27][24] ) );
  DFFR_X1 \pc_target_reg[27][26]  ( .D(n5620), .CK(Clk), .RN(n3867), .Q(
        \pc_target[27][26] ) );
  DFFR_X1 \pc_target_reg[27][28]  ( .D(n5619), .CK(Clk), .RN(n3867), .Q(
        \pc_target[27][28] ) );
  DFFR_X1 \pc_target_reg[27][30]  ( .D(n5618), .CK(Clk), .RN(n3868), .Q(
        \pc_target[27][30] ) );
  DFFR_X1 \pc_target_reg[28][31]  ( .D(n5617), .CK(Clk), .RN(n3865), .QN(n175)
         );
  DFFR_X1 \pc_target_reg[28][29]  ( .D(n5616), .CK(Clk), .RN(n3868), .QN(n174)
         );
  DFFR_X1 \pc_target_reg[28][27]  ( .D(n5615), .CK(Clk), .RN(n3868), .QN(n173)
         );
  DFFR_X1 \pc_target_reg[28][25]  ( .D(n5614), .CK(Clk), .RN(n3868), .QN(n172)
         );
  DFFR_X1 \pc_target_reg[28][23]  ( .D(n5613), .CK(Clk), .RN(n3868), .QN(n171)
         );
  DFFR_X1 \pc_target_reg[28][21]  ( .D(n5612), .CK(Clk), .RN(n3868), .QN(n170)
         );
  DFFR_X1 \pc_target_reg[28][19]  ( .D(n5611), .CK(Clk), .RN(n3868), .QN(n169)
         );
  DFFR_X1 \pc_target_reg[28][17]  ( .D(n5610), .CK(Clk), .RN(n3868), .QN(n168)
         );
  DFFR_X1 \pc_target_reg[28][15]  ( .D(n5609), .CK(Clk), .RN(n3868), .QN(n167)
         );
  DFFR_X1 \pc_target_reg[28][13]  ( .D(n5608), .CK(Clk), .RN(n3868), .QN(n166)
         );
  DFFR_X1 \pc_target_reg[28][11]  ( .D(n5607), .CK(Clk), .RN(n3868), .QN(n165)
         );
  DFFR_X1 \pc_target_reg[28][9]  ( .D(n5606), .CK(Clk), .RN(n3868), .QN(n164)
         );
  DFFR_X1 \pc_target_reg[28][7]  ( .D(n5605), .CK(Clk), .RN(n3868), .QN(n163)
         );
  DFFR_X1 \pc_target_reg[28][5]  ( .D(n5604), .CK(Clk), .RN(n3868), .QN(n162)
         );
  DFFR_X1 \pc_target_reg[28][3]  ( .D(n5603), .CK(Clk), .RN(n3868), .QN(n161)
         );
  DFFR_X1 \pc_target_reg[28][1]  ( .D(n5602), .CK(Clk), .RN(n3869), .QN(n160)
         );
  DFFR_X1 \pc_target_reg[28][0]  ( .D(n5601), .CK(Clk), .RN(n3869), .QN(n159)
         );
  DFFR_X1 \pc_target_reg[28][2]  ( .D(n5600), .CK(Clk), .RN(n3869), .QN(n158)
         );
  DFFR_X1 \pc_target_reg[28][4]  ( .D(n5599), .CK(Clk), .RN(n3869), .QN(n157)
         );
  DFFR_X1 \pc_target_reg[28][6]  ( .D(n5598), .CK(Clk), .RN(n3869), .QN(n156)
         );
  DFFR_X1 \pc_target_reg[28][8]  ( .D(n5597), .CK(Clk), .RN(n3869), .QN(n155)
         );
  DFFR_X1 \pc_target_reg[28][10]  ( .D(n5596), .CK(Clk), .RN(n3869), .QN(n154)
         );
  DFFR_X1 \pc_target_reg[28][12]  ( .D(n5595), .CK(Clk), .RN(n3869), .QN(n153)
         );
  DFFR_X1 \pc_target_reg[28][14]  ( .D(n5594), .CK(Clk), .RN(n3869), .QN(n152)
         );
  DFFR_X1 \pc_target_reg[28][16]  ( .D(n5593), .CK(Clk), .RN(n3869), .QN(n151)
         );
  DFFR_X1 \pc_target_reg[28][18]  ( .D(n5592), .CK(Clk), .RN(n3869), .QN(n150)
         );
  DFFR_X1 \pc_target_reg[28][20]  ( .D(n5591), .CK(Clk), .RN(n3869), .QN(n149)
         );
  DFFR_X1 \pc_target_reg[28][22]  ( .D(n5590), .CK(Clk), .RN(n3869), .QN(n148)
         );
  DFFR_X1 \pc_target_reg[28][24]  ( .D(n5589), .CK(Clk), .RN(n3869), .QN(n147)
         );
  DFFR_X1 \pc_target_reg[28][26]  ( .D(n5588), .CK(Clk), .RN(n3869), .QN(n146)
         );
  DFFR_X1 \pc_target_reg[28][28]  ( .D(n5587), .CK(Clk), .RN(n3870), .QN(n145)
         );
  DFFR_X1 \pc_target_reg[29][31]  ( .D(n5585), .CK(Clk), .RN(n3865), .QN(n140)
         );
  DFFR_X1 \pc_target_reg[29][29]  ( .D(n5584), .CK(Clk), .RN(n3870), .QN(n138)
         );
  DFFR_X1 \pc_target_reg[29][27]  ( .D(n5583), .CK(Clk), .RN(n3870), .QN(n136)
         );
  DFFR_X1 \pc_target_reg[29][25]  ( .D(n5582), .CK(Clk), .RN(n3870), .QN(n134)
         );
  DFFR_X1 \pc_target_reg[29][23]  ( .D(n5581), .CK(Clk), .RN(n3870), .QN(n132)
         );
  DFFR_X1 \pc_target_reg[29][21]  ( .D(n5580), .CK(Clk), .RN(n3870), .QN(n130)
         );
  DFFR_X1 \pc_target_reg[29][19]  ( .D(n5579), .CK(Clk), .RN(n3870), .QN(n128)
         );
  DFFR_X1 \pc_target_reg[29][17]  ( .D(n5578), .CK(Clk), .RN(n3870), .QN(n126)
         );
  DFFR_X1 \pc_target_reg[29][15]  ( .D(n5577), .CK(Clk), .RN(n3870), .QN(n124)
         );
  DFFR_X1 \pc_target_reg[29][13]  ( .D(n5576), .CK(Clk), .RN(n3870), .QN(n122)
         );
  DFFR_X1 \pc_target_reg[29][11]  ( .D(n5575), .CK(Clk), .RN(n3870), .QN(n120)
         );
  DFFR_X1 \pc_target_reg[29][9]  ( .D(n5574), .CK(Clk), .RN(n3870), .QN(n118)
         );
  DFFR_X1 \pc_target_reg[29][7]  ( .D(n5573), .CK(Clk), .RN(n3870), .QN(n116)
         );
  DFFR_X1 \pc_target_reg[29][5]  ( .D(n5572), .CK(Clk), .RN(n3870), .QN(n114)
         );
  DFFR_X1 \pc_target_reg[29][3]  ( .D(n5571), .CK(Clk), .RN(n3870), .QN(n112)
         );
  DFFR_X1 \pc_target_reg[29][1]  ( .D(n5570), .CK(Clk), .RN(n3871), .QN(n110)
         );
  DFFR_X1 \pc_target_reg[29][0]  ( .D(n5569), .CK(Clk), .RN(n3871), .QN(n108)
         );
  DFFR_X1 \pc_target_reg[29][2]  ( .D(n5568), .CK(Clk), .RN(n3871), .QN(n106)
         );
  DFFR_X1 \pc_target_reg[29][4]  ( .D(n5567), .CK(Clk), .RN(n3871), .QN(n104)
         );
  DFFR_X1 \pc_target_reg[29][6]  ( .D(n5566), .CK(Clk), .RN(n3871), .QN(n102)
         );
  DFFR_X1 \pc_target_reg[29][8]  ( .D(n5565), .CK(Clk), .RN(n3871), .QN(n100)
         );
  DFFR_X1 \pc_target_reg[29][10]  ( .D(n5564), .CK(Clk), .RN(n3871), .QN(n98)
         );
  DFFR_X1 \pc_target_reg[29][12]  ( .D(n5563), .CK(Clk), .RN(n3871), .QN(n96)
         );
  DFFR_X1 \pc_target_reg[29][14]  ( .D(n5562), .CK(Clk), .RN(n3871), .QN(n94)
         );
  DFFR_X1 \pc_target_reg[29][16]  ( .D(n5561), .CK(Clk), .RN(n3871), .QN(n92)
         );
  DFFR_X1 \pc_target_reg[29][18]  ( .D(n5560), .CK(Clk), .RN(n3871), .QN(n90)
         );
  DFFR_X1 \pc_target_reg[29][20]  ( .D(n5559), .CK(Clk), .RN(n3859), .QN(n88)
         );
  DFFR_X1 \pc_target_reg[29][22]  ( .D(n5558), .CK(Clk), .RN(n3855), .QN(n86)
         );
  DFFR_X1 \pc_target_reg[29][24]  ( .D(n5557), .CK(Clk), .RN(n3855), .QN(n84)
         );
  DFFR_X1 \pc_target_reg[29][26]  ( .D(n5556), .CK(Clk), .RN(n3855), .QN(n82)
         );
  DFFR_X1 \pc_target_reg[29][28]  ( .D(n5555), .CK(Clk), .RN(n3855), .QN(n80)
         );
  DFFR_X1 \pc_target_reg[30][31]  ( .D(n5553), .CK(Clk), .RN(n3867), .Q(
        \pc_target[30][31] ) );
  DFFR_X1 \pc_target_reg[30][29]  ( .D(n5552), .CK(Clk), .RN(n3871), .Q(
        \pc_target[30][29] ) );
  DFFR_X1 \pc_target_reg[30][27]  ( .D(n5551), .CK(Clk), .RN(n3871), .Q(
        \pc_target[30][27] ) );
  DFFR_X1 \pc_target_reg[30][25]  ( .D(n5550), .CK(Clk), .RN(n3855), .Q(
        \pc_target[30][25] ) );
  DFFR_X1 \pc_target_reg[30][23]  ( .D(n5549), .CK(Clk), .RN(n3856), .Q(
        \pc_target[30][23] ) );
  DFFR_X1 \pc_target_reg[30][21]  ( .D(n5548), .CK(Clk), .RN(n3856), .Q(
        \pc_target[30][21] ) );
  DFFR_X1 \pc_target_reg[30][19]  ( .D(n5547), .CK(Clk), .RN(n3856), .Q(
        \pc_target[30][19] ) );
  DFFR_X1 \pc_target_reg[30][17]  ( .D(n5546), .CK(Clk), .RN(n3856), .Q(
        \pc_target[30][17] ) );
  DFFR_X1 \pc_target_reg[30][15]  ( .D(n5545), .CK(Clk), .RN(n3856), .Q(
        \pc_target[30][15] ) );
  DFFR_X1 \pc_target_reg[30][13]  ( .D(n5544), .CK(Clk), .RN(n3856), .Q(
        \pc_target[30][13] ) );
  DFFR_X1 \pc_target_reg[30][11]  ( .D(n5543), .CK(Clk), .RN(n3856), .Q(
        \pc_target[30][11] ) );
  DFFR_X1 \pc_target_reg[30][9]  ( .D(n5542), .CK(Clk), .RN(n3856), .Q(
        \pc_target[30][9] ) );
  DFFR_X1 \pc_target_reg[30][7]  ( .D(n5541), .CK(Clk), .RN(n3856), .Q(
        \pc_target[30][7] ) );
  DFFR_X1 \pc_target_reg[30][5]  ( .D(n5540), .CK(Clk), .RN(n3856), .Q(
        \pc_target[30][5] ) );
  DFFR_X1 \pc_target_reg[30][3]  ( .D(n5539), .CK(Clk), .RN(n3856), .Q(
        \pc_target[30][3] ) );
  DFFR_X1 \pc_target_reg[30][1]  ( .D(n5538), .CK(Clk), .RN(n3856), .Q(
        \pc_target[30][1] ) );
  DFFR_X1 \pc_target_reg[30][0]  ( .D(n5537), .CK(Clk), .RN(n3857), .Q(
        \pc_target[30][0] ) );
  DFFR_X1 \pc_target_reg[30][2]  ( .D(n5536), .CK(Clk), .RN(n3856), .Q(
        \pc_target[30][2] ) );
  DFFR_X1 \pc_target_reg[30][4]  ( .D(n5535), .CK(Clk), .RN(n3856), .Q(
        \pc_target[30][4] ) );
  DFFR_X1 \pc_target_reg[30][6]  ( .D(n5534), .CK(Clk), .RN(n3856), .Q(
        \pc_target[30][6] ) );
  DFFR_X1 \pc_target_reg[30][8]  ( .D(n5533), .CK(Clk), .RN(n3857), .Q(
        \pc_target[30][8] ) );
  DFFR_X1 \pc_target_reg[30][10]  ( .D(n5532), .CK(Clk), .RN(n3857), .Q(
        \pc_target[30][10] ) );
  DFFR_X1 \pc_target_reg[30][12]  ( .D(n5531), .CK(Clk), .RN(n3857), .Q(
        \pc_target[30][12] ) );
  DFFR_X1 \pc_target_reg[30][14]  ( .D(n5530), .CK(Clk), .RN(n3857), .Q(
        \pc_target[30][14] ) );
  DFFR_X1 \pc_target_reg[30][16]  ( .D(n5529), .CK(Clk), .RN(n3857), .Q(
        \pc_target[30][16] ) );
  DFFR_X1 \pc_target_reg[30][18]  ( .D(n5528), .CK(Clk), .RN(n3857), .Q(
        \pc_target[30][18] ) );
  DFFR_X1 \pc_target_reg[30][20]  ( .D(n5527), .CK(Clk), .RN(n3857), .Q(
        \pc_target[30][20] ) );
  DFFR_X1 \pc_target_reg[30][22]  ( .D(n5526), .CK(Clk), .RN(n3857), .Q(
        \pc_target[30][22] ) );
  DFFR_X1 \pc_target_reg[30][24]  ( .D(n5525), .CK(Clk), .RN(n3857), .Q(
        \pc_target[30][24] ) );
  DFFR_X1 \pc_target_reg[30][26]  ( .D(n5524), .CK(Clk), .RN(n3857), .Q(
        \pc_target[30][26] ) );
  DFFR_X1 \pc_target_reg[30][28]  ( .D(n5523), .CK(Clk), .RN(n3857), .Q(
        \pc_target[30][28] ) );
  DFFR_X1 \pc_target_reg[30][30]  ( .D(n5522), .CK(Clk), .RN(n3857), .Q(
        \pc_target[30][30] ) );
  DFFR_X1 \pc_target_reg[31][31]  ( .D(n5521), .CK(Clk), .RN(n3863), .Q(
        \pc_target[31][31] ) );
  DLH_X1 \OUT_PC_target_reg[31]  ( .G(Enable), .D(N96), .Q(OUT_PC_target[31])
         );
  DFFR_X1 \pc_target_reg[31][29]  ( .D(n5520), .CK(Clk), .RN(n3857), .Q(
        \pc_target[31][29] ) );
  DLH_X1 \OUT_PC_target_reg[29]  ( .G(Enable), .D(N98), .Q(OUT_PC_target[29])
         );
  DFFR_X1 \pc_target_reg[31][27]  ( .D(n5519), .CK(Clk), .RN(n3857), .Q(
        \pc_target[31][27] ) );
  DLH_X1 \OUT_PC_target_reg[27]  ( .G(Enable), .D(N100), .Q(OUT_PC_target[27])
         );
  DFFR_X1 \pc_target_reg[31][25]  ( .D(n5518), .CK(Clk), .RN(n3858), .Q(
        \pc_target[31][25] ) );
  DLH_X1 \OUT_PC_target_reg[25]  ( .G(Enable), .D(N102), .Q(OUT_PC_target[25])
         );
  DFFR_X1 \pc_target_reg[31][23]  ( .D(n5517), .CK(Clk), .RN(n3858), .Q(
        \pc_target[31][23] ) );
  DLH_X1 \OUT_PC_target_reg[23]  ( .G(Enable), .D(N104), .Q(OUT_PC_target[23])
         );
  DFFR_X1 \pc_target_reg[31][21]  ( .D(n5516), .CK(Clk), .RN(n3858), .Q(
        \pc_target[31][21] ) );
  DLH_X1 \OUT_PC_target_reg[21]  ( .G(Enable), .D(N106), .Q(OUT_PC_target[21])
         );
  DFFR_X1 \pc_target_reg[31][19]  ( .D(n5515), .CK(Clk), .RN(n3858), .Q(
        \pc_target[31][19] ) );
  DLH_X1 \OUT_PC_target_reg[19]  ( .G(Enable), .D(N108), .Q(OUT_PC_target[19])
         );
  DFFR_X1 \pc_target_reg[31][17]  ( .D(n5514), .CK(Clk), .RN(n3858), .Q(
        \pc_target[31][17] ) );
  DLH_X1 \OUT_PC_target_reg[17]  ( .G(Enable), .D(N110), .Q(OUT_PC_target[17])
         );
  DFFR_X1 \pc_target_reg[31][15]  ( .D(n5513), .CK(Clk), .RN(n3858), .Q(
        \pc_target[31][15] ) );
  DLH_X1 \OUT_PC_target_reg[15]  ( .G(Enable), .D(N112), .Q(OUT_PC_target[15])
         );
  DFFR_X1 \pc_target_reg[31][13]  ( .D(n5512), .CK(Clk), .RN(n3858), .Q(
        \pc_target[31][13] ) );
  DLH_X1 \OUT_PC_target_reg[13]  ( .G(Enable), .D(N114), .Q(OUT_PC_target[13])
         );
  DFFR_X1 \pc_target_reg[31][11]  ( .D(n5511), .CK(Clk), .RN(n3858), .Q(
        \pc_target[31][11] ) );
  DLH_X1 \OUT_PC_target_reg[11]  ( .G(Enable), .D(N116), .Q(OUT_PC_target[11])
         );
  DFFR_X1 \pc_target_reg[31][9]  ( .D(n5510), .CK(Clk), .RN(n3858), .Q(
        \pc_target[31][9] ) );
  DLH_X1 \OUT_PC_target_reg[9]  ( .G(Enable), .D(N118), .Q(OUT_PC_target[9])
         );
  DFFR_X1 \pc_target_reg[31][7]  ( .D(n5509), .CK(Clk), .RN(n3858), .Q(
        \pc_target[31][7] ) );
  DLH_X1 \OUT_PC_target_reg[7]  ( .G(Enable), .D(N120), .Q(OUT_PC_target[7])
         );
  DFFR_X1 \pc_target_reg[31][5]  ( .D(n5508), .CK(Clk), .RN(n3858), .Q(
        \pc_target[31][5] ) );
  DLH_X1 \OUT_PC_target_reg[5]  ( .G(Enable), .D(N122), .Q(OUT_PC_target[5])
         );
  DFFR_X1 \pc_target_reg[31][3]  ( .D(n5507), .CK(Clk), .RN(n3860), .Q(
        \pc_target[31][3] ) );
  DLH_X1 \OUT_PC_target_reg[3]  ( .G(Enable), .D(N124), .Q(OUT_PC_target[3])
         );
  DFFR_X1 \pc_target_reg[31][1]  ( .D(n5506), .CK(Clk), .RN(n3860), .Q(
        \pc_target[31][1] ) );
  DLH_X1 \OUT_PC_target_reg[1]  ( .G(Enable), .D(N126), .Q(OUT_PC_target[1])
         );
  DFFR_X1 \pc_target_reg[31][0]  ( .D(n5505), .CK(Clk), .RN(n3861), .Q(
        \pc_target[31][0] ) );
  DLH_X1 \OUT_PC_target_reg[0]  ( .G(Enable), .D(N127), .Q(OUT_PC_target[0])
         );
  DFFR_X1 \pc_target_reg[31][2]  ( .D(n5504), .CK(Clk), .RN(n3860), .Q(
        \pc_target[31][2] ) );
  DLH_X1 \OUT_PC_target_reg[2]  ( .G(Enable), .D(N125), .Q(OUT_PC_target[2])
         );
  DFFR_X1 \pc_target_reg[31][4]  ( .D(n5503), .CK(Clk), .RN(n3861), .Q(
        \pc_target[31][4] ) );
  DLH_X1 \OUT_PC_target_reg[4]  ( .G(Enable), .D(N123), .Q(OUT_PC_target[4])
         );
  DFFR_X1 \pc_target_reg[31][6]  ( .D(n5502), .CK(Clk), .RN(n3861), .Q(
        \pc_target[31][6] ) );
  DLH_X1 \OUT_PC_target_reg[6]  ( .G(Enable), .D(N121), .Q(OUT_PC_target[6])
         );
  DFFR_X1 \pc_target_reg[31][8]  ( .D(n5501), .CK(Clk), .RN(n3861), .Q(
        \pc_target[31][8] ) );
  DLH_X1 \OUT_PC_target_reg[8]  ( .G(Enable), .D(N119), .Q(OUT_PC_target[8])
         );
  DFFR_X1 \pc_target_reg[31][10]  ( .D(n5500), .CK(Clk), .RN(n3861), .Q(
        \pc_target[31][10] ) );
  DLH_X1 \OUT_PC_target_reg[10]  ( .G(Enable), .D(N117), .Q(OUT_PC_target[10])
         );
  DFFR_X1 \pc_target_reg[31][12]  ( .D(n5499), .CK(Clk), .RN(n3861), .Q(
        \pc_target[31][12] ) );
  DLH_X1 \OUT_PC_target_reg[12]  ( .G(Enable), .D(N115), .Q(OUT_PC_target[12])
         );
  DFFR_X1 \pc_target_reg[31][14]  ( .D(n5498), .CK(Clk), .RN(n3861), .Q(
        \pc_target[31][14] ) );
  DLH_X1 \OUT_PC_target_reg[14]  ( .G(Enable), .D(N113), .Q(OUT_PC_target[14])
         );
  DFFR_X1 \pc_target_reg[31][16]  ( .D(n5497), .CK(Clk), .RN(n3861), .Q(
        \pc_target[31][16] ) );
  DLH_X1 \OUT_PC_target_reg[16]  ( .G(Enable), .D(N111), .Q(OUT_PC_target[16])
         );
  DFFR_X1 \pc_target_reg[31][18]  ( .D(n5496), .CK(Clk), .RN(n3861), .Q(
        \pc_target[31][18] ) );
  DLH_X1 \OUT_PC_target_reg[18]  ( .G(Enable), .D(N109), .Q(OUT_PC_target[18])
         );
  DFFR_X1 \pc_target_reg[31][20]  ( .D(n5495), .CK(Clk), .RN(n3863), .Q(
        \pc_target[31][20] ) );
  DLH_X1 \OUT_PC_target_reg[20]  ( .G(Enable), .D(N107), .Q(OUT_PC_target[20])
         );
  DFFR_X1 \pc_target_reg[31][22]  ( .D(n5494), .CK(Clk), .RN(n3863), .Q(
        \pc_target[31][22] ) );
  DLH_X1 \OUT_PC_target_reg[22]  ( .G(Enable), .D(N105), .Q(OUT_PC_target[22])
         );
  DFFR_X1 \pc_target_reg[31][24]  ( .D(n5493), .CK(Clk), .RN(n3863), .Q(
        \pc_target[31][24] ) );
  DLH_X1 \OUT_PC_target_reg[24]  ( .G(Enable), .D(N103), .Q(OUT_PC_target[24])
         );
  DFFR_X1 \pc_target_reg[31][26]  ( .D(n5492), .CK(Clk), .RN(n3863), .Q(
        \pc_target[31][26] ) );
  DLH_X1 \OUT_PC_target_reg[26]  ( .G(Enable), .D(N101), .Q(OUT_PC_target[26])
         );
  DFFR_X1 \pc_target_reg[31][28]  ( .D(n5491), .CK(Clk), .RN(n3864), .Q(
        \pc_target[31][28] ) );
  DLH_X1 \OUT_PC_target_reg[28]  ( .G(Enable), .D(N99), .Q(OUT_PC_target[28])
         );
  DFFR_X1 \pc_target_reg[31][30]  ( .D(n5490), .CK(Clk), .RN(n3864), .Q(
        \pc_target[31][30] ) );
  DLH_X1 \OUT_PC_target_reg[30]  ( .G(Enable), .D(N97), .Q(OUT_PC_target[30])
         );
  INV_X1 U3 ( .A(n4), .ZN(n5490) );
  AOI22_X1 U5 ( .A1(n5), .A2(Set_target[30]), .B1(n6), .B2(\pc_target[31][30] ), .ZN(n4) );
  INV_X1 U6 ( .A(n7), .ZN(n5491) );
  AOI22_X1 U7 ( .A1(n5), .A2(Set_target[28]), .B1(n6), .B2(\pc_target[31][28] ), .ZN(n7) );
  INV_X1 U8 ( .A(n8), .ZN(n5492) );
  AOI22_X1 U9 ( .A1(n5), .A2(Set_target[26]), .B1(n6), .B2(\pc_target[31][26] ), .ZN(n8) );
  INV_X1 U10 ( .A(n9), .ZN(n5493) );
  AOI22_X1 U11 ( .A1(n5), .A2(Set_target[24]), .B1(n6), .B2(
        \pc_target[31][24] ), .ZN(n9) );
  INV_X1 U12 ( .A(n10), .ZN(n5494) );
  AOI22_X1 U13 ( .A1(n5), .A2(Set_target[22]), .B1(n6), .B2(
        \pc_target[31][22] ), .ZN(n10) );
  INV_X1 U14 ( .A(n11), .ZN(n5495) );
  AOI22_X1 U15 ( .A1(n5), .A2(Set_target[20]), .B1(n6), .B2(
        \pc_target[31][20] ), .ZN(n11) );
  INV_X1 U16 ( .A(n12), .ZN(n5496) );
  AOI22_X1 U17 ( .A1(n5), .A2(Set_target[18]), .B1(n6), .B2(
        \pc_target[31][18] ), .ZN(n12) );
  INV_X1 U18 ( .A(n13), .ZN(n5497) );
  AOI22_X1 U19 ( .A1(n5), .A2(Set_target[16]), .B1(n6), .B2(
        \pc_target[31][16] ), .ZN(n13) );
  INV_X1 U20 ( .A(n14), .ZN(n5498) );
  AOI22_X1 U21 ( .A1(n5), .A2(Set_target[14]), .B1(n6), .B2(
        \pc_target[31][14] ), .ZN(n14) );
  INV_X1 U22 ( .A(n15), .ZN(n5499) );
  AOI22_X1 U23 ( .A1(n5), .A2(Set_target[12]), .B1(n6), .B2(
        \pc_target[31][12] ), .ZN(n15) );
  INV_X1 U24 ( .A(n16), .ZN(n5500) );
  AOI22_X1 U25 ( .A1(n5), .A2(Set_target[10]), .B1(n6), .B2(
        \pc_target[31][10] ), .ZN(n16) );
  INV_X1 U26 ( .A(n17), .ZN(n5501) );
  AOI22_X1 U27 ( .A1(n5), .A2(Set_target[8]), .B1(n6), .B2(\pc_target[31][8] ), 
        .ZN(n17) );
  INV_X1 U28 ( .A(n18), .ZN(n5502) );
  AOI22_X1 U29 ( .A1(n5), .A2(Set_target[6]), .B1(n6), .B2(\pc_target[31][6] ), 
        .ZN(n18) );
  INV_X1 U30 ( .A(n19), .ZN(n5503) );
  AOI22_X1 U31 ( .A1(n5), .A2(Set_target[4]), .B1(n6), .B2(\pc_target[31][4] ), 
        .ZN(n19) );
  INV_X1 U32 ( .A(n20), .ZN(n5504) );
  AOI22_X1 U33 ( .A1(n5), .A2(Set_target[2]), .B1(n6), .B2(\pc_target[31][2] ), 
        .ZN(n20) );
  INV_X1 U34 ( .A(n21), .ZN(n5505) );
  AOI22_X1 U35 ( .A1(n5), .A2(Set_target[0]), .B1(n6), .B2(\pc_target[31][0] ), 
        .ZN(n21) );
  INV_X1 U36 ( .A(n22), .ZN(n5506) );
  AOI22_X1 U37 ( .A1(n5), .A2(Set_target[1]), .B1(n6), .B2(\pc_target[31][1] ), 
        .ZN(n22) );
  INV_X1 U38 ( .A(n23), .ZN(n5507) );
  AOI22_X1 U39 ( .A1(n5), .A2(Set_target[3]), .B1(n6), .B2(\pc_target[31][3] ), 
        .ZN(n23) );
  INV_X1 U40 ( .A(n24), .ZN(n5508) );
  AOI22_X1 U41 ( .A1(n5), .A2(Set_target[5]), .B1(n6), .B2(\pc_target[31][5] ), 
        .ZN(n24) );
  INV_X1 U42 ( .A(n25), .ZN(n5509) );
  AOI22_X1 U43 ( .A1(n5), .A2(Set_target[7]), .B1(n6), .B2(\pc_target[31][7] ), 
        .ZN(n25) );
  INV_X1 U44 ( .A(n26), .ZN(n5510) );
  AOI22_X1 U45 ( .A1(n5), .A2(Set_target[9]), .B1(n6), .B2(\pc_target[31][9] ), 
        .ZN(n26) );
  INV_X1 U46 ( .A(n27), .ZN(n5511) );
  AOI22_X1 U47 ( .A1(n5), .A2(Set_target[11]), .B1(n6), .B2(
        \pc_target[31][11] ), .ZN(n27) );
  INV_X1 U48 ( .A(n28), .ZN(n5512) );
  AOI22_X1 U49 ( .A1(n5), .A2(Set_target[13]), .B1(n6), .B2(
        \pc_target[31][13] ), .ZN(n28) );
  INV_X1 U50 ( .A(n29), .ZN(n5513) );
  AOI22_X1 U51 ( .A1(n5), .A2(Set_target[15]), .B1(n6), .B2(
        \pc_target[31][15] ), .ZN(n29) );
  INV_X1 U52 ( .A(n30), .ZN(n5514) );
  AOI22_X1 U53 ( .A1(n5), .A2(Set_target[17]), .B1(n6), .B2(
        \pc_target[31][17] ), .ZN(n30) );
  INV_X1 U54 ( .A(n31), .ZN(n5515) );
  AOI22_X1 U55 ( .A1(n5), .A2(Set_target[19]), .B1(n6), .B2(
        \pc_target[31][19] ), .ZN(n31) );
  INV_X1 U56 ( .A(n32), .ZN(n5516) );
  AOI22_X1 U57 ( .A1(n5), .A2(Set_target[21]), .B1(n6), .B2(
        \pc_target[31][21] ), .ZN(n32) );
  INV_X1 U58 ( .A(n33), .ZN(n5517) );
  AOI22_X1 U59 ( .A1(n5), .A2(Set_target[23]), .B1(n6), .B2(
        \pc_target[31][23] ), .ZN(n33) );
  INV_X1 U60 ( .A(n34), .ZN(n5518) );
  AOI22_X1 U61 ( .A1(n5), .A2(Set_target[25]), .B1(n6), .B2(
        \pc_target[31][25] ), .ZN(n34) );
  INV_X1 U62 ( .A(n35), .ZN(n5519) );
  AOI22_X1 U63 ( .A1(n5), .A2(Set_target[27]), .B1(n6), .B2(
        \pc_target[31][27] ), .ZN(n35) );
  INV_X1 U64 ( .A(n36), .ZN(n5520) );
  AOI22_X1 U65 ( .A1(n5), .A2(Set_target[29]), .B1(n6), .B2(
        \pc_target[31][29] ), .ZN(n36) );
  INV_X1 U66 ( .A(n37), .ZN(n5521) );
  AOI22_X1 U67 ( .A1(n5), .A2(Set_target[31]), .B1(n6), .B2(
        \pc_target[31][31] ), .ZN(n37) );
  INV_X1 U70 ( .A(n40), .ZN(n5522) );
  AOI22_X1 U71 ( .A1(Set_target[30]), .A2(n3798), .B1(n42), .B2(
        \pc_target[30][30] ), .ZN(n40) );
  INV_X1 U72 ( .A(n43), .ZN(n5523) );
  AOI22_X1 U73 ( .A1(Set_target[28]), .A2(n3798), .B1(n42), .B2(
        \pc_target[30][28] ), .ZN(n43) );
  INV_X1 U74 ( .A(n44), .ZN(n5524) );
  AOI22_X1 U75 ( .A1(Set_target[26]), .A2(n3798), .B1(n42), .B2(
        \pc_target[30][26] ), .ZN(n44) );
  INV_X1 U76 ( .A(n45), .ZN(n5525) );
  AOI22_X1 U77 ( .A1(Set_target[24]), .A2(n3798), .B1(n42), .B2(
        \pc_target[30][24] ), .ZN(n45) );
  INV_X1 U78 ( .A(n46), .ZN(n5526) );
  AOI22_X1 U79 ( .A1(Set_target[22]), .A2(n3798), .B1(n42), .B2(
        \pc_target[30][22] ), .ZN(n46) );
  INV_X1 U80 ( .A(n47), .ZN(n5527) );
  AOI22_X1 U81 ( .A1(Set_target[20]), .A2(n3798), .B1(n42), .B2(
        \pc_target[30][20] ), .ZN(n47) );
  INV_X1 U82 ( .A(n48), .ZN(n5528) );
  AOI22_X1 U83 ( .A1(Set_target[18]), .A2(n3798), .B1(n42), .B2(
        \pc_target[30][18] ), .ZN(n48) );
  INV_X1 U84 ( .A(n49), .ZN(n5529) );
  AOI22_X1 U85 ( .A1(Set_target[16]), .A2(n3798), .B1(n42), .B2(
        \pc_target[30][16] ), .ZN(n49) );
  INV_X1 U86 ( .A(n50), .ZN(n5530) );
  AOI22_X1 U87 ( .A1(Set_target[14]), .A2(n3798), .B1(n42), .B2(
        \pc_target[30][14] ), .ZN(n50) );
  INV_X1 U88 ( .A(n51), .ZN(n5531) );
  AOI22_X1 U89 ( .A1(Set_target[12]), .A2(n3798), .B1(n42), .B2(
        \pc_target[30][12] ), .ZN(n51) );
  INV_X1 U90 ( .A(n52), .ZN(n5532) );
  AOI22_X1 U91 ( .A1(Set_target[10]), .A2(n3798), .B1(n42), .B2(
        \pc_target[30][10] ), .ZN(n52) );
  INV_X1 U92 ( .A(n53), .ZN(n5533) );
  AOI22_X1 U93 ( .A1(Set_target[8]), .A2(n3798), .B1(n42), .B2(
        \pc_target[30][8] ), .ZN(n53) );
  INV_X1 U94 ( .A(n54), .ZN(n5534) );
  AOI22_X1 U95 ( .A1(Set_target[6]), .A2(n3798), .B1(n42), .B2(
        \pc_target[30][6] ), .ZN(n54) );
  INV_X1 U96 ( .A(n55), .ZN(n5535) );
  AOI22_X1 U97 ( .A1(Set_target[4]), .A2(n3798), .B1(n42), .B2(
        \pc_target[30][4] ), .ZN(n55) );
  INV_X1 U98 ( .A(n56), .ZN(n5536) );
  AOI22_X1 U99 ( .A1(Set_target[2]), .A2(n3798), .B1(n42), .B2(
        \pc_target[30][2] ), .ZN(n56) );
  INV_X1 U100 ( .A(n57), .ZN(n5537) );
  AOI22_X1 U101 ( .A1(Set_target[0]), .A2(n3798), .B1(n42), .B2(
        \pc_target[30][0] ), .ZN(n57) );
  INV_X1 U102 ( .A(n58), .ZN(n5538) );
  AOI22_X1 U103 ( .A1(Set_target[1]), .A2(n3798), .B1(n42), .B2(
        \pc_target[30][1] ), .ZN(n58) );
  INV_X1 U104 ( .A(n59), .ZN(n5539) );
  AOI22_X1 U105 ( .A1(Set_target[3]), .A2(n3798), .B1(n42), .B2(
        \pc_target[30][3] ), .ZN(n59) );
  INV_X1 U106 ( .A(n60), .ZN(n5540) );
  AOI22_X1 U107 ( .A1(Set_target[5]), .A2(n3798), .B1(n42), .B2(
        \pc_target[30][5] ), .ZN(n60) );
  INV_X1 U108 ( .A(n61), .ZN(n5541) );
  AOI22_X1 U109 ( .A1(Set_target[7]), .A2(n3798), .B1(n42), .B2(
        \pc_target[30][7] ), .ZN(n61) );
  INV_X1 U110 ( .A(n62), .ZN(n5542) );
  AOI22_X1 U111 ( .A1(Set_target[9]), .A2(n3798), .B1(n42), .B2(
        \pc_target[30][9] ), .ZN(n62) );
  INV_X1 U112 ( .A(n63), .ZN(n5543) );
  AOI22_X1 U113 ( .A1(Set_target[11]), .A2(n3798), .B1(n42), .B2(
        \pc_target[30][11] ), .ZN(n63) );
  INV_X1 U114 ( .A(n64), .ZN(n5544) );
  AOI22_X1 U115 ( .A1(Set_target[13]), .A2(n3798), .B1(n42), .B2(
        \pc_target[30][13] ), .ZN(n64) );
  INV_X1 U116 ( .A(n65), .ZN(n5545) );
  AOI22_X1 U117 ( .A1(Set_target[15]), .A2(n3798), .B1(n42), .B2(
        \pc_target[30][15] ), .ZN(n65) );
  INV_X1 U118 ( .A(n66), .ZN(n5546) );
  AOI22_X1 U119 ( .A1(Set_target[17]), .A2(n3798), .B1(n42), .B2(
        \pc_target[30][17] ), .ZN(n66) );
  INV_X1 U120 ( .A(n67), .ZN(n5547) );
  AOI22_X1 U121 ( .A1(Set_target[19]), .A2(n3798), .B1(n42), .B2(
        \pc_target[30][19] ), .ZN(n67) );
  INV_X1 U122 ( .A(n68), .ZN(n5548) );
  AOI22_X1 U123 ( .A1(Set_target[21]), .A2(n3798), .B1(n42), .B2(
        \pc_target[30][21] ), .ZN(n68) );
  INV_X1 U124 ( .A(n69), .ZN(n5549) );
  AOI22_X1 U125 ( .A1(Set_target[23]), .A2(n3798), .B1(n42), .B2(
        \pc_target[30][23] ), .ZN(n69) );
  INV_X1 U126 ( .A(n70), .ZN(n5550) );
  AOI22_X1 U127 ( .A1(Set_target[25]), .A2(n3798), .B1(n42), .B2(
        \pc_target[30][25] ), .ZN(n70) );
  INV_X1 U128 ( .A(n71), .ZN(n5551) );
  AOI22_X1 U129 ( .A1(Set_target[27]), .A2(n3798), .B1(n42), .B2(
        \pc_target[30][27] ), .ZN(n71) );
  INV_X1 U130 ( .A(n72), .ZN(n5552) );
  AOI22_X1 U131 ( .A1(Set_target[29]), .A2(n3798), .B1(n42), .B2(
        \pc_target[30][29] ), .ZN(n72) );
  INV_X1 U132 ( .A(n73), .ZN(n5553) );
  AOI22_X1 U133 ( .A1(Set_target[31]), .A2(n3798), .B1(n42), .B2(
        \pc_target[30][31] ), .ZN(n73) );
  OAI22_X1 U136 ( .A1(n75), .A2(n76), .B1(n77), .B2(n78), .ZN(n5554) );
  OAI22_X1 U137 ( .A1(n79), .A2(n76), .B1(n77), .B2(n80), .ZN(n5555) );
  OAI22_X1 U138 ( .A1(n81), .A2(n76), .B1(n77), .B2(n82), .ZN(n5556) );
  OAI22_X1 U139 ( .A1(n83), .A2(n76), .B1(n77), .B2(n84), .ZN(n5557) );
  OAI22_X1 U140 ( .A1(n85), .A2(n76), .B1(n77), .B2(n86), .ZN(n5558) );
  OAI22_X1 U141 ( .A1(n87), .A2(n76), .B1(n77), .B2(n88), .ZN(n5559) );
  OAI22_X1 U142 ( .A1(n89), .A2(n76), .B1(n77), .B2(n90), .ZN(n5560) );
  OAI22_X1 U143 ( .A1(n91), .A2(n76), .B1(n77), .B2(n92), .ZN(n5561) );
  OAI22_X1 U144 ( .A1(n93), .A2(n76), .B1(n77), .B2(n94), .ZN(n5562) );
  OAI22_X1 U145 ( .A1(n95), .A2(n76), .B1(n77), .B2(n96), .ZN(n5563) );
  OAI22_X1 U146 ( .A1(n97), .A2(n76), .B1(n77), .B2(n98), .ZN(n5564) );
  OAI22_X1 U147 ( .A1(n99), .A2(n76), .B1(n77), .B2(n100), .ZN(n5565) );
  OAI22_X1 U148 ( .A1(n101), .A2(n76), .B1(n77), .B2(n102), .ZN(n5566) );
  OAI22_X1 U149 ( .A1(n103), .A2(n76), .B1(n77), .B2(n104), .ZN(n5567) );
  OAI22_X1 U150 ( .A1(n105), .A2(n76), .B1(n77), .B2(n106), .ZN(n5568) );
  OAI22_X1 U151 ( .A1(n107), .A2(n76), .B1(n77), .B2(n108), .ZN(n5569) );
  OAI22_X1 U152 ( .A1(n109), .A2(n76), .B1(n77), .B2(n110), .ZN(n5570) );
  OAI22_X1 U153 ( .A1(n111), .A2(n76), .B1(n77), .B2(n112), .ZN(n5571) );
  OAI22_X1 U154 ( .A1(n113), .A2(n76), .B1(n77), .B2(n114), .ZN(n5572) );
  OAI22_X1 U155 ( .A1(n115), .A2(n76), .B1(n77), .B2(n116), .ZN(n5573) );
  OAI22_X1 U156 ( .A1(n117), .A2(n76), .B1(n77), .B2(n118), .ZN(n5574) );
  OAI22_X1 U157 ( .A1(n119), .A2(n76), .B1(n77), .B2(n120), .ZN(n5575) );
  OAI22_X1 U158 ( .A1(n121), .A2(n76), .B1(n77), .B2(n122), .ZN(n5576) );
  OAI22_X1 U159 ( .A1(n123), .A2(n76), .B1(n77), .B2(n124), .ZN(n5577) );
  OAI22_X1 U160 ( .A1(n125), .A2(n76), .B1(n77), .B2(n126), .ZN(n5578) );
  OAI22_X1 U161 ( .A1(n127), .A2(n76), .B1(n77), .B2(n128), .ZN(n5579) );
  OAI22_X1 U162 ( .A1(n129), .A2(n76), .B1(n77), .B2(n130), .ZN(n5580) );
  OAI22_X1 U163 ( .A1(n131), .A2(n76), .B1(n77), .B2(n132), .ZN(n5581) );
  OAI22_X1 U164 ( .A1(n133), .A2(n76), .B1(n77), .B2(n134), .ZN(n5582) );
  OAI22_X1 U165 ( .A1(n135), .A2(n76), .B1(n77), .B2(n136), .ZN(n5583) );
  OAI22_X1 U166 ( .A1(n137), .A2(n76), .B1(n77), .B2(n138), .ZN(n5584) );
  OAI22_X1 U167 ( .A1(n139), .A2(n76), .B1(n77), .B2(n140), .ZN(n5585) );
  OAI22_X1 U170 ( .A1(n75), .A2(n142), .B1(n143), .B2(n144), .ZN(n5586) );
  OAI22_X1 U171 ( .A1(n79), .A2(n142), .B1(n143), .B2(n145), .ZN(n5587) );
  OAI22_X1 U172 ( .A1(n81), .A2(n142), .B1(n143), .B2(n146), .ZN(n5588) );
  OAI22_X1 U173 ( .A1(n83), .A2(n142), .B1(n143), .B2(n147), .ZN(n5589) );
  OAI22_X1 U174 ( .A1(n85), .A2(n142), .B1(n143), .B2(n148), .ZN(n5590) );
  OAI22_X1 U175 ( .A1(n87), .A2(n142), .B1(n143), .B2(n149), .ZN(n5591) );
  OAI22_X1 U176 ( .A1(n89), .A2(n142), .B1(n143), .B2(n150), .ZN(n5592) );
  OAI22_X1 U177 ( .A1(n91), .A2(n142), .B1(n143), .B2(n151), .ZN(n5593) );
  OAI22_X1 U178 ( .A1(n93), .A2(n142), .B1(n143), .B2(n152), .ZN(n5594) );
  OAI22_X1 U179 ( .A1(n95), .A2(n142), .B1(n143), .B2(n153), .ZN(n5595) );
  OAI22_X1 U180 ( .A1(n97), .A2(n142), .B1(n143), .B2(n154), .ZN(n5596) );
  OAI22_X1 U181 ( .A1(n99), .A2(n142), .B1(n143), .B2(n155), .ZN(n5597) );
  OAI22_X1 U182 ( .A1(n101), .A2(n142), .B1(n143), .B2(n156), .ZN(n5598) );
  OAI22_X1 U183 ( .A1(n103), .A2(n142), .B1(n143), .B2(n157), .ZN(n5599) );
  OAI22_X1 U184 ( .A1(n105), .A2(n142), .B1(n143), .B2(n158), .ZN(n5600) );
  OAI22_X1 U185 ( .A1(n107), .A2(n142), .B1(n143), .B2(n159), .ZN(n5601) );
  OAI22_X1 U186 ( .A1(n109), .A2(n142), .B1(n143), .B2(n160), .ZN(n5602) );
  OAI22_X1 U187 ( .A1(n111), .A2(n142), .B1(n143), .B2(n161), .ZN(n5603) );
  OAI22_X1 U188 ( .A1(n113), .A2(n142), .B1(n143), .B2(n162), .ZN(n5604) );
  OAI22_X1 U189 ( .A1(n115), .A2(n142), .B1(n143), .B2(n163), .ZN(n5605) );
  OAI22_X1 U190 ( .A1(n117), .A2(n142), .B1(n143), .B2(n164), .ZN(n5606) );
  OAI22_X1 U191 ( .A1(n119), .A2(n142), .B1(n143), .B2(n165), .ZN(n5607) );
  OAI22_X1 U192 ( .A1(n121), .A2(n142), .B1(n143), .B2(n166), .ZN(n5608) );
  OAI22_X1 U193 ( .A1(n123), .A2(n142), .B1(n143), .B2(n167), .ZN(n5609) );
  OAI22_X1 U194 ( .A1(n125), .A2(n142), .B1(n143), .B2(n168), .ZN(n5610) );
  OAI22_X1 U195 ( .A1(n127), .A2(n142), .B1(n143), .B2(n169), .ZN(n5611) );
  OAI22_X1 U196 ( .A1(n129), .A2(n142), .B1(n143), .B2(n170), .ZN(n5612) );
  OAI22_X1 U197 ( .A1(n131), .A2(n142), .B1(n143), .B2(n171), .ZN(n5613) );
  OAI22_X1 U198 ( .A1(n133), .A2(n142), .B1(n143), .B2(n172), .ZN(n5614) );
  OAI22_X1 U199 ( .A1(n135), .A2(n142), .B1(n143), .B2(n173), .ZN(n5615) );
  OAI22_X1 U200 ( .A1(n137), .A2(n142), .B1(n143), .B2(n174), .ZN(n5616) );
  OAI22_X1 U201 ( .A1(n139), .A2(n142), .B1(n143), .B2(n175), .ZN(n5617) );
  INV_X1 U205 ( .A(n179), .ZN(n5618) );
  AOI22_X1 U206 ( .A1(Set_target[30]), .A2(n3797), .B1(n181), .B2(
        \pc_target[27][30] ), .ZN(n179) );
  INV_X1 U207 ( .A(n182), .ZN(n5619) );
  AOI22_X1 U208 ( .A1(Set_target[28]), .A2(n3797), .B1(n181), .B2(
        \pc_target[27][28] ), .ZN(n182) );
  INV_X1 U209 ( .A(n183), .ZN(n5620) );
  AOI22_X1 U210 ( .A1(Set_target[26]), .A2(n3797), .B1(n181), .B2(
        \pc_target[27][26] ), .ZN(n183) );
  INV_X1 U211 ( .A(n184), .ZN(n5621) );
  AOI22_X1 U212 ( .A1(Set_target[24]), .A2(n3797), .B1(n181), .B2(
        \pc_target[27][24] ), .ZN(n184) );
  INV_X1 U213 ( .A(n185), .ZN(n5622) );
  AOI22_X1 U214 ( .A1(Set_target[22]), .A2(n3797), .B1(n181), .B2(
        \pc_target[27][22] ), .ZN(n185) );
  INV_X1 U215 ( .A(n186), .ZN(n5623) );
  AOI22_X1 U216 ( .A1(Set_target[20]), .A2(n3797), .B1(n181), .B2(
        \pc_target[27][20] ), .ZN(n186) );
  INV_X1 U217 ( .A(n187), .ZN(n5624) );
  AOI22_X1 U218 ( .A1(Set_target[18]), .A2(n3797), .B1(n181), .B2(
        \pc_target[27][18] ), .ZN(n187) );
  INV_X1 U219 ( .A(n188), .ZN(n5625) );
  AOI22_X1 U220 ( .A1(Set_target[16]), .A2(n3797), .B1(n181), .B2(
        \pc_target[27][16] ), .ZN(n188) );
  INV_X1 U221 ( .A(n189), .ZN(n5626) );
  AOI22_X1 U222 ( .A1(Set_target[14]), .A2(n3797), .B1(n181), .B2(
        \pc_target[27][14] ), .ZN(n189) );
  INV_X1 U223 ( .A(n190), .ZN(n5627) );
  AOI22_X1 U224 ( .A1(Set_target[12]), .A2(n3797), .B1(n181), .B2(
        \pc_target[27][12] ), .ZN(n190) );
  INV_X1 U225 ( .A(n191), .ZN(n5628) );
  AOI22_X1 U226 ( .A1(Set_target[10]), .A2(n3797), .B1(n181), .B2(
        \pc_target[27][10] ), .ZN(n191) );
  INV_X1 U227 ( .A(n192), .ZN(n5629) );
  AOI22_X1 U228 ( .A1(Set_target[8]), .A2(n3797), .B1(n181), .B2(
        \pc_target[27][8] ), .ZN(n192) );
  INV_X1 U229 ( .A(n193), .ZN(n5630) );
  AOI22_X1 U230 ( .A1(Set_target[6]), .A2(n3797), .B1(n181), .B2(
        \pc_target[27][6] ), .ZN(n193) );
  INV_X1 U231 ( .A(n194), .ZN(n5631) );
  AOI22_X1 U232 ( .A1(Set_target[4]), .A2(n3797), .B1(n181), .B2(
        \pc_target[27][4] ), .ZN(n194) );
  INV_X1 U233 ( .A(n195), .ZN(n5632) );
  AOI22_X1 U234 ( .A1(Set_target[2]), .A2(n3797), .B1(n181), .B2(
        \pc_target[27][2] ), .ZN(n195) );
  INV_X1 U235 ( .A(n196), .ZN(n5633) );
  AOI22_X1 U236 ( .A1(Set_target[0]), .A2(n3797), .B1(n181), .B2(
        \pc_target[27][0] ), .ZN(n196) );
  INV_X1 U237 ( .A(n197), .ZN(n5634) );
  AOI22_X1 U238 ( .A1(Set_target[1]), .A2(n3797), .B1(n181), .B2(
        \pc_target[27][1] ), .ZN(n197) );
  INV_X1 U239 ( .A(n198), .ZN(n5635) );
  AOI22_X1 U240 ( .A1(Set_target[3]), .A2(n3797), .B1(n181), .B2(
        \pc_target[27][3] ), .ZN(n198) );
  INV_X1 U241 ( .A(n199), .ZN(n5636) );
  AOI22_X1 U242 ( .A1(Set_target[5]), .A2(n3797), .B1(n181), .B2(
        \pc_target[27][5] ), .ZN(n199) );
  INV_X1 U243 ( .A(n200), .ZN(n5637) );
  AOI22_X1 U244 ( .A1(Set_target[7]), .A2(n3797), .B1(n181), .B2(
        \pc_target[27][7] ), .ZN(n200) );
  INV_X1 U245 ( .A(n201), .ZN(n5638) );
  AOI22_X1 U246 ( .A1(Set_target[9]), .A2(n3797), .B1(n181), .B2(
        \pc_target[27][9] ), .ZN(n201) );
  INV_X1 U247 ( .A(n202), .ZN(n5639) );
  AOI22_X1 U248 ( .A1(Set_target[11]), .A2(n3797), .B1(n181), .B2(
        \pc_target[27][11] ), .ZN(n202) );
  INV_X1 U249 ( .A(n203), .ZN(n5640) );
  AOI22_X1 U250 ( .A1(Set_target[13]), .A2(n3797), .B1(n181), .B2(
        \pc_target[27][13] ), .ZN(n203) );
  INV_X1 U251 ( .A(n204), .ZN(n5641) );
  AOI22_X1 U252 ( .A1(Set_target[15]), .A2(n3797), .B1(n181), .B2(
        \pc_target[27][15] ), .ZN(n204) );
  INV_X1 U253 ( .A(n205), .ZN(n5642) );
  AOI22_X1 U254 ( .A1(Set_target[17]), .A2(n3797), .B1(n181), .B2(
        \pc_target[27][17] ), .ZN(n205) );
  INV_X1 U255 ( .A(n206), .ZN(n5643) );
  AOI22_X1 U256 ( .A1(Set_target[19]), .A2(n3797), .B1(n181), .B2(
        \pc_target[27][19] ), .ZN(n206) );
  INV_X1 U257 ( .A(n207), .ZN(n5644) );
  AOI22_X1 U258 ( .A1(Set_target[21]), .A2(n3797), .B1(n181), .B2(
        \pc_target[27][21] ), .ZN(n207) );
  INV_X1 U259 ( .A(n208), .ZN(n5645) );
  AOI22_X1 U260 ( .A1(Set_target[23]), .A2(n3797), .B1(n181), .B2(
        \pc_target[27][23] ), .ZN(n208) );
  INV_X1 U261 ( .A(n209), .ZN(n5646) );
  AOI22_X1 U262 ( .A1(Set_target[25]), .A2(n3797), .B1(n181), .B2(
        \pc_target[27][25] ), .ZN(n209) );
  INV_X1 U263 ( .A(n210), .ZN(n5647) );
  AOI22_X1 U264 ( .A1(Set_target[27]), .A2(n3797), .B1(n181), .B2(
        \pc_target[27][27] ), .ZN(n210) );
  INV_X1 U265 ( .A(n211), .ZN(n5648) );
  AOI22_X1 U266 ( .A1(Set_target[29]), .A2(n3797), .B1(n181), .B2(
        \pc_target[27][29] ), .ZN(n211) );
  INV_X1 U267 ( .A(n212), .ZN(n5649) );
  AOI22_X1 U268 ( .A1(Set_target[31]), .A2(n3797), .B1(n181), .B2(
        \pc_target[27][31] ), .ZN(n212) );
  INV_X1 U271 ( .A(n214), .ZN(n5650) );
  AOI22_X1 U272 ( .A1(Set_target[30]), .A2(n215), .B1(n216), .B2(
        \pc_target[26][30] ), .ZN(n214) );
  INV_X1 U273 ( .A(n217), .ZN(n5651) );
  AOI22_X1 U274 ( .A1(Set_target[28]), .A2(n215), .B1(n216), .B2(
        \pc_target[26][28] ), .ZN(n217) );
  INV_X1 U275 ( .A(n218), .ZN(n5652) );
  AOI22_X1 U276 ( .A1(Set_target[26]), .A2(n215), .B1(n216), .B2(
        \pc_target[26][26] ), .ZN(n218) );
  INV_X1 U277 ( .A(n219), .ZN(n5653) );
  AOI22_X1 U278 ( .A1(Set_target[24]), .A2(n215), .B1(n216), .B2(
        \pc_target[26][24] ), .ZN(n219) );
  INV_X1 U279 ( .A(n220), .ZN(n5654) );
  AOI22_X1 U280 ( .A1(Set_target[22]), .A2(n215), .B1(n216), .B2(
        \pc_target[26][22] ), .ZN(n220) );
  INV_X1 U281 ( .A(n221), .ZN(n5655) );
  AOI22_X1 U282 ( .A1(Set_target[20]), .A2(n215), .B1(n216), .B2(
        \pc_target[26][20] ), .ZN(n221) );
  INV_X1 U283 ( .A(n222), .ZN(n5656) );
  AOI22_X1 U284 ( .A1(Set_target[18]), .A2(n215), .B1(n216), .B2(
        \pc_target[26][18] ), .ZN(n222) );
  INV_X1 U285 ( .A(n223), .ZN(n5657) );
  AOI22_X1 U286 ( .A1(Set_target[16]), .A2(n215), .B1(n216), .B2(
        \pc_target[26][16] ), .ZN(n223) );
  INV_X1 U287 ( .A(n224), .ZN(n5658) );
  AOI22_X1 U288 ( .A1(Set_target[14]), .A2(n215), .B1(n216), .B2(
        \pc_target[26][14] ), .ZN(n224) );
  INV_X1 U289 ( .A(n225), .ZN(n5659) );
  AOI22_X1 U290 ( .A1(Set_target[12]), .A2(n215), .B1(n216), .B2(
        \pc_target[26][12] ), .ZN(n225) );
  INV_X1 U291 ( .A(n226), .ZN(n5660) );
  AOI22_X1 U292 ( .A1(Set_target[10]), .A2(n215), .B1(n216), .B2(
        \pc_target[26][10] ), .ZN(n226) );
  INV_X1 U293 ( .A(n227), .ZN(n5661) );
  AOI22_X1 U294 ( .A1(Set_target[8]), .A2(n215), .B1(n216), .B2(
        \pc_target[26][8] ), .ZN(n227) );
  INV_X1 U295 ( .A(n228), .ZN(n5662) );
  AOI22_X1 U296 ( .A1(Set_target[6]), .A2(n215), .B1(n216), .B2(
        \pc_target[26][6] ), .ZN(n228) );
  INV_X1 U297 ( .A(n229), .ZN(n5663) );
  AOI22_X1 U298 ( .A1(Set_target[4]), .A2(n215), .B1(n216), .B2(
        \pc_target[26][4] ), .ZN(n229) );
  INV_X1 U299 ( .A(n230), .ZN(n5664) );
  AOI22_X1 U300 ( .A1(Set_target[2]), .A2(n215), .B1(n216), .B2(
        \pc_target[26][2] ), .ZN(n230) );
  INV_X1 U301 ( .A(n231), .ZN(n5665) );
  AOI22_X1 U302 ( .A1(Set_target[0]), .A2(n215), .B1(n216), .B2(
        \pc_target[26][0] ), .ZN(n231) );
  INV_X1 U303 ( .A(n232), .ZN(n5666) );
  AOI22_X1 U304 ( .A1(Set_target[1]), .A2(n215), .B1(n216), .B2(
        \pc_target[26][1] ), .ZN(n232) );
  INV_X1 U305 ( .A(n233), .ZN(n5667) );
  AOI22_X1 U306 ( .A1(Set_target[3]), .A2(n215), .B1(n216), .B2(
        \pc_target[26][3] ), .ZN(n233) );
  INV_X1 U307 ( .A(n234), .ZN(n5668) );
  AOI22_X1 U308 ( .A1(Set_target[5]), .A2(n215), .B1(n216), .B2(
        \pc_target[26][5] ), .ZN(n234) );
  INV_X1 U309 ( .A(n235), .ZN(n5669) );
  AOI22_X1 U310 ( .A1(Set_target[7]), .A2(n215), .B1(n216), .B2(
        \pc_target[26][7] ), .ZN(n235) );
  INV_X1 U311 ( .A(n236), .ZN(n5670) );
  AOI22_X1 U312 ( .A1(Set_target[9]), .A2(n215), .B1(n216), .B2(
        \pc_target[26][9] ), .ZN(n236) );
  INV_X1 U313 ( .A(n237), .ZN(n5671) );
  AOI22_X1 U314 ( .A1(Set_target[11]), .A2(n215), .B1(n216), .B2(
        \pc_target[26][11] ), .ZN(n237) );
  INV_X1 U315 ( .A(n238), .ZN(n5672) );
  AOI22_X1 U316 ( .A1(Set_target[13]), .A2(n215), .B1(n216), .B2(
        \pc_target[26][13] ), .ZN(n238) );
  INV_X1 U317 ( .A(n239), .ZN(n5673) );
  AOI22_X1 U318 ( .A1(Set_target[15]), .A2(n215), .B1(n216), .B2(
        \pc_target[26][15] ), .ZN(n239) );
  INV_X1 U319 ( .A(n240), .ZN(n5674) );
  AOI22_X1 U320 ( .A1(Set_target[17]), .A2(n215), .B1(n216), .B2(
        \pc_target[26][17] ), .ZN(n240) );
  INV_X1 U321 ( .A(n241), .ZN(n5675) );
  AOI22_X1 U322 ( .A1(Set_target[19]), .A2(n215), .B1(n216), .B2(
        \pc_target[26][19] ), .ZN(n241) );
  INV_X1 U323 ( .A(n242), .ZN(n5676) );
  AOI22_X1 U324 ( .A1(Set_target[21]), .A2(n215), .B1(n216), .B2(
        \pc_target[26][21] ), .ZN(n242) );
  INV_X1 U325 ( .A(n243), .ZN(n5677) );
  AOI22_X1 U326 ( .A1(Set_target[23]), .A2(n215), .B1(n216), .B2(
        \pc_target[26][23] ), .ZN(n243) );
  INV_X1 U327 ( .A(n244), .ZN(n5678) );
  AOI22_X1 U328 ( .A1(Set_target[25]), .A2(n215), .B1(n216), .B2(
        \pc_target[26][25] ), .ZN(n244) );
  INV_X1 U329 ( .A(n245), .ZN(n5679) );
  AOI22_X1 U330 ( .A1(Set_target[27]), .A2(n215), .B1(n216), .B2(
        \pc_target[26][27] ), .ZN(n245) );
  INV_X1 U331 ( .A(n246), .ZN(n5680) );
  AOI22_X1 U332 ( .A1(Set_target[29]), .A2(n215), .B1(n216), .B2(
        \pc_target[26][29] ), .ZN(n246) );
  INV_X1 U333 ( .A(n247), .ZN(n5681) );
  AOI22_X1 U334 ( .A1(Set_target[31]), .A2(n215), .B1(n216), .B2(
        \pc_target[26][31] ), .ZN(n247) );
  OAI22_X1 U337 ( .A1(n75), .A2(n248), .B1(n249), .B2(n250), .ZN(n5682) );
  OAI22_X1 U338 ( .A1(n79), .A2(n248), .B1(n249), .B2(n251), .ZN(n5683) );
  OAI22_X1 U339 ( .A1(n81), .A2(n248), .B1(n249), .B2(n252), .ZN(n5684) );
  OAI22_X1 U340 ( .A1(n83), .A2(n248), .B1(n249), .B2(n253), .ZN(n5685) );
  OAI22_X1 U341 ( .A1(n85), .A2(n248), .B1(n249), .B2(n254), .ZN(n5686) );
  OAI22_X1 U342 ( .A1(n87), .A2(n248), .B1(n249), .B2(n255), .ZN(n5687) );
  OAI22_X1 U343 ( .A1(n89), .A2(n248), .B1(n249), .B2(n256), .ZN(n5688) );
  OAI22_X1 U344 ( .A1(n91), .A2(n248), .B1(n249), .B2(n257), .ZN(n5689) );
  OAI22_X1 U345 ( .A1(n93), .A2(n248), .B1(n249), .B2(n258), .ZN(n5690) );
  OAI22_X1 U346 ( .A1(n95), .A2(n248), .B1(n249), .B2(n259), .ZN(n5691) );
  OAI22_X1 U347 ( .A1(n97), .A2(n248), .B1(n249), .B2(n260), .ZN(n5692) );
  OAI22_X1 U348 ( .A1(n99), .A2(n248), .B1(n249), .B2(n261), .ZN(n5693) );
  OAI22_X1 U349 ( .A1(n101), .A2(n248), .B1(n249), .B2(n262), .ZN(n5694) );
  OAI22_X1 U350 ( .A1(n103), .A2(n248), .B1(n249), .B2(n263), .ZN(n5695) );
  OAI22_X1 U351 ( .A1(n105), .A2(n248), .B1(n249), .B2(n264), .ZN(n5696) );
  OAI22_X1 U352 ( .A1(n107), .A2(n248), .B1(n249), .B2(n265), .ZN(n5697) );
  OAI22_X1 U353 ( .A1(n109), .A2(n248), .B1(n249), .B2(n266), .ZN(n5698) );
  OAI22_X1 U354 ( .A1(n111), .A2(n248), .B1(n249), .B2(n267), .ZN(n5699) );
  OAI22_X1 U355 ( .A1(n113), .A2(n248), .B1(n249), .B2(n268), .ZN(n5700) );
  OAI22_X1 U356 ( .A1(n115), .A2(n248), .B1(n249), .B2(n269), .ZN(n5701) );
  OAI22_X1 U357 ( .A1(n117), .A2(n248), .B1(n249), .B2(n270), .ZN(n5702) );
  OAI22_X1 U358 ( .A1(n119), .A2(n248), .B1(n249), .B2(n271), .ZN(n5703) );
  OAI22_X1 U359 ( .A1(n121), .A2(n248), .B1(n249), .B2(n272), .ZN(n5704) );
  OAI22_X1 U360 ( .A1(n123), .A2(n248), .B1(n249), .B2(n273), .ZN(n5705) );
  OAI22_X1 U361 ( .A1(n125), .A2(n248), .B1(n249), .B2(n274), .ZN(n5706) );
  OAI22_X1 U362 ( .A1(n127), .A2(n248), .B1(n249), .B2(n275), .ZN(n5707) );
  OAI22_X1 U363 ( .A1(n129), .A2(n248), .B1(n249), .B2(n276), .ZN(n5708) );
  OAI22_X1 U364 ( .A1(n131), .A2(n248), .B1(n249), .B2(n277), .ZN(n5709) );
  OAI22_X1 U365 ( .A1(n133), .A2(n248), .B1(n249), .B2(n278), .ZN(n5710) );
  OAI22_X1 U366 ( .A1(n135), .A2(n248), .B1(n249), .B2(n279), .ZN(n5711) );
  OAI22_X1 U367 ( .A1(n137), .A2(n248), .B1(n249), .B2(n280), .ZN(n5712) );
  OAI22_X1 U368 ( .A1(n139), .A2(n248), .B1(n249), .B2(n281), .ZN(n5713) );
  OAI22_X1 U371 ( .A1(n75), .A2(n282), .B1(n3444), .B2(n284), .ZN(n5714) );
  OAI22_X1 U372 ( .A1(n79), .A2(n282), .B1(n3444), .B2(n285), .ZN(n5715) );
  OAI22_X1 U373 ( .A1(n81), .A2(n282), .B1(n3444), .B2(n286), .ZN(n5716) );
  OAI22_X1 U374 ( .A1(n83), .A2(n282), .B1(n3444), .B2(n287), .ZN(n5717) );
  OAI22_X1 U375 ( .A1(n85), .A2(n282), .B1(n3444), .B2(n288), .ZN(n5718) );
  OAI22_X1 U376 ( .A1(n87), .A2(n282), .B1(n3444), .B2(n289), .ZN(n5719) );
  OAI22_X1 U377 ( .A1(n89), .A2(n282), .B1(n3444), .B2(n290), .ZN(n5720) );
  OAI22_X1 U378 ( .A1(n91), .A2(n282), .B1(n3444), .B2(n291), .ZN(n5721) );
  OAI22_X1 U379 ( .A1(n93), .A2(n282), .B1(n3444), .B2(n292), .ZN(n5722) );
  OAI22_X1 U380 ( .A1(n95), .A2(n282), .B1(n3444), .B2(n293), .ZN(n5723) );
  OAI22_X1 U381 ( .A1(n97), .A2(n282), .B1(n3444), .B2(n294), .ZN(n5724) );
  OAI22_X1 U382 ( .A1(n99), .A2(n282), .B1(n3444), .B2(n295), .ZN(n5725) );
  OAI22_X1 U383 ( .A1(n101), .A2(n282), .B1(n3444), .B2(n296), .ZN(n5726) );
  OAI22_X1 U384 ( .A1(n103), .A2(n282), .B1(n3444), .B2(n297), .ZN(n5727) );
  OAI22_X1 U385 ( .A1(n105), .A2(n282), .B1(n3444), .B2(n298), .ZN(n5728) );
  OAI22_X1 U386 ( .A1(n107), .A2(n282), .B1(n3444), .B2(n299), .ZN(n5729) );
  OAI22_X1 U387 ( .A1(n109), .A2(n282), .B1(n3444), .B2(n300), .ZN(n5730) );
  OAI22_X1 U388 ( .A1(n111), .A2(n282), .B1(n3444), .B2(n301), .ZN(n5731) );
  OAI22_X1 U389 ( .A1(n113), .A2(n282), .B1(n3444), .B2(n302), .ZN(n5732) );
  OAI22_X1 U390 ( .A1(n115), .A2(n282), .B1(n3444), .B2(n303), .ZN(n5733) );
  OAI22_X1 U391 ( .A1(n117), .A2(n282), .B1(n3444), .B2(n304), .ZN(n5734) );
  OAI22_X1 U392 ( .A1(n119), .A2(n282), .B1(n3444), .B2(n305), .ZN(n5735) );
  OAI22_X1 U393 ( .A1(n121), .A2(n282), .B1(n3444), .B2(n306), .ZN(n5736) );
  OAI22_X1 U394 ( .A1(n123), .A2(n282), .B1(n3444), .B2(n307), .ZN(n5737) );
  OAI22_X1 U395 ( .A1(n125), .A2(n282), .B1(n3444), .B2(n308), .ZN(n5738) );
  OAI22_X1 U396 ( .A1(n127), .A2(n282), .B1(n3444), .B2(n309), .ZN(n5739) );
  OAI22_X1 U397 ( .A1(n129), .A2(n282), .B1(n3444), .B2(n310), .ZN(n5740) );
  OAI22_X1 U398 ( .A1(n131), .A2(n282), .B1(n3444), .B2(n311), .ZN(n5741) );
  OAI22_X1 U399 ( .A1(n133), .A2(n282), .B1(n3444), .B2(n312), .ZN(n5742) );
  OAI22_X1 U400 ( .A1(n135), .A2(n282), .B1(n3444), .B2(n313), .ZN(n5743) );
  OAI22_X1 U401 ( .A1(n137), .A2(n282), .B1(n3444), .B2(n314), .ZN(n5744) );
  OAI22_X1 U402 ( .A1(n139), .A2(n282), .B1(n3444), .B2(n315), .ZN(n5745) );
  OAI22_X1 U406 ( .A1(n75), .A2(n317), .B1(n318), .B2(n319), .ZN(n5746) );
  OAI22_X1 U407 ( .A1(n79), .A2(n317), .B1(n318), .B2(n320), .ZN(n5747) );
  OAI22_X1 U408 ( .A1(n81), .A2(n317), .B1(n318), .B2(n321), .ZN(n5748) );
  OAI22_X1 U409 ( .A1(n83), .A2(n317), .B1(n318), .B2(n322), .ZN(n5749) );
  OAI22_X1 U410 ( .A1(n85), .A2(n317), .B1(n318), .B2(n323), .ZN(n5750) );
  OAI22_X1 U411 ( .A1(n87), .A2(n317), .B1(n318), .B2(n324), .ZN(n5751) );
  OAI22_X1 U412 ( .A1(n89), .A2(n317), .B1(n318), .B2(n325), .ZN(n5752) );
  OAI22_X1 U413 ( .A1(n91), .A2(n317), .B1(n318), .B2(n326), .ZN(n5753) );
  OAI22_X1 U414 ( .A1(n93), .A2(n317), .B1(n318), .B2(n327), .ZN(n5754) );
  OAI22_X1 U415 ( .A1(n95), .A2(n317), .B1(n318), .B2(n328), .ZN(n5755) );
  OAI22_X1 U416 ( .A1(n97), .A2(n317), .B1(n318), .B2(n329), .ZN(n5756) );
  OAI22_X1 U417 ( .A1(n99), .A2(n317), .B1(n318), .B2(n330), .ZN(n5757) );
  OAI22_X1 U418 ( .A1(n101), .A2(n317), .B1(n318), .B2(n331), .ZN(n5758) );
  OAI22_X1 U419 ( .A1(n103), .A2(n317), .B1(n318), .B2(n332), .ZN(n5759) );
  OAI22_X1 U420 ( .A1(n105), .A2(n317), .B1(n318), .B2(n333), .ZN(n5760) );
  OAI22_X1 U421 ( .A1(n107), .A2(n317), .B1(n318), .B2(n334), .ZN(n5761) );
  OAI22_X1 U422 ( .A1(n109), .A2(n317), .B1(n318), .B2(n335), .ZN(n5762) );
  OAI22_X1 U423 ( .A1(n111), .A2(n317), .B1(n318), .B2(n336), .ZN(n5763) );
  OAI22_X1 U424 ( .A1(n113), .A2(n317), .B1(n318), .B2(n337), .ZN(n5764) );
  OAI22_X1 U425 ( .A1(n115), .A2(n317), .B1(n318), .B2(n338), .ZN(n5765) );
  OAI22_X1 U426 ( .A1(n117), .A2(n317), .B1(n318), .B2(n339), .ZN(n5766) );
  OAI22_X1 U427 ( .A1(n119), .A2(n317), .B1(n318), .B2(n340), .ZN(n5767) );
  OAI22_X1 U428 ( .A1(n121), .A2(n317), .B1(n318), .B2(n341), .ZN(n5768) );
  OAI22_X1 U429 ( .A1(n123), .A2(n317), .B1(n318), .B2(n342), .ZN(n5769) );
  OAI22_X1 U430 ( .A1(n125), .A2(n317), .B1(n318), .B2(n343), .ZN(n5770) );
  OAI22_X1 U431 ( .A1(n127), .A2(n317), .B1(n318), .B2(n344), .ZN(n5771) );
  OAI22_X1 U432 ( .A1(n129), .A2(n317), .B1(n318), .B2(n345), .ZN(n5772) );
  OAI22_X1 U433 ( .A1(n131), .A2(n317), .B1(n318), .B2(n346), .ZN(n5773) );
  OAI22_X1 U434 ( .A1(n133), .A2(n317), .B1(n318), .B2(n347), .ZN(n5774) );
  OAI22_X1 U435 ( .A1(n135), .A2(n317), .B1(n318), .B2(n348), .ZN(n5775) );
  OAI22_X1 U436 ( .A1(n137), .A2(n317), .B1(n318), .B2(n349), .ZN(n5776) );
  OAI22_X1 U437 ( .A1(n139), .A2(n317), .B1(n318), .B2(n350), .ZN(n5777) );
  OAI22_X1 U440 ( .A1(n75), .A2(n352), .B1(n353), .B2(n354), .ZN(n5778) );
  OAI22_X1 U441 ( .A1(n79), .A2(n352), .B1(n353), .B2(n355), .ZN(n5779) );
  OAI22_X1 U442 ( .A1(n81), .A2(n352), .B1(n353), .B2(n356), .ZN(n5780) );
  OAI22_X1 U443 ( .A1(n83), .A2(n352), .B1(n353), .B2(n357), .ZN(n5781) );
  OAI22_X1 U444 ( .A1(n85), .A2(n352), .B1(n353), .B2(n358), .ZN(n5782) );
  OAI22_X1 U445 ( .A1(n87), .A2(n352), .B1(n353), .B2(n359), .ZN(n5783) );
  OAI22_X1 U446 ( .A1(n89), .A2(n352), .B1(n353), .B2(n360), .ZN(n5784) );
  OAI22_X1 U447 ( .A1(n91), .A2(n352), .B1(n353), .B2(n361), .ZN(n5785) );
  OAI22_X1 U448 ( .A1(n93), .A2(n352), .B1(n353), .B2(n362), .ZN(n5786) );
  OAI22_X1 U449 ( .A1(n95), .A2(n352), .B1(n353), .B2(n363), .ZN(n5787) );
  OAI22_X1 U450 ( .A1(n97), .A2(n352), .B1(n353), .B2(n364), .ZN(n5788) );
  OAI22_X1 U451 ( .A1(n99), .A2(n352), .B1(n353), .B2(n365), .ZN(n5789) );
  OAI22_X1 U452 ( .A1(n101), .A2(n352), .B1(n353), .B2(n366), .ZN(n5790) );
  OAI22_X1 U453 ( .A1(n103), .A2(n352), .B1(n353), .B2(n367), .ZN(n5791) );
  OAI22_X1 U454 ( .A1(n105), .A2(n352), .B1(n353), .B2(n368), .ZN(n5792) );
  OAI22_X1 U455 ( .A1(n107), .A2(n352), .B1(n353), .B2(n369), .ZN(n5793) );
  OAI22_X1 U456 ( .A1(n109), .A2(n352), .B1(n353), .B2(n370), .ZN(n5794) );
  OAI22_X1 U457 ( .A1(n111), .A2(n352), .B1(n353), .B2(n371), .ZN(n5795) );
  OAI22_X1 U458 ( .A1(n113), .A2(n352), .B1(n353), .B2(n372), .ZN(n5796) );
  OAI22_X1 U459 ( .A1(n115), .A2(n352), .B1(n353), .B2(n373), .ZN(n5797) );
  OAI22_X1 U460 ( .A1(n117), .A2(n352), .B1(n353), .B2(n374), .ZN(n5798) );
  OAI22_X1 U461 ( .A1(n119), .A2(n352), .B1(n353), .B2(n375), .ZN(n5799) );
  OAI22_X1 U462 ( .A1(n121), .A2(n352), .B1(n353), .B2(n376), .ZN(n5800) );
  OAI22_X1 U463 ( .A1(n123), .A2(n352), .B1(n353), .B2(n377), .ZN(n5801) );
  OAI22_X1 U464 ( .A1(n125), .A2(n352), .B1(n353), .B2(n378), .ZN(n5802) );
  OAI22_X1 U465 ( .A1(n127), .A2(n352), .B1(n353), .B2(n379), .ZN(n5803) );
  OAI22_X1 U466 ( .A1(n129), .A2(n352), .B1(n353), .B2(n380), .ZN(n5804) );
  OAI22_X1 U467 ( .A1(n131), .A2(n352), .B1(n353), .B2(n381), .ZN(n5805) );
  OAI22_X1 U468 ( .A1(n133), .A2(n352), .B1(n353), .B2(n382), .ZN(n5806) );
  OAI22_X1 U469 ( .A1(n135), .A2(n352), .B1(n353), .B2(n383), .ZN(n5807) );
  OAI22_X1 U470 ( .A1(n137), .A2(n352), .B1(n353), .B2(n384), .ZN(n5808) );
  OAI22_X1 U471 ( .A1(n139), .A2(n352), .B1(n353), .B2(n385), .ZN(n5809) );
  INV_X1 U474 ( .A(n386), .ZN(n5810) );
  AOI22_X1 U475 ( .A1(Set_target[30]), .A2(n3799), .B1(n388), .B2(
        \pc_target[21][30] ), .ZN(n386) );
  INV_X1 U476 ( .A(n389), .ZN(n5811) );
  AOI22_X1 U477 ( .A1(Set_target[28]), .A2(n3799), .B1(n388), .B2(
        \pc_target[21][28] ), .ZN(n389) );
  INV_X1 U478 ( .A(n390), .ZN(n5812) );
  AOI22_X1 U479 ( .A1(Set_target[26]), .A2(n3799), .B1(n388), .B2(
        \pc_target[21][26] ), .ZN(n390) );
  INV_X1 U480 ( .A(n391), .ZN(n5813) );
  AOI22_X1 U481 ( .A1(Set_target[24]), .A2(n3799), .B1(n388), .B2(
        \pc_target[21][24] ), .ZN(n391) );
  INV_X1 U482 ( .A(n392), .ZN(n5814) );
  AOI22_X1 U483 ( .A1(Set_target[22]), .A2(n3799), .B1(n388), .B2(
        \pc_target[21][22] ), .ZN(n392) );
  INV_X1 U484 ( .A(n393), .ZN(n5815) );
  AOI22_X1 U485 ( .A1(Set_target[20]), .A2(n3799), .B1(n388), .B2(
        \pc_target[21][20] ), .ZN(n393) );
  INV_X1 U486 ( .A(n394), .ZN(n5816) );
  AOI22_X1 U487 ( .A1(Set_target[18]), .A2(n3799), .B1(n388), .B2(
        \pc_target[21][18] ), .ZN(n394) );
  INV_X1 U488 ( .A(n395), .ZN(n5817) );
  AOI22_X1 U489 ( .A1(Set_target[16]), .A2(n3799), .B1(n388), .B2(
        \pc_target[21][16] ), .ZN(n395) );
  INV_X1 U490 ( .A(n396), .ZN(n5818) );
  AOI22_X1 U491 ( .A1(Set_target[14]), .A2(n3799), .B1(n388), .B2(
        \pc_target[21][14] ), .ZN(n396) );
  INV_X1 U492 ( .A(n397), .ZN(n5819) );
  AOI22_X1 U493 ( .A1(Set_target[12]), .A2(n3799), .B1(n388), .B2(
        \pc_target[21][12] ), .ZN(n397) );
  INV_X1 U494 ( .A(n398), .ZN(n5820) );
  AOI22_X1 U495 ( .A1(Set_target[10]), .A2(n3799), .B1(n388), .B2(
        \pc_target[21][10] ), .ZN(n398) );
  INV_X1 U496 ( .A(n399), .ZN(n5821) );
  AOI22_X1 U497 ( .A1(Set_target[8]), .A2(n3799), .B1(n388), .B2(
        \pc_target[21][8] ), .ZN(n399) );
  INV_X1 U498 ( .A(n400), .ZN(n5822) );
  AOI22_X1 U499 ( .A1(Set_target[6]), .A2(n3799), .B1(n388), .B2(
        \pc_target[21][6] ), .ZN(n400) );
  INV_X1 U500 ( .A(n401), .ZN(n5823) );
  AOI22_X1 U501 ( .A1(Set_target[4]), .A2(n3799), .B1(n388), .B2(
        \pc_target[21][4] ), .ZN(n401) );
  INV_X1 U502 ( .A(n402), .ZN(n5824) );
  AOI22_X1 U503 ( .A1(Set_target[2]), .A2(n3799), .B1(n388), .B2(
        \pc_target[21][2] ), .ZN(n402) );
  INV_X1 U504 ( .A(n403), .ZN(n5825) );
  AOI22_X1 U505 ( .A1(Set_target[0]), .A2(n3799), .B1(n388), .B2(
        \pc_target[21][0] ), .ZN(n403) );
  INV_X1 U506 ( .A(n404), .ZN(n5826) );
  AOI22_X1 U507 ( .A1(Set_target[1]), .A2(n3799), .B1(n388), .B2(
        \pc_target[21][1] ), .ZN(n404) );
  INV_X1 U508 ( .A(n405), .ZN(n5827) );
  AOI22_X1 U509 ( .A1(Set_target[3]), .A2(n3799), .B1(n388), .B2(
        \pc_target[21][3] ), .ZN(n405) );
  INV_X1 U510 ( .A(n406), .ZN(n5828) );
  AOI22_X1 U511 ( .A1(Set_target[5]), .A2(n3799), .B1(n388), .B2(
        \pc_target[21][5] ), .ZN(n406) );
  INV_X1 U512 ( .A(n407), .ZN(n5829) );
  AOI22_X1 U513 ( .A1(Set_target[7]), .A2(n3799), .B1(n388), .B2(
        \pc_target[21][7] ), .ZN(n407) );
  INV_X1 U514 ( .A(n408), .ZN(n5830) );
  AOI22_X1 U515 ( .A1(Set_target[9]), .A2(n3799), .B1(n388), .B2(
        \pc_target[21][9] ), .ZN(n408) );
  INV_X1 U516 ( .A(n409), .ZN(n5831) );
  AOI22_X1 U517 ( .A1(Set_target[11]), .A2(n3799), .B1(n388), .B2(
        \pc_target[21][11] ), .ZN(n409) );
  INV_X1 U518 ( .A(n410), .ZN(n5832) );
  AOI22_X1 U519 ( .A1(Set_target[13]), .A2(n3799), .B1(n388), .B2(
        \pc_target[21][13] ), .ZN(n410) );
  INV_X1 U520 ( .A(n411), .ZN(n5833) );
  AOI22_X1 U521 ( .A1(Set_target[15]), .A2(n3799), .B1(n388), .B2(
        \pc_target[21][15] ), .ZN(n411) );
  INV_X1 U522 ( .A(n412), .ZN(n5834) );
  AOI22_X1 U523 ( .A1(Set_target[17]), .A2(n3799), .B1(n388), .B2(
        \pc_target[21][17] ), .ZN(n412) );
  INV_X1 U524 ( .A(n413), .ZN(n5835) );
  AOI22_X1 U525 ( .A1(Set_target[19]), .A2(n3799), .B1(n388), .B2(
        \pc_target[21][19] ), .ZN(n413) );
  INV_X1 U526 ( .A(n414), .ZN(n5836) );
  AOI22_X1 U527 ( .A1(Set_target[21]), .A2(n3799), .B1(n388), .B2(
        \pc_target[21][21] ), .ZN(n414) );
  INV_X1 U528 ( .A(n415), .ZN(n5837) );
  AOI22_X1 U529 ( .A1(Set_target[23]), .A2(n3799), .B1(n388), .B2(
        \pc_target[21][23] ), .ZN(n415) );
  INV_X1 U530 ( .A(n416), .ZN(n5838) );
  AOI22_X1 U531 ( .A1(Set_target[25]), .A2(n3799), .B1(n388), .B2(
        \pc_target[21][25] ), .ZN(n416) );
  INV_X1 U532 ( .A(n417), .ZN(n5839) );
  AOI22_X1 U533 ( .A1(Set_target[27]), .A2(n3799), .B1(n388), .B2(
        \pc_target[21][27] ), .ZN(n417) );
  INV_X1 U534 ( .A(n418), .ZN(n5840) );
  AOI22_X1 U535 ( .A1(Set_target[29]), .A2(n3799), .B1(n388), .B2(
        \pc_target[21][29] ), .ZN(n418) );
  INV_X1 U536 ( .A(n419), .ZN(n5841) );
  AOI22_X1 U537 ( .A1(Set_target[31]), .A2(n3799), .B1(n388), .B2(
        \pc_target[21][31] ), .ZN(n419) );
  INV_X1 U540 ( .A(n420), .ZN(n5842) );
  AOI22_X1 U541 ( .A1(Set_target[30]), .A2(n421), .B1(n422), .B2(
        \pc_target[20][30] ), .ZN(n420) );
  INV_X1 U542 ( .A(n423), .ZN(n5843) );
  AOI22_X1 U543 ( .A1(Set_target[28]), .A2(n421), .B1(n422), .B2(
        \pc_target[20][28] ), .ZN(n423) );
  INV_X1 U544 ( .A(n424), .ZN(n5844) );
  AOI22_X1 U545 ( .A1(Set_target[26]), .A2(n421), .B1(n422), .B2(
        \pc_target[20][26] ), .ZN(n424) );
  INV_X1 U546 ( .A(n425), .ZN(n5845) );
  AOI22_X1 U547 ( .A1(Set_target[24]), .A2(n421), .B1(n422), .B2(
        \pc_target[20][24] ), .ZN(n425) );
  INV_X1 U548 ( .A(n426), .ZN(n5846) );
  AOI22_X1 U549 ( .A1(Set_target[22]), .A2(n421), .B1(n422), .B2(
        \pc_target[20][22] ), .ZN(n426) );
  INV_X1 U550 ( .A(n427), .ZN(n5847) );
  AOI22_X1 U551 ( .A1(Set_target[20]), .A2(n421), .B1(n422), .B2(
        \pc_target[20][20] ), .ZN(n427) );
  INV_X1 U552 ( .A(n428), .ZN(n5848) );
  AOI22_X1 U553 ( .A1(Set_target[18]), .A2(n421), .B1(n422), .B2(
        \pc_target[20][18] ), .ZN(n428) );
  INV_X1 U554 ( .A(n429), .ZN(n5849) );
  AOI22_X1 U555 ( .A1(Set_target[16]), .A2(n421), .B1(n422), .B2(
        \pc_target[20][16] ), .ZN(n429) );
  INV_X1 U556 ( .A(n430), .ZN(n5850) );
  AOI22_X1 U557 ( .A1(Set_target[14]), .A2(n421), .B1(n422), .B2(
        \pc_target[20][14] ), .ZN(n430) );
  INV_X1 U558 ( .A(n431), .ZN(n5851) );
  AOI22_X1 U559 ( .A1(Set_target[12]), .A2(n421), .B1(n422), .B2(
        \pc_target[20][12] ), .ZN(n431) );
  INV_X1 U560 ( .A(n432), .ZN(n5852) );
  AOI22_X1 U561 ( .A1(Set_target[10]), .A2(n421), .B1(n422), .B2(
        \pc_target[20][10] ), .ZN(n432) );
  INV_X1 U562 ( .A(n433), .ZN(n5853) );
  AOI22_X1 U563 ( .A1(Set_target[8]), .A2(n421), .B1(n422), .B2(
        \pc_target[20][8] ), .ZN(n433) );
  INV_X1 U564 ( .A(n434), .ZN(n5854) );
  AOI22_X1 U565 ( .A1(Set_target[6]), .A2(n421), .B1(n422), .B2(
        \pc_target[20][6] ), .ZN(n434) );
  INV_X1 U566 ( .A(n435), .ZN(n5855) );
  AOI22_X1 U567 ( .A1(Set_target[4]), .A2(n421), .B1(n422), .B2(
        \pc_target[20][4] ), .ZN(n435) );
  INV_X1 U568 ( .A(n436), .ZN(n5856) );
  AOI22_X1 U569 ( .A1(Set_target[2]), .A2(n421), .B1(n422), .B2(
        \pc_target[20][2] ), .ZN(n436) );
  INV_X1 U570 ( .A(n437), .ZN(n5857) );
  AOI22_X1 U571 ( .A1(Set_target[0]), .A2(n421), .B1(n422), .B2(
        \pc_target[20][0] ), .ZN(n437) );
  INV_X1 U572 ( .A(n438), .ZN(n5858) );
  AOI22_X1 U573 ( .A1(Set_target[1]), .A2(n421), .B1(n422), .B2(
        \pc_target[20][1] ), .ZN(n438) );
  INV_X1 U574 ( .A(n439), .ZN(n5859) );
  AOI22_X1 U575 ( .A1(Set_target[3]), .A2(n421), .B1(n422), .B2(
        \pc_target[20][3] ), .ZN(n439) );
  INV_X1 U576 ( .A(n440), .ZN(n5860) );
  AOI22_X1 U577 ( .A1(Set_target[5]), .A2(n421), .B1(n422), .B2(
        \pc_target[20][5] ), .ZN(n440) );
  INV_X1 U578 ( .A(n441), .ZN(n5861) );
  AOI22_X1 U579 ( .A1(Set_target[7]), .A2(n421), .B1(n422), .B2(
        \pc_target[20][7] ), .ZN(n441) );
  INV_X1 U580 ( .A(n442), .ZN(n5862) );
  AOI22_X1 U581 ( .A1(Set_target[9]), .A2(n421), .B1(n422), .B2(
        \pc_target[20][9] ), .ZN(n442) );
  INV_X1 U582 ( .A(n443), .ZN(n5863) );
  AOI22_X1 U583 ( .A1(Set_target[11]), .A2(n421), .B1(n422), .B2(
        \pc_target[20][11] ), .ZN(n443) );
  INV_X1 U584 ( .A(n444), .ZN(n5864) );
  AOI22_X1 U585 ( .A1(Set_target[13]), .A2(n421), .B1(n422), .B2(
        \pc_target[20][13] ), .ZN(n444) );
  INV_X1 U586 ( .A(n445), .ZN(n5865) );
  AOI22_X1 U587 ( .A1(Set_target[15]), .A2(n421), .B1(n422), .B2(
        \pc_target[20][15] ), .ZN(n445) );
  INV_X1 U588 ( .A(n446), .ZN(n5866) );
  AOI22_X1 U589 ( .A1(Set_target[17]), .A2(n421), .B1(n422), .B2(
        \pc_target[20][17] ), .ZN(n446) );
  INV_X1 U590 ( .A(n447), .ZN(n5867) );
  AOI22_X1 U591 ( .A1(Set_target[19]), .A2(n421), .B1(n422), .B2(
        \pc_target[20][19] ), .ZN(n447) );
  INV_X1 U592 ( .A(n448), .ZN(n5868) );
  AOI22_X1 U593 ( .A1(Set_target[21]), .A2(n421), .B1(n422), .B2(
        \pc_target[20][21] ), .ZN(n448) );
  INV_X1 U594 ( .A(n449), .ZN(n5869) );
  AOI22_X1 U595 ( .A1(Set_target[23]), .A2(n421), .B1(n422), .B2(
        \pc_target[20][23] ), .ZN(n449) );
  INV_X1 U596 ( .A(n450), .ZN(n5870) );
  AOI22_X1 U597 ( .A1(Set_target[25]), .A2(n421), .B1(n422), .B2(
        \pc_target[20][25] ), .ZN(n450) );
  INV_X1 U598 ( .A(n451), .ZN(n5871) );
  AOI22_X1 U599 ( .A1(Set_target[27]), .A2(n421), .B1(n422), .B2(
        \pc_target[20][27] ), .ZN(n451) );
  INV_X1 U600 ( .A(n452), .ZN(n5872) );
  AOI22_X1 U601 ( .A1(Set_target[29]), .A2(n421), .B1(n422), .B2(
        \pc_target[20][29] ), .ZN(n452) );
  INV_X1 U602 ( .A(n453), .ZN(n5873) );
  AOI22_X1 U603 ( .A1(Set_target[31]), .A2(n421), .B1(n422), .B2(
        \pc_target[20][31] ), .ZN(n453) );
  INV_X1 U607 ( .A(n455), .ZN(n5874) );
  AOI22_X1 U608 ( .A1(Set_target[30]), .A2(n456), .B1(n457), .B2(
        \pc_target[19][30] ), .ZN(n455) );
  INV_X1 U609 ( .A(n458), .ZN(n5875) );
  AOI22_X1 U610 ( .A1(Set_target[28]), .A2(n456), .B1(n457), .B2(
        \pc_target[19][28] ), .ZN(n458) );
  INV_X1 U611 ( .A(n459), .ZN(n5876) );
  AOI22_X1 U612 ( .A1(Set_target[26]), .A2(n456), .B1(n457), .B2(
        \pc_target[19][26] ), .ZN(n459) );
  INV_X1 U613 ( .A(n460), .ZN(n5877) );
  AOI22_X1 U614 ( .A1(Set_target[24]), .A2(n456), .B1(n457), .B2(
        \pc_target[19][24] ), .ZN(n460) );
  INV_X1 U615 ( .A(n461), .ZN(n5878) );
  AOI22_X1 U616 ( .A1(Set_target[22]), .A2(n456), .B1(n457), .B2(
        \pc_target[19][22] ), .ZN(n461) );
  INV_X1 U617 ( .A(n462), .ZN(n5879) );
  AOI22_X1 U618 ( .A1(Set_target[20]), .A2(n456), .B1(n457), .B2(
        \pc_target[19][20] ), .ZN(n462) );
  INV_X1 U619 ( .A(n463), .ZN(n5880) );
  AOI22_X1 U620 ( .A1(Set_target[18]), .A2(n456), .B1(n457), .B2(
        \pc_target[19][18] ), .ZN(n463) );
  INV_X1 U621 ( .A(n464), .ZN(n5881) );
  AOI22_X1 U622 ( .A1(Set_target[16]), .A2(n456), .B1(n457), .B2(
        \pc_target[19][16] ), .ZN(n464) );
  INV_X1 U623 ( .A(n465), .ZN(n5882) );
  AOI22_X1 U624 ( .A1(Set_target[14]), .A2(n456), .B1(n457), .B2(
        \pc_target[19][14] ), .ZN(n465) );
  INV_X1 U625 ( .A(n466), .ZN(n5883) );
  AOI22_X1 U626 ( .A1(Set_target[12]), .A2(n456), .B1(n457), .B2(
        \pc_target[19][12] ), .ZN(n466) );
  INV_X1 U627 ( .A(n467), .ZN(n5884) );
  AOI22_X1 U628 ( .A1(Set_target[10]), .A2(n456), .B1(n457), .B2(
        \pc_target[19][10] ), .ZN(n467) );
  INV_X1 U629 ( .A(n468), .ZN(n5885) );
  AOI22_X1 U630 ( .A1(Set_target[8]), .A2(n456), .B1(n457), .B2(
        \pc_target[19][8] ), .ZN(n468) );
  INV_X1 U631 ( .A(n469), .ZN(n5886) );
  AOI22_X1 U632 ( .A1(Set_target[6]), .A2(n456), .B1(n457), .B2(
        \pc_target[19][6] ), .ZN(n469) );
  INV_X1 U633 ( .A(n470), .ZN(n5887) );
  AOI22_X1 U634 ( .A1(Set_target[4]), .A2(n456), .B1(n457), .B2(
        \pc_target[19][4] ), .ZN(n470) );
  INV_X1 U635 ( .A(n471), .ZN(n5888) );
  AOI22_X1 U636 ( .A1(Set_target[2]), .A2(n456), .B1(n457), .B2(
        \pc_target[19][2] ), .ZN(n471) );
  INV_X1 U637 ( .A(n472), .ZN(n5889) );
  AOI22_X1 U638 ( .A1(Set_target[0]), .A2(n456), .B1(n457), .B2(
        \pc_target[19][0] ), .ZN(n472) );
  INV_X1 U639 ( .A(n473), .ZN(n5890) );
  AOI22_X1 U640 ( .A1(Set_target[1]), .A2(n456), .B1(n457), .B2(
        \pc_target[19][1] ), .ZN(n473) );
  INV_X1 U641 ( .A(n474), .ZN(n5891) );
  AOI22_X1 U642 ( .A1(Set_target[3]), .A2(n456), .B1(n457), .B2(
        \pc_target[19][3] ), .ZN(n474) );
  INV_X1 U643 ( .A(n475), .ZN(n5892) );
  AOI22_X1 U644 ( .A1(Set_target[5]), .A2(n456), .B1(n457), .B2(
        \pc_target[19][5] ), .ZN(n475) );
  INV_X1 U645 ( .A(n476), .ZN(n5893) );
  AOI22_X1 U646 ( .A1(Set_target[7]), .A2(n456), .B1(n457), .B2(
        \pc_target[19][7] ), .ZN(n476) );
  INV_X1 U647 ( .A(n477), .ZN(n5894) );
  AOI22_X1 U648 ( .A1(Set_target[9]), .A2(n456), .B1(n457), .B2(
        \pc_target[19][9] ), .ZN(n477) );
  INV_X1 U649 ( .A(n478), .ZN(n5895) );
  AOI22_X1 U650 ( .A1(Set_target[11]), .A2(n456), .B1(n457), .B2(
        \pc_target[19][11] ), .ZN(n478) );
  INV_X1 U651 ( .A(n479), .ZN(n5896) );
  AOI22_X1 U652 ( .A1(Set_target[13]), .A2(n456), .B1(n457), .B2(
        \pc_target[19][13] ), .ZN(n479) );
  INV_X1 U653 ( .A(n480), .ZN(n5897) );
  AOI22_X1 U654 ( .A1(Set_target[15]), .A2(n456), .B1(n457), .B2(
        \pc_target[19][15] ), .ZN(n480) );
  INV_X1 U655 ( .A(n481), .ZN(n5898) );
  AOI22_X1 U656 ( .A1(Set_target[17]), .A2(n456), .B1(n457), .B2(
        \pc_target[19][17] ), .ZN(n481) );
  INV_X1 U657 ( .A(n482), .ZN(n5899) );
  AOI22_X1 U658 ( .A1(Set_target[19]), .A2(n456), .B1(n457), .B2(
        \pc_target[19][19] ), .ZN(n482) );
  INV_X1 U659 ( .A(n483), .ZN(n5900) );
  AOI22_X1 U660 ( .A1(Set_target[21]), .A2(n456), .B1(n457), .B2(
        \pc_target[19][21] ), .ZN(n483) );
  INV_X1 U661 ( .A(n484), .ZN(n5901) );
  AOI22_X1 U662 ( .A1(Set_target[23]), .A2(n456), .B1(n457), .B2(
        \pc_target[19][23] ), .ZN(n484) );
  INV_X1 U663 ( .A(n485), .ZN(n5902) );
  AOI22_X1 U664 ( .A1(Set_target[25]), .A2(n456), .B1(n457), .B2(
        \pc_target[19][25] ), .ZN(n485) );
  INV_X1 U665 ( .A(n486), .ZN(n5903) );
  AOI22_X1 U666 ( .A1(Set_target[27]), .A2(n456), .B1(n457), .B2(
        \pc_target[19][27] ), .ZN(n486) );
  INV_X1 U667 ( .A(n487), .ZN(n5904) );
  AOI22_X1 U668 ( .A1(Set_target[29]), .A2(n456), .B1(n457), .B2(
        \pc_target[19][29] ), .ZN(n487) );
  INV_X1 U669 ( .A(n488), .ZN(n5905) );
  AOI22_X1 U670 ( .A1(Set_target[31]), .A2(n456), .B1(n457), .B2(
        \pc_target[19][31] ), .ZN(n488) );
  INV_X1 U673 ( .A(n490), .ZN(n5906) );
  AOI22_X1 U674 ( .A1(Set_target[30]), .A2(n491), .B1(n492), .B2(
        \pc_target[18][30] ), .ZN(n490) );
  INV_X1 U675 ( .A(n493), .ZN(n5907) );
  AOI22_X1 U676 ( .A1(Set_target[28]), .A2(n491), .B1(n492), .B2(
        \pc_target[18][28] ), .ZN(n493) );
  INV_X1 U677 ( .A(n494), .ZN(n5908) );
  AOI22_X1 U678 ( .A1(Set_target[26]), .A2(n491), .B1(n492), .B2(
        \pc_target[18][26] ), .ZN(n494) );
  INV_X1 U679 ( .A(n495), .ZN(n5909) );
  AOI22_X1 U680 ( .A1(Set_target[24]), .A2(n491), .B1(n492), .B2(
        \pc_target[18][24] ), .ZN(n495) );
  INV_X1 U681 ( .A(n496), .ZN(n5910) );
  AOI22_X1 U682 ( .A1(Set_target[22]), .A2(n491), .B1(n492), .B2(
        \pc_target[18][22] ), .ZN(n496) );
  INV_X1 U683 ( .A(n497), .ZN(n5911) );
  AOI22_X1 U684 ( .A1(Set_target[20]), .A2(n491), .B1(n492), .B2(
        \pc_target[18][20] ), .ZN(n497) );
  INV_X1 U685 ( .A(n498), .ZN(n5912) );
  AOI22_X1 U686 ( .A1(Set_target[18]), .A2(n491), .B1(n492), .B2(
        \pc_target[18][18] ), .ZN(n498) );
  INV_X1 U687 ( .A(n499), .ZN(n5913) );
  AOI22_X1 U688 ( .A1(Set_target[16]), .A2(n491), .B1(n492), .B2(
        \pc_target[18][16] ), .ZN(n499) );
  INV_X1 U689 ( .A(n500), .ZN(n5914) );
  AOI22_X1 U690 ( .A1(Set_target[14]), .A2(n491), .B1(n492), .B2(
        \pc_target[18][14] ), .ZN(n500) );
  INV_X1 U691 ( .A(n501), .ZN(n5915) );
  AOI22_X1 U692 ( .A1(Set_target[12]), .A2(n491), .B1(n492), .B2(
        \pc_target[18][12] ), .ZN(n501) );
  INV_X1 U693 ( .A(n502), .ZN(n5916) );
  AOI22_X1 U694 ( .A1(Set_target[10]), .A2(n491), .B1(n492), .B2(
        \pc_target[18][10] ), .ZN(n502) );
  INV_X1 U695 ( .A(n503), .ZN(n5917) );
  AOI22_X1 U696 ( .A1(Set_target[8]), .A2(n491), .B1(n492), .B2(
        \pc_target[18][8] ), .ZN(n503) );
  INV_X1 U697 ( .A(n504), .ZN(n5918) );
  AOI22_X1 U698 ( .A1(Set_target[6]), .A2(n491), .B1(n492), .B2(
        \pc_target[18][6] ), .ZN(n504) );
  INV_X1 U699 ( .A(n505), .ZN(n5919) );
  AOI22_X1 U700 ( .A1(Set_target[4]), .A2(n491), .B1(n492), .B2(
        \pc_target[18][4] ), .ZN(n505) );
  INV_X1 U701 ( .A(n506), .ZN(n5920) );
  AOI22_X1 U702 ( .A1(Set_target[2]), .A2(n491), .B1(n492), .B2(
        \pc_target[18][2] ), .ZN(n506) );
  INV_X1 U703 ( .A(n507), .ZN(n5921) );
  AOI22_X1 U704 ( .A1(Set_target[0]), .A2(n491), .B1(n492), .B2(
        \pc_target[18][0] ), .ZN(n507) );
  INV_X1 U705 ( .A(n508), .ZN(n5922) );
  AOI22_X1 U706 ( .A1(Set_target[1]), .A2(n491), .B1(n492), .B2(
        \pc_target[18][1] ), .ZN(n508) );
  INV_X1 U707 ( .A(n509), .ZN(n5923) );
  AOI22_X1 U708 ( .A1(Set_target[3]), .A2(n491), .B1(n492), .B2(
        \pc_target[18][3] ), .ZN(n509) );
  INV_X1 U709 ( .A(n510), .ZN(n5924) );
  AOI22_X1 U710 ( .A1(Set_target[5]), .A2(n491), .B1(n492), .B2(
        \pc_target[18][5] ), .ZN(n510) );
  INV_X1 U711 ( .A(n511), .ZN(n5925) );
  AOI22_X1 U712 ( .A1(Set_target[7]), .A2(n491), .B1(n492), .B2(
        \pc_target[18][7] ), .ZN(n511) );
  INV_X1 U713 ( .A(n512), .ZN(n5926) );
  AOI22_X1 U714 ( .A1(Set_target[9]), .A2(n491), .B1(n492), .B2(
        \pc_target[18][9] ), .ZN(n512) );
  INV_X1 U715 ( .A(n513), .ZN(n5927) );
  AOI22_X1 U716 ( .A1(Set_target[11]), .A2(n491), .B1(n492), .B2(
        \pc_target[18][11] ), .ZN(n513) );
  INV_X1 U717 ( .A(n514), .ZN(n5928) );
  AOI22_X1 U718 ( .A1(Set_target[13]), .A2(n491), .B1(n492), .B2(
        \pc_target[18][13] ), .ZN(n514) );
  INV_X1 U719 ( .A(n515), .ZN(n5929) );
  AOI22_X1 U720 ( .A1(Set_target[15]), .A2(n491), .B1(n492), .B2(
        \pc_target[18][15] ), .ZN(n515) );
  INV_X1 U721 ( .A(n516), .ZN(n5930) );
  AOI22_X1 U722 ( .A1(Set_target[17]), .A2(n491), .B1(n492), .B2(
        \pc_target[18][17] ), .ZN(n516) );
  INV_X1 U723 ( .A(n517), .ZN(n5931) );
  AOI22_X1 U724 ( .A1(Set_target[19]), .A2(n491), .B1(n492), .B2(
        \pc_target[18][19] ), .ZN(n517) );
  INV_X1 U725 ( .A(n518), .ZN(n5932) );
  AOI22_X1 U726 ( .A1(Set_target[21]), .A2(n491), .B1(n492), .B2(
        \pc_target[18][21] ), .ZN(n518) );
  INV_X1 U727 ( .A(n519), .ZN(n5933) );
  AOI22_X1 U728 ( .A1(Set_target[23]), .A2(n491), .B1(n492), .B2(
        \pc_target[18][23] ), .ZN(n519) );
  INV_X1 U729 ( .A(n520), .ZN(n5934) );
  AOI22_X1 U730 ( .A1(Set_target[25]), .A2(n491), .B1(n492), .B2(
        \pc_target[18][25] ), .ZN(n520) );
  INV_X1 U731 ( .A(n521), .ZN(n5935) );
  AOI22_X1 U732 ( .A1(Set_target[27]), .A2(n491), .B1(n492), .B2(
        \pc_target[18][27] ), .ZN(n521) );
  INV_X1 U733 ( .A(n522), .ZN(n5936) );
  AOI22_X1 U734 ( .A1(Set_target[29]), .A2(n491), .B1(n492), .B2(
        \pc_target[18][29] ), .ZN(n522) );
  INV_X1 U735 ( .A(n523), .ZN(n5937) );
  AOI22_X1 U736 ( .A1(Set_target[31]), .A2(n491), .B1(n492), .B2(
        \pc_target[18][31] ), .ZN(n523) );
  OAI22_X1 U739 ( .A1(n75), .A2(n524), .B1(n3445), .B2(n526), .ZN(n5938) );
  OAI22_X1 U740 ( .A1(n79), .A2(n524), .B1(n3445), .B2(n527), .ZN(n5939) );
  OAI22_X1 U741 ( .A1(n81), .A2(n524), .B1(n3445), .B2(n528), .ZN(n5940) );
  OAI22_X1 U742 ( .A1(n83), .A2(n524), .B1(n3445), .B2(n529), .ZN(n5941) );
  OAI22_X1 U743 ( .A1(n85), .A2(n524), .B1(n3445), .B2(n530), .ZN(n5942) );
  OAI22_X1 U744 ( .A1(n87), .A2(n524), .B1(n3445), .B2(n531), .ZN(n5943) );
  OAI22_X1 U745 ( .A1(n89), .A2(n524), .B1(n3445), .B2(n532), .ZN(n5944) );
  OAI22_X1 U746 ( .A1(n91), .A2(n524), .B1(n3445), .B2(n533), .ZN(n5945) );
  OAI22_X1 U747 ( .A1(n93), .A2(n524), .B1(n3445), .B2(n534), .ZN(n5946) );
  OAI22_X1 U748 ( .A1(n95), .A2(n524), .B1(n3445), .B2(n535), .ZN(n5947) );
  OAI22_X1 U749 ( .A1(n97), .A2(n524), .B1(n3445), .B2(n536), .ZN(n5948) );
  OAI22_X1 U750 ( .A1(n99), .A2(n524), .B1(n3445), .B2(n537), .ZN(n5949) );
  OAI22_X1 U751 ( .A1(n101), .A2(n524), .B1(n3445), .B2(n538), .ZN(n5950) );
  OAI22_X1 U752 ( .A1(n103), .A2(n524), .B1(n3445), .B2(n539), .ZN(n5951) );
  OAI22_X1 U753 ( .A1(n105), .A2(n524), .B1(n3445), .B2(n540), .ZN(n5952) );
  OAI22_X1 U754 ( .A1(n107), .A2(n524), .B1(n3445), .B2(n541), .ZN(n5953) );
  OAI22_X1 U755 ( .A1(n109), .A2(n524), .B1(n3445), .B2(n542), .ZN(n5954) );
  OAI22_X1 U756 ( .A1(n111), .A2(n524), .B1(n3445), .B2(n543), .ZN(n5955) );
  OAI22_X1 U757 ( .A1(n113), .A2(n524), .B1(n3445), .B2(n544), .ZN(n5956) );
  OAI22_X1 U758 ( .A1(n115), .A2(n524), .B1(n3445), .B2(n545), .ZN(n5957) );
  OAI22_X1 U759 ( .A1(n117), .A2(n524), .B1(n3445), .B2(n546), .ZN(n5958) );
  OAI22_X1 U760 ( .A1(n119), .A2(n524), .B1(n3445), .B2(n547), .ZN(n5959) );
  OAI22_X1 U761 ( .A1(n121), .A2(n524), .B1(n3445), .B2(n548), .ZN(n5960) );
  OAI22_X1 U762 ( .A1(n123), .A2(n524), .B1(n3445), .B2(n549), .ZN(n5961) );
  OAI22_X1 U763 ( .A1(n125), .A2(n524), .B1(n3445), .B2(n550), .ZN(n5962) );
  OAI22_X1 U764 ( .A1(n127), .A2(n524), .B1(n3445), .B2(n551), .ZN(n5963) );
  OAI22_X1 U765 ( .A1(n129), .A2(n524), .B1(n3445), .B2(n552), .ZN(n5964) );
  OAI22_X1 U766 ( .A1(n131), .A2(n524), .B1(n3445), .B2(n553), .ZN(n5965) );
  OAI22_X1 U767 ( .A1(n133), .A2(n524), .B1(n3445), .B2(n554), .ZN(n5966) );
  OAI22_X1 U768 ( .A1(n135), .A2(n524), .B1(n3445), .B2(n555), .ZN(n5967) );
  OAI22_X1 U769 ( .A1(n137), .A2(n524), .B1(n3445), .B2(n556), .ZN(n5968) );
  OAI22_X1 U770 ( .A1(n139), .A2(n524), .B1(n3445), .B2(n557), .ZN(n5969) );
  OAI22_X1 U773 ( .A1(n75), .A2(n1463), .B1(n559), .B2(n560), .ZN(n5970) );
  OAI22_X1 U774 ( .A1(n79), .A2(n1481), .B1(n559), .B2(n561), .ZN(n5971) );
  OAI22_X1 U775 ( .A1(n81), .A2(n1481), .B1(n559), .B2(n562), .ZN(n5972) );
  OAI22_X1 U776 ( .A1(n83), .A2(n1481), .B1(n559), .B2(n563), .ZN(n5973) );
  OAI22_X1 U778 ( .A1(n87), .A2(n1463), .B1(n559), .B2(n565), .ZN(n5975) );
  OAI22_X1 U779 ( .A1(n89), .A2(n1481), .B1(n559), .B2(n566), .ZN(n5976) );
  OAI22_X1 U780 ( .A1(n91), .A2(n1463), .B1(n559), .B2(n567), .ZN(n5977) );
  OAI22_X1 U781 ( .A1(n93), .A2(n1481), .B1(n559), .B2(n568), .ZN(n5978) );
  OAI22_X1 U782 ( .A1(n95), .A2(n1463), .B1(n559), .B2(n569), .ZN(n5979) );
  OAI22_X1 U783 ( .A1(n97), .A2(n1481), .B1(n559), .B2(n570), .ZN(n5980) );
  OAI22_X1 U784 ( .A1(n99), .A2(n1481), .B1(n559), .B2(n571), .ZN(n5981) );
  OAI22_X1 U785 ( .A1(n101), .A2(n1481), .B1(n559), .B2(n572), .ZN(n5982) );
  OAI22_X1 U786 ( .A1(n103), .A2(n1481), .B1(n559), .B2(n573), .ZN(n5983) );
  OAI22_X1 U787 ( .A1(n105), .A2(n1481), .B1(n559), .B2(n574), .ZN(n5984) );
  OAI22_X1 U788 ( .A1(n107), .A2(n1481), .B1(n559), .B2(n575), .ZN(n5985) );
  OAI22_X1 U789 ( .A1(n109), .A2(n1481), .B1(n559), .B2(n576), .ZN(n5986) );
  OAI22_X1 U790 ( .A1(n111), .A2(n1481), .B1(n559), .B2(n577), .ZN(n5987) );
  OAI22_X1 U791 ( .A1(n113), .A2(n1481), .B1(n559), .B2(n578), .ZN(n5988) );
  OAI22_X1 U792 ( .A1(n115), .A2(n1481), .B1(n559), .B2(n579), .ZN(n5989) );
  OAI22_X1 U793 ( .A1(n117), .A2(n1481), .B1(n559), .B2(n580), .ZN(n5990) );
  OAI22_X1 U794 ( .A1(n119), .A2(n1481), .B1(n559), .B2(n581), .ZN(n5991) );
  OAI22_X1 U795 ( .A1(n121), .A2(n1481), .B1(n559), .B2(n582), .ZN(n5992) );
  OAI22_X1 U796 ( .A1(n123), .A2(n1481), .B1(n559), .B2(n583), .ZN(n5993) );
  OAI22_X1 U797 ( .A1(n125), .A2(n1481), .B1(n559), .B2(n584), .ZN(n5994) );
  OAI22_X1 U798 ( .A1(n127), .A2(n1481), .B1(n559), .B2(n585), .ZN(n5995) );
  OAI22_X1 U799 ( .A1(n129), .A2(n1481), .B1(n559), .B2(n586), .ZN(n5996) );
  OAI22_X1 U800 ( .A1(n131), .A2(n1481), .B1(n559), .B2(n587), .ZN(n5997) );
  OAI22_X1 U801 ( .A1(n133), .A2(n1481), .B1(n559), .B2(n588), .ZN(n5998) );
  OAI22_X1 U802 ( .A1(n135), .A2(n1463), .B1(n559), .B2(n589), .ZN(n5999) );
  OAI22_X1 U803 ( .A1(n137), .A2(n1481), .B1(n559), .B2(n590), .ZN(n6000) );
  OAI22_X1 U804 ( .A1(n139), .A2(n1481), .B1(n559), .B2(n591), .ZN(n6001) );
  INV_X1 U809 ( .A(n594), .ZN(n6002) );
  AOI22_X1 U810 ( .A1(Set_target[30]), .A2(n595), .B1(n596), .B2(
        \pc_target[15][30] ), .ZN(n594) );
  INV_X1 U811 ( .A(n597), .ZN(n6003) );
  AOI22_X1 U812 ( .A1(Set_target[28]), .A2(n595), .B1(n596), .B2(
        \pc_target[15][28] ), .ZN(n597) );
  INV_X1 U813 ( .A(n598), .ZN(n6004) );
  AOI22_X1 U814 ( .A1(Set_target[26]), .A2(n595), .B1(n596), .B2(
        \pc_target[15][26] ), .ZN(n598) );
  INV_X1 U815 ( .A(n599), .ZN(n6005) );
  AOI22_X1 U816 ( .A1(Set_target[24]), .A2(n595), .B1(n596), .B2(
        \pc_target[15][24] ), .ZN(n599) );
  INV_X1 U817 ( .A(n600), .ZN(n6006) );
  AOI22_X1 U818 ( .A1(Set_target[22]), .A2(n595), .B1(n596), .B2(
        \pc_target[15][22] ), .ZN(n600) );
  INV_X1 U819 ( .A(n601), .ZN(n6007) );
  AOI22_X1 U820 ( .A1(Set_target[20]), .A2(n595), .B1(n596), .B2(
        \pc_target[15][20] ), .ZN(n601) );
  INV_X1 U821 ( .A(n602), .ZN(n6008) );
  AOI22_X1 U822 ( .A1(Set_target[18]), .A2(n595), .B1(n596), .B2(
        \pc_target[15][18] ), .ZN(n602) );
  INV_X1 U823 ( .A(n603), .ZN(n6009) );
  AOI22_X1 U824 ( .A1(Set_target[16]), .A2(n595), .B1(n596), .B2(
        \pc_target[15][16] ), .ZN(n603) );
  INV_X1 U825 ( .A(n604), .ZN(n6010) );
  AOI22_X1 U826 ( .A1(Set_target[14]), .A2(n595), .B1(n596), .B2(
        \pc_target[15][14] ), .ZN(n604) );
  INV_X1 U827 ( .A(n605), .ZN(n6011) );
  AOI22_X1 U828 ( .A1(Set_target[12]), .A2(n595), .B1(n596), .B2(
        \pc_target[15][12] ), .ZN(n605) );
  INV_X1 U829 ( .A(n606), .ZN(n6012) );
  AOI22_X1 U830 ( .A1(Set_target[10]), .A2(n595), .B1(n596), .B2(
        \pc_target[15][10] ), .ZN(n606) );
  INV_X1 U831 ( .A(n607), .ZN(n6013) );
  AOI22_X1 U832 ( .A1(Set_target[8]), .A2(n595), .B1(n596), .B2(
        \pc_target[15][8] ), .ZN(n607) );
  INV_X1 U833 ( .A(n608), .ZN(n6014) );
  AOI22_X1 U834 ( .A1(Set_target[6]), .A2(n595), .B1(n596), .B2(
        \pc_target[15][6] ), .ZN(n608) );
  INV_X1 U835 ( .A(n609), .ZN(n6015) );
  AOI22_X1 U836 ( .A1(Set_target[4]), .A2(n595), .B1(n596), .B2(
        \pc_target[15][4] ), .ZN(n609) );
  INV_X1 U837 ( .A(n610), .ZN(n6016) );
  AOI22_X1 U838 ( .A1(Set_target[2]), .A2(n595), .B1(n596), .B2(
        \pc_target[15][2] ), .ZN(n610) );
  INV_X1 U839 ( .A(n611), .ZN(n6017) );
  AOI22_X1 U840 ( .A1(Set_target[0]), .A2(n595), .B1(n596), .B2(
        \pc_target[15][0] ), .ZN(n611) );
  INV_X1 U841 ( .A(n612), .ZN(n6018) );
  AOI22_X1 U842 ( .A1(Set_target[1]), .A2(n595), .B1(n596), .B2(
        \pc_target[15][1] ), .ZN(n612) );
  INV_X1 U843 ( .A(n613), .ZN(n6019) );
  AOI22_X1 U844 ( .A1(Set_target[3]), .A2(n595), .B1(n596), .B2(
        \pc_target[15][3] ), .ZN(n613) );
  INV_X1 U845 ( .A(n614), .ZN(n6020) );
  AOI22_X1 U846 ( .A1(Set_target[5]), .A2(n595), .B1(n596), .B2(
        \pc_target[15][5] ), .ZN(n614) );
  INV_X1 U847 ( .A(n615), .ZN(n6021) );
  AOI22_X1 U848 ( .A1(Set_target[7]), .A2(n595), .B1(n596), .B2(
        \pc_target[15][7] ), .ZN(n615) );
  INV_X1 U849 ( .A(n616), .ZN(n6022) );
  AOI22_X1 U850 ( .A1(Set_target[9]), .A2(n595), .B1(n596), .B2(
        \pc_target[15][9] ), .ZN(n616) );
  INV_X1 U851 ( .A(n617), .ZN(n6023) );
  AOI22_X1 U852 ( .A1(Set_target[11]), .A2(n595), .B1(n596), .B2(
        \pc_target[15][11] ), .ZN(n617) );
  INV_X1 U853 ( .A(n618), .ZN(n6024) );
  AOI22_X1 U854 ( .A1(Set_target[13]), .A2(n595), .B1(n596), .B2(
        \pc_target[15][13] ), .ZN(n618) );
  INV_X1 U855 ( .A(n619), .ZN(n6025) );
  AOI22_X1 U856 ( .A1(Set_target[15]), .A2(n595), .B1(n596), .B2(
        \pc_target[15][15] ), .ZN(n619) );
  INV_X1 U857 ( .A(n620), .ZN(n6026) );
  AOI22_X1 U858 ( .A1(Set_target[17]), .A2(n595), .B1(n596), .B2(
        \pc_target[15][17] ), .ZN(n620) );
  INV_X1 U859 ( .A(n621), .ZN(n6027) );
  AOI22_X1 U860 ( .A1(Set_target[19]), .A2(n595), .B1(n596), .B2(
        \pc_target[15][19] ), .ZN(n621) );
  INV_X1 U861 ( .A(n622), .ZN(n6028) );
  AOI22_X1 U862 ( .A1(Set_target[21]), .A2(n595), .B1(n596), .B2(
        \pc_target[15][21] ), .ZN(n622) );
  INV_X1 U863 ( .A(n623), .ZN(n6029) );
  AOI22_X1 U864 ( .A1(Set_target[23]), .A2(n595), .B1(n596), .B2(
        \pc_target[15][23] ), .ZN(n623) );
  INV_X1 U865 ( .A(n624), .ZN(n6030) );
  AOI22_X1 U866 ( .A1(Set_target[25]), .A2(n595), .B1(n596), .B2(
        \pc_target[15][25] ), .ZN(n624) );
  INV_X1 U867 ( .A(n625), .ZN(n6031) );
  AOI22_X1 U868 ( .A1(Set_target[27]), .A2(n595), .B1(n596), .B2(
        \pc_target[15][27] ), .ZN(n625) );
  INV_X1 U869 ( .A(n626), .ZN(n6032) );
  AOI22_X1 U870 ( .A1(Set_target[29]), .A2(n595), .B1(n596), .B2(
        \pc_target[15][29] ), .ZN(n626) );
  INV_X1 U871 ( .A(n627), .ZN(n6033) );
  AOI22_X1 U872 ( .A1(Set_target[31]), .A2(n595), .B1(n596), .B2(
        \pc_target[15][31] ), .ZN(n627) );
  INV_X1 U875 ( .A(n629), .ZN(n6034) );
  AOI22_X1 U876 ( .A1(Set_target[30]), .A2(n630), .B1(n631), .B2(
        \pc_target[14][30] ), .ZN(n629) );
  INV_X1 U877 ( .A(n632), .ZN(n6035) );
  AOI22_X1 U878 ( .A1(Set_target[28]), .A2(n630), .B1(n631), .B2(
        \pc_target[14][28] ), .ZN(n632) );
  INV_X1 U879 ( .A(n633), .ZN(n6036) );
  AOI22_X1 U880 ( .A1(Set_target[26]), .A2(n630), .B1(n631), .B2(
        \pc_target[14][26] ), .ZN(n633) );
  INV_X1 U881 ( .A(n634), .ZN(n6037) );
  AOI22_X1 U882 ( .A1(Set_target[24]), .A2(n630), .B1(n631), .B2(
        \pc_target[14][24] ), .ZN(n634) );
  INV_X1 U883 ( .A(n635), .ZN(n6038) );
  AOI22_X1 U884 ( .A1(Set_target[22]), .A2(n630), .B1(n631), .B2(
        \pc_target[14][22] ), .ZN(n635) );
  INV_X1 U885 ( .A(n636), .ZN(n6039) );
  AOI22_X1 U886 ( .A1(Set_target[20]), .A2(n630), .B1(n631), .B2(
        \pc_target[14][20] ), .ZN(n636) );
  INV_X1 U887 ( .A(n637), .ZN(n6040) );
  AOI22_X1 U888 ( .A1(Set_target[18]), .A2(n630), .B1(n631), .B2(
        \pc_target[14][18] ), .ZN(n637) );
  INV_X1 U889 ( .A(n638), .ZN(n6041) );
  AOI22_X1 U890 ( .A1(Set_target[16]), .A2(n630), .B1(n631), .B2(
        \pc_target[14][16] ), .ZN(n638) );
  INV_X1 U891 ( .A(n639), .ZN(n6042) );
  AOI22_X1 U892 ( .A1(Set_target[14]), .A2(n630), .B1(n631), .B2(
        \pc_target[14][14] ), .ZN(n639) );
  INV_X1 U893 ( .A(n640), .ZN(n6043) );
  AOI22_X1 U894 ( .A1(Set_target[12]), .A2(n630), .B1(n631), .B2(
        \pc_target[14][12] ), .ZN(n640) );
  INV_X1 U895 ( .A(n641), .ZN(n6044) );
  AOI22_X1 U896 ( .A1(Set_target[10]), .A2(n630), .B1(n631), .B2(
        \pc_target[14][10] ), .ZN(n641) );
  INV_X1 U897 ( .A(n642), .ZN(n6045) );
  AOI22_X1 U898 ( .A1(Set_target[8]), .A2(n630), .B1(n631), .B2(
        \pc_target[14][8] ), .ZN(n642) );
  INV_X1 U899 ( .A(n643), .ZN(n6046) );
  AOI22_X1 U900 ( .A1(Set_target[6]), .A2(n630), .B1(n631), .B2(
        \pc_target[14][6] ), .ZN(n643) );
  INV_X1 U901 ( .A(n644), .ZN(n6047) );
  AOI22_X1 U902 ( .A1(Set_target[4]), .A2(n630), .B1(n631), .B2(
        \pc_target[14][4] ), .ZN(n644) );
  INV_X1 U903 ( .A(n645), .ZN(n6048) );
  AOI22_X1 U904 ( .A1(Set_target[2]), .A2(n630), .B1(n631), .B2(
        \pc_target[14][2] ), .ZN(n645) );
  INV_X1 U905 ( .A(n646), .ZN(n6049) );
  AOI22_X1 U906 ( .A1(Set_target[0]), .A2(n630), .B1(n631), .B2(
        \pc_target[14][0] ), .ZN(n646) );
  INV_X1 U907 ( .A(n647), .ZN(n6050) );
  AOI22_X1 U908 ( .A1(Set_target[1]), .A2(n630), .B1(n631), .B2(
        \pc_target[14][1] ), .ZN(n647) );
  INV_X1 U909 ( .A(n648), .ZN(n6051) );
  AOI22_X1 U910 ( .A1(Set_target[3]), .A2(n630), .B1(n631), .B2(
        \pc_target[14][3] ), .ZN(n648) );
  INV_X1 U911 ( .A(n649), .ZN(n6052) );
  AOI22_X1 U912 ( .A1(Set_target[5]), .A2(n630), .B1(n631), .B2(
        \pc_target[14][5] ), .ZN(n649) );
  INV_X1 U913 ( .A(n650), .ZN(n6053) );
  AOI22_X1 U914 ( .A1(Set_target[7]), .A2(n630), .B1(n631), .B2(
        \pc_target[14][7] ), .ZN(n650) );
  INV_X1 U915 ( .A(n651), .ZN(n6054) );
  AOI22_X1 U916 ( .A1(Set_target[9]), .A2(n630), .B1(n631), .B2(
        \pc_target[14][9] ), .ZN(n651) );
  INV_X1 U917 ( .A(n652), .ZN(n6055) );
  AOI22_X1 U918 ( .A1(Set_target[11]), .A2(n630), .B1(n631), .B2(
        \pc_target[14][11] ), .ZN(n652) );
  INV_X1 U919 ( .A(n653), .ZN(n6056) );
  AOI22_X1 U920 ( .A1(Set_target[13]), .A2(n630), .B1(n631), .B2(
        \pc_target[14][13] ), .ZN(n653) );
  INV_X1 U921 ( .A(n654), .ZN(n6057) );
  AOI22_X1 U922 ( .A1(Set_target[15]), .A2(n630), .B1(n631), .B2(
        \pc_target[14][15] ), .ZN(n654) );
  INV_X1 U923 ( .A(n655), .ZN(n6058) );
  AOI22_X1 U924 ( .A1(Set_target[17]), .A2(n630), .B1(n631), .B2(
        \pc_target[14][17] ), .ZN(n655) );
  INV_X1 U925 ( .A(n656), .ZN(n6059) );
  AOI22_X1 U926 ( .A1(Set_target[19]), .A2(n630), .B1(n631), .B2(
        \pc_target[14][19] ), .ZN(n656) );
  INV_X1 U927 ( .A(n657), .ZN(n6060) );
  AOI22_X1 U928 ( .A1(Set_target[21]), .A2(n630), .B1(n631), .B2(
        \pc_target[14][21] ), .ZN(n657) );
  INV_X1 U929 ( .A(n658), .ZN(n6061) );
  AOI22_X1 U930 ( .A1(Set_target[23]), .A2(n630), .B1(n631), .B2(
        \pc_target[14][23] ), .ZN(n658) );
  INV_X1 U931 ( .A(n659), .ZN(n6062) );
  AOI22_X1 U932 ( .A1(Set_target[25]), .A2(n630), .B1(n631), .B2(
        \pc_target[14][25] ), .ZN(n659) );
  INV_X1 U933 ( .A(n660), .ZN(n6063) );
  AOI22_X1 U934 ( .A1(Set_target[27]), .A2(n630), .B1(n631), .B2(
        \pc_target[14][27] ), .ZN(n660) );
  INV_X1 U935 ( .A(n661), .ZN(n6064) );
  AOI22_X1 U936 ( .A1(Set_target[29]), .A2(n630), .B1(n631), .B2(
        \pc_target[14][29] ), .ZN(n661) );
  INV_X1 U937 ( .A(n662), .ZN(n6065) );
  AOI22_X1 U938 ( .A1(Set_target[31]), .A2(n630), .B1(n631), .B2(
        \pc_target[14][31] ), .ZN(n662) );
  OAI22_X1 U941 ( .A1(n75), .A2(n663), .B1(n664), .B2(n665), .ZN(n6066) );
  OAI22_X1 U942 ( .A1(n79), .A2(n663), .B1(n664), .B2(n666), .ZN(n6067) );
  OAI22_X1 U943 ( .A1(n81), .A2(n663), .B1(n664), .B2(n667), .ZN(n6068) );
  OAI22_X1 U944 ( .A1(n83), .A2(n663), .B1(n664), .B2(n668), .ZN(n6069) );
  OAI22_X1 U945 ( .A1(n85), .A2(n663), .B1(n664), .B2(n669), .ZN(n6070) );
  OAI22_X1 U946 ( .A1(n87), .A2(n663), .B1(n664), .B2(n670), .ZN(n6071) );
  OAI22_X1 U947 ( .A1(n89), .A2(n663), .B1(n664), .B2(n671), .ZN(n6072) );
  OAI22_X1 U948 ( .A1(n91), .A2(n663), .B1(n664), .B2(n672), .ZN(n6073) );
  OAI22_X1 U949 ( .A1(n93), .A2(n663), .B1(n664), .B2(n673), .ZN(n6074) );
  OAI22_X1 U950 ( .A1(n95), .A2(n663), .B1(n664), .B2(n674), .ZN(n6075) );
  OAI22_X1 U951 ( .A1(n97), .A2(n663), .B1(n664), .B2(n675), .ZN(n6076) );
  OAI22_X1 U952 ( .A1(n99), .A2(n663), .B1(n664), .B2(n676), .ZN(n6077) );
  OAI22_X1 U953 ( .A1(n101), .A2(n663), .B1(n664), .B2(n677), .ZN(n6078) );
  OAI22_X1 U954 ( .A1(n103), .A2(n663), .B1(n664), .B2(n678), .ZN(n6079) );
  OAI22_X1 U955 ( .A1(n105), .A2(n663), .B1(n664), .B2(n679), .ZN(n6080) );
  OAI22_X1 U956 ( .A1(n107), .A2(n663), .B1(n664), .B2(n680), .ZN(n6081) );
  OAI22_X1 U957 ( .A1(n109), .A2(n663), .B1(n664), .B2(n681), .ZN(n6082) );
  OAI22_X1 U958 ( .A1(n111), .A2(n663), .B1(n664), .B2(n682), .ZN(n6083) );
  OAI22_X1 U959 ( .A1(n113), .A2(n663), .B1(n664), .B2(n683), .ZN(n6084) );
  OAI22_X1 U960 ( .A1(n115), .A2(n663), .B1(n664), .B2(n684), .ZN(n6085) );
  OAI22_X1 U961 ( .A1(n117), .A2(n663), .B1(n664), .B2(n685), .ZN(n6086) );
  OAI22_X1 U962 ( .A1(n119), .A2(n663), .B1(n664), .B2(n686), .ZN(n6087) );
  OAI22_X1 U963 ( .A1(n121), .A2(n663), .B1(n664), .B2(n687), .ZN(n6088) );
  OAI22_X1 U964 ( .A1(n123), .A2(n663), .B1(n664), .B2(n688), .ZN(n6089) );
  OAI22_X1 U965 ( .A1(n125), .A2(n663), .B1(n664), .B2(n689), .ZN(n6090) );
  OAI22_X1 U966 ( .A1(n127), .A2(n663), .B1(n664), .B2(n690), .ZN(n6091) );
  OAI22_X1 U967 ( .A1(n129), .A2(n663), .B1(n664), .B2(n691), .ZN(n6092) );
  OAI22_X1 U968 ( .A1(n131), .A2(n663), .B1(n664), .B2(n692), .ZN(n6093) );
  OAI22_X1 U969 ( .A1(n133), .A2(n663), .B1(n664), .B2(n693), .ZN(n6094) );
  OAI22_X1 U970 ( .A1(n135), .A2(n663), .B1(n664), .B2(n694), .ZN(n6095) );
  OAI22_X1 U971 ( .A1(n137), .A2(n663), .B1(n664), .B2(n695), .ZN(n6096) );
  OAI22_X1 U972 ( .A1(n139), .A2(n663), .B1(n664), .B2(n696), .ZN(n6097) );
  OAI22_X1 U975 ( .A1(n75), .A2(n697), .B1(n698), .B2(n699), .ZN(n6098) );
  OAI22_X1 U976 ( .A1(n79), .A2(n697), .B1(n698), .B2(n700), .ZN(n6099) );
  OAI22_X1 U977 ( .A1(n81), .A2(n697), .B1(n698), .B2(n701), .ZN(n6100) );
  OAI22_X1 U978 ( .A1(n83), .A2(n697), .B1(n698), .B2(n702), .ZN(n6101) );
  OAI22_X1 U979 ( .A1(n85), .A2(n697), .B1(n698), .B2(n703), .ZN(n6102) );
  OAI22_X1 U980 ( .A1(n87), .A2(n697), .B1(n698), .B2(n704), .ZN(n6103) );
  OAI22_X1 U981 ( .A1(n89), .A2(n697), .B1(n698), .B2(n705), .ZN(n6104) );
  OAI22_X1 U982 ( .A1(n91), .A2(n697), .B1(n698), .B2(n706), .ZN(n6105) );
  OAI22_X1 U983 ( .A1(n93), .A2(n697), .B1(n698), .B2(n707), .ZN(n6106) );
  OAI22_X1 U984 ( .A1(n95), .A2(n697), .B1(n698), .B2(n708), .ZN(n6107) );
  OAI22_X1 U985 ( .A1(n97), .A2(n697), .B1(n698), .B2(n709), .ZN(n6108) );
  OAI22_X1 U986 ( .A1(n99), .A2(n697), .B1(n698), .B2(n710), .ZN(n6109) );
  OAI22_X1 U987 ( .A1(n101), .A2(n697), .B1(n698), .B2(n711), .ZN(n6110) );
  OAI22_X1 U988 ( .A1(n103), .A2(n697), .B1(n698), .B2(n712), .ZN(n6111) );
  OAI22_X1 U989 ( .A1(n105), .A2(n697), .B1(n698), .B2(n713), .ZN(n6112) );
  OAI22_X1 U990 ( .A1(n107), .A2(n697), .B1(n698), .B2(n714), .ZN(n6113) );
  OAI22_X1 U991 ( .A1(n109), .A2(n697), .B1(n698), .B2(n715), .ZN(n6114) );
  OAI22_X1 U992 ( .A1(n111), .A2(n697), .B1(n698), .B2(n716), .ZN(n6115) );
  OAI22_X1 U993 ( .A1(n113), .A2(n697), .B1(n698), .B2(n717), .ZN(n6116) );
  OAI22_X1 U994 ( .A1(n115), .A2(n697), .B1(n698), .B2(n718), .ZN(n6117) );
  OAI22_X1 U995 ( .A1(n117), .A2(n697), .B1(n698), .B2(n719), .ZN(n6118) );
  OAI22_X1 U996 ( .A1(n119), .A2(n697), .B1(n698), .B2(n720), .ZN(n6119) );
  OAI22_X1 U997 ( .A1(n121), .A2(n697), .B1(n698), .B2(n721), .ZN(n6120) );
  OAI22_X1 U998 ( .A1(n123), .A2(n697), .B1(n698), .B2(n722), .ZN(n6121) );
  OAI22_X1 U999 ( .A1(n125), .A2(n697), .B1(n698), .B2(n723), .ZN(n6122) );
  OAI22_X1 U1000 ( .A1(n127), .A2(n697), .B1(n698), .B2(n724), .ZN(n6123) );
  OAI22_X1 U1001 ( .A1(n129), .A2(n697), .B1(n698), .B2(n725), .ZN(n6124) );
  OAI22_X1 U1002 ( .A1(n131), .A2(n697), .B1(n698), .B2(n726), .ZN(n6125) );
  OAI22_X1 U1003 ( .A1(n133), .A2(n697), .B1(n698), .B2(n727), .ZN(n6126) );
  OAI22_X1 U1004 ( .A1(n135), .A2(n697), .B1(n698), .B2(n728), .ZN(n6127) );
  OAI22_X1 U1005 ( .A1(n137), .A2(n697), .B1(n698), .B2(n729), .ZN(n6128) );
  OAI22_X1 U1006 ( .A1(n139), .A2(n697), .B1(n698), .B2(n730), .ZN(n6129) );
  INV_X1 U1010 ( .A(n732), .ZN(n6130) );
  AOI22_X1 U1011 ( .A1(Set_target[30]), .A2(n733), .B1(n734), .B2(
        \pc_target[11][30] ), .ZN(n732) );
  INV_X1 U1012 ( .A(n735), .ZN(n6131) );
  AOI22_X1 U1013 ( .A1(Set_target[28]), .A2(n733), .B1(n734), .B2(
        \pc_target[11][28] ), .ZN(n735) );
  INV_X1 U1014 ( .A(n736), .ZN(n6132) );
  AOI22_X1 U1015 ( .A1(Set_target[26]), .A2(n733), .B1(n734), .B2(
        \pc_target[11][26] ), .ZN(n736) );
  INV_X1 U1016 ( .A(n737), .ZN(n6133) );
  AOI22_X1 U1017 ( .A1(Set_target[24]), .A2(n733), .B1(n734), .B2(
        \pc_target[11][24] ), .ZN(n737) );
  INV_X1 U1018 ( .A(n738), .ZN(n6134) );
  AOI22_X1 U1019 ( .A1(Set_target[22]), .A2(n733), .B1(n734), .B2(
        \pc_target[11][22] ), .ZN(n738) );
  INV_X1 U1020 ( .A(n739), .ZN(n6135) );
  AOI22_X1 U1021 ( .A1(Set_target[20]), .A2(n733), .B1(n734), .B2(
        \pc_target[11][20] ), .ZN(n739) );
  INV_X1 U1022 ( .A(n740), .ZN(n6136) );
  AOI22_X1 U1023 ( .A1(Set_target[18]), .A2(n733), .B1(n734), .B2(
        \pc_target[11][18] ), .ZN(n740) );
  INV_X1 U1024 ( .A(n741), .ZN(n6137) );
  AOI22_X1 U1025 ( .A1(Set_target[16]), .A2(n733), .B1(n734), .B2(
        \pc_target[11][16] ), .ZN(n741) );
  INV_X1 U1026 ( .A(n742), .ZN(n6138) );
  AOI22_X1 U1027 ( .A1(Set_target[14]), .A2(n733), .B1(n734), .B2(
        \pc_target[11][14] ), .ZN(n742) );
  INV_X1 U1028 ( .A(n743), .ZN(n6139) );
  AOI22_X1 U1029 ( .A1(Set_target[12]), .A2(n733), .B1(n734), .B2(
        \pc_target[11][12] ), .ZN(n743) );
  INV_X1 U1030 ( .A(n744), .ZN(n6140) );
  AOI22_X1 U1031 ( .A1(Set_target[10]), .A2(n733), .B1(n734), .B2(
        \pc_target[11][10] ), .ZN(n744) );
  INV_X1 U1032 ( .A(n745), .ZN(n6141) );
  AOI22_X1 U1033 ( .A1(Set_target[8]), .A2(n733), .B1(n734), .B2(
        \pc_target[11][8] ), .ZN(n745) );
  INV_X1 U1034 ( .A(n746), .ZN(n6142) );
  AOI22_X1 U1035 ( .A1(Set_target[6]), .A2(n733), .B1(n734), .B2(
        \pc_target[11][6] ), .ZN(n746) );
  INV_X1 U1036 ( .A(n747), .ZN(n6143) );
  AOI22_X1 U1037 ( .A1(Set_target[4]), .A2(n733), .B1(n734), .B2(
        \pc_target[11][4] ), .ZN(n747) );
  INV_X1 U1038 ( .A(n748), .ZN(n6144) );
  AOI22_X1 U1039 ( .A1(Set_target[2]), .A2(n733), .B1(n734), .B2(
        \pc_target[11][2] ), .ZN(n748) );
  INV_X1 U1040 ( .A(n749), .ZN(n6145) );
  AOI22_X1 U1041 ( .A1(Set_target[0]), .A2(n733), .B1(n734), .B2(
        \pc_target[11][0] ), .ZN(n749) );
  INV_X1 U1042 ( .A(n750), .ZN(n6146) );
  AOI22_X1 U1043 ( .A1(Set_target[1]), .A2(n733), .B1(n734), .B2(
        \pc_target[11][1] ), .ZN(n750) );
  INV_X1 U1044 ( .A(n751), .ZN(n6147) );
  AOI22_X1 U1045 ( .A1(Set_target[3]), .A2(n733), .B1(n734), .B2(
        \pc_target[11][3] ), .ZN(n751) );
  INV_X1 U1046 ( .A(n752), .ZN(n6148) );
  AOI22_X1 U1047 ( .A1(Set_target[5]), .A2(n733), .B1(n734), .B2(
        \pc_target[11][5] ), .ZN(n752) );
  INV_X1 U1048 ( .A(n753), .ZN(n6149) );
  AOI22_X1 U1049 ( .A1(Set_target[7]), .A2(n733), .B1(n734), .B2(
        \pc_target[11][7] ), .ZN(n753) );
  INV_X1 U1050 ( .A(n754), .ZN(n6150) );
  AOI22_X1 U1051 ( .A1(Set_target[9]), .A2(n733), .B1(n734), .B2(
        \pc_target[11][9] ), .ZN(n754) );
  INV_X1 U1052 ( .A(n755), .ZN(n6151) );
  AOI22_X1 U1053 ( .A1(Set_target[11]), .A2(n733), .B1(n734), .B2(
        \pc_target[11][11] ), .ZN(n755) );
  INV_X1 U1054 ( .A(n756), .ZN(n6152) );
  AOI22_X1 U1055 ( .A1(Set_target[13]), .A2(n733), .B1(n734), .B2(
        \pc_target[11][13] ), .ZN(n756) );
  INV_X1 U1056 ( .A(n757), .ZN(n6153) );
  AOI22_X1 U1057 ( .A1(Set_target[15]), .A2(n733), .B1(n734), .B2(
        \pc_target[11][15] ), .ZN(n757) );
  INV_X1 U1058 ( .A(n758), .ZN(n6154) );
  AOI22_X1 U1059 ( .A1(Set_target[17]), .A2(n733), .B1(n734), .B2(
        \pc_target[11][17] ), .ZN(n758) );
  INV_X1 U1060 ( .A(n759), .ZN(n6155) );
  AOI22_X1 U1061 ( .A1(Set_target[19]), .A2(n733), .B1(n734), .B2(
        \pc_target[11][19] ), .ZN(n759) );
  INV_X1 U1062 ( .A(n760), .ZN(n6156) );
  AOI22_X1 U1063 ( .A1(Set_target[21]), .A2(n733), .B1(n734), .B2(
        \pc_target[11][21] ), .ZN(n760) );
  INV_X1 U1064 ( .A(n761), .ZN(n6157) );
  AOI22_X1 U1065 ( .A1(Set_target[23]), .A2(n733), .B1(n734), .B2(
        \pc_target[11][23] ), .ZN(n761) );
  INV_X1 U1066 ( .A(n762), .ZN(n6158) );
  AOI22_X1 U1067 ( .A1(Set_target[25]), .A2(n733), .B1(n734), .B2(
        \pc_target[11][25] ), .ZN(n762) );
  INV_X1 U1068 ( .A(n763), .ZN(n6159) );
  AOI22_X1 U1069 ( .A1(Set_target[27]), .A2(n733), .B1(n734), .B2(
        \pc_target[11][27] ), .ZN(n763) );
  INV_X1 U1070 ( .A(n764), .ZN(n6160) );
  AOI22_X1 U1071 ( .A1(Set_target[29]), .A2(n733), .B1(n734), .B2(
        \pc_target[11][29] ), .ZN(n764) );
  INV_X1 U1072 ( .A(n765), .ZN(n6161) );
  AOI22_X1 U1073 ( .A1(Set_target[31]), .A2(n733), .B1(n734), .B2(
        \pc_target[11][31] ), .ZN(n765) );
  INV_X1 U1076 ( .A(n767), .ZN(n6162) );
  AOI22_X1 U1077 ( .A1(Set_target[30]), .A2(n3446), .B1(n769), .B2(
        \pc_target[10][30] ), .ZN(n767) );
  INV_X1 U1078 ( .A(n770), .ZN(n6163) );
  AOI22_X1 U1079 ( .A1(Set_target[28]), .A2(n3446), .B1(n769), .B2(
        \pc_target[10][28] ), .ZN(n770) );
  INV_X1 U1080 ( .A(n771), .ZN(n6164) );
  AOI22_X1 U1081 ( .A1(Set_target[26]), .A2(n3446), .B1(n769), .B2(
        \pc_target[10][26] ), .ZN(n771) );
  INV_X1 U1082 ( .A(n772), .ZN(n6165) );
  AOI22_X1 U1083 ( .A1(Set_target[24]), .A2(n3446), .B1(n769), .B2(
        \pc_target[10][24] ), .ZN(n772) );
  INV_X1 U1084 ( .A(n773), .ZN(n6166) );
  AOI22_X1 U1085 ( .A1(Set_target[22]), .A2(n3446), .B1(n769), .B2(
        \pc_target[10][22] ), .ZN(n773) );
  INV_X1 U1086 ( .A(n774), .ZN(n6167) );
  AOI22_X1 U1087 ( .A1(Set_target[20]), .A2(n3446), .B1(n769), .B2(
        \pc_target[10][20] ), .ZN(n774) );
  INV_X1 U1088 ( .A(n775), .ZN(n6168) );
  AOI22_X1 U1089 ( .A1(Set_target[18]), .A2(n3446), .B1(n769), .B2(
        \pc_target[10][18] ), .ZN(n775) );
  INV_X1 U1090 ( .A(n776), .ZN(n6169) );
  AOI22_X1 U1091 ( .A1(Set_target[16]), .A2(n3446), .B1(n769), .B2(
        \pc_target[10][16] ), .ZN(n776) );
  INV_X1 U1092 ( .A(n777), .ZN(n6170) );
  AOI22_X1 U1093 ( .A1(Set_target[14]), .A2(n3446), .B1(n769), .B2(
        \pc_target[10][14] ), .ZN(n777) );
  INV_X1 U1094 ( .A(n778), .ZN(n6171) );
  AOI22_X1 U1095 ( .A1(Set_target[12]), .A2(n3446), .B1(n769), .B2(
        \pc_target[10][12] ), .ZN(n778) );
  INV_X1 U1096 ( .A(n779), .ZN(n6172) );
  AOI22_X1 U1097 ( .A1(Set_target[10]), .A2(n3446), .B1(n769), .B2(
        \pc_target[10][10] ), .ZN(n779) );
  INV_X1 U1098 ( .A(n780), .ZN(n6173) );
  AOI22_X1 U1099 ( .A1(Set_target[8]), .A2(n3446), .B1(n769), .B2(
        \pc_target[10][8] ), .ZN(n780) );
  INV_X1 U1100 ( .A(n781), .ZN(n6174) );
  AOI22_X1 U1101 ( .A1(Set_target[6]), .A2(n3446), .B1(n769), .B2(
        \pc_target[10][6] ), .ZN(n781) );
  INV_X1 U1102 ( .A(n782), .ZN(n6175) );
  AOI22_X1 U1103 ( .A1(Set_target[4]), .A2(n3446), .B1(n769), .B2(
        \pc_target[10][4] ), .ZN(n782) );
  INV_X1 U1104 ( .A(n783), .ZN(n6176) );
  AOI22_X1 U1105 ( .A1(Set_target[2]), .A2(n3446), .B1(n769), .B2(
        \pc_target[10][2] ), .ZN(n783) );
  INV_X1 U1106 ( .A(n784), .ZN(n6177) );
  AOI22_X1 U1107 ( .A1(Set_target[0]), .A2(n3446), .B1(n769), .B2(
        \pc_target[10][0] ), .ZN(n784) );
  INV_X1 U1108 ( .A(n785), .ZN(n6178) );
  AOI22_X1 U1109 ( .A1(Set_target[1]), .A2(n3446), .B1(n769), .B2(
        \pc_target[10][1] ), .ZN(n785) );
  INV_X1 U1110 ( .A(n786), .ZN(n6179) );
  AOI22_X1 U1111 ( .A1(Set_target[3]), .A2(n3446), .B1(n769), .B2(
        \pc_target[10][3] ), .ZN(n786) );
  INV_X1 U1112 ( .A(n787), .ZN(n6180) );
  AOI22_X1 U1113 ( .A1(Set_target[5]), .A2(n3446), .B1(n769), .B2(
        \pc_target[10][5] ), .ZN(n787) );
  INV_X1 U1114 ( .A(n788), .ZN(n6181) );
  AOI22_X1 U1115 ( .A1(Set_target[7]), .A2(n3446), .B1(n769), .B2(
        \pc_target[10][7] ), .ZN(n788) );
  INV_X1 U1116 ( .A(n789), .ZN(n6182) );
  AOI22_X1 U1117 ( .A1(Set_target[9]), .A2(n3446), .B1(n769), .B2(
        \pc_target[10][9] ), .ZN(n789) );
  INV_X1 U1118 ( .A(n790), .ZN(n6183) );
  AOI22_X1 U1119 ( .A1(Set_target[11]), .A2(n3446), .B1(n769), .B2(
        \pc_target[10][11] ), .ZN(n790) );
  INV_X1 U1120 ( .A(n791), .ZN(n6184) );
  AOI22_X1 U1121 ( .A1(Set_target[13]), .A2(n3446), .B1(n769), .B2(
        \pc_target[10][13] ), .ZN(n791) );
  INV_X1 U1122 ( .A(n792), .ZN(n6185) );
  AOI22_X1 U1123 ( .A1(Set_target[15]), .A2(n3446), .B1(n769), .B2(
        \pc_target[10][15] ), .ZN(n792) );
  INV_X1 U1124 ( .A(n793), .ZN(n6186) );
  AOI22_X1 U1125 ( .A1(Set_target[17]), .A2(n3446), .B1(n769), .B2(
        \pc_target[10][17] ), .ZN(n793) );
  INV_X1 U1126 ( .A(n794), .ZN(n6187) );
  AOI22_X1 U1127 ( .A1(Set_target[19]), .A2(n3446), .B1(n769), .B2(
        \pc_target[10][19] ), .ZN(n794) );
  INV_X1 U1128 ( .A(n795), .ZN(n6188) );
  AOI22_X1 U1129 ( .A1(Set_target[21]), .A2(n3446), .B1(n769), .B2(
        \pc_target[10][21] ), .ZN(n795) );
  INV_X1 U1130 ( .A(n796), .ZN(n6189) );
  AOI22_X1 U1131 ( .A1(Set_target[23]), .A2(n3446), .B1(n769), .B2(
        \pc_target[10][23] ), .ZN(n796) );
  INV_X1 U1132 ( .A(n797), .ZN(n6190) );
  AOI22_X1 U1133 ( .A1(Set_target[25]), .A2(n3446), .B1(n769), .B2(
        \pc_target[10][25] ), .ZN(n797) );
  INV_X1 U1134 ( .A(n798), .ZN(n6191) );
  AOI22_X1 U1135 ( .A1(Set_target[27]), .A2(n3446), .B1(n769), .B2(
        \pc_target[10][27] ), .ZN(n798) );
  INV_X1 U1136 ( .A(n799), .ZN(n6192) );
  AOI22_X1 U1137 ( .A1(Set_target[29]), .A2(n3446), .B1(n769), .B2(
        \pc_target[10][29] ), .ZN(n799) );
  INV_X1 U1138 ( .A(n800), .ZN(n6193) );
  AOI22_X1 U1139 ( .A1(Set_target[31]), .A2(n3446), .B1(n769), .B2(
        \pc_target[10][31] ), .ZN(n800) );
  OAI22_X1 U1142 ( .A1(n75), .A2(n801), .B1(n3442), .B2(n803), .ZN(n6194) );
  OAI22_X1 U1143 ( .A1(n79), .A2(n801), .B1(n3442), .B2(n804), .ZN(n6195) );
  OAI22_X1 U1144 ( .A1(n81), .A2(n801), .B1(n3442), .B2(n805), .ZN(n6196) );
  OAI22_X1 U1145 ( .A1(n83), .A2(n801), .B1(n3442), .B2(n806), .ZN(n6197) );
  OAI22_X1 U1146 ( .A1(n85), .A2(n801), .B1(n3442), .B2(n807), .ZN(n6198) );
  OAI22_X1 U1147 ( .A1(n87), .A2(n801), .B1(n3442), .B2(n808), .ZN(n6199) );
  OAI22_X1 U1148 ( .A1(n89), .A2(n801), .B1(n3442), .B2(n809), .ZN(n6200) );
  OAI22_X1 U1149 ( .A1(n91), .A2(n801), .B1(n3442), .B2(n810), .ZN(n6201) );
  OAI22_X1 U1150 ( .A1(n93), .A2(n801), .B1(n3442), .B2(n811), .ZN(n6202) );
  OAI22_X1 U1151 ( .A1(n95), .A2(n801), .B1(n3442), .B2(n812), .ZN(n6203) );
  OAI22_X1 U1152 ( .A1(n97), .A2(n801), .B1(n3442), .B2(n813), .ZN(n6204) );
  OAI22_X1 U1153 ( .A1(n99), .A2(n801), .B1(n3442), .B2(n814), .ZN(n6205) );
  OAI22_X1 U1154 ( .A1(n101), .A2(n801), .B1(n3442), .B2(n815), .ZN(n6206) );
  OAI22_X1 U1155 ( .A1(n103), .A2(n801), .B1(n3442), .B2(n816), .ZN(n6207) );
  OAI22_X1 U1156 ( .A1(n105), .A2(n801), .B1(n3442), .B2(n817), .ZN(n6208) );
  OAI22_X1 U1157 ( .A1(n107), .A2(n801), .B1(n3442), .B2(n818), .ZN(n6209) );
  OAI22_X1 U1158 ( .A1(n109), .A2(n801), .B1(n3442), .B2(n819), .ZN(n6210) );
  OAI22_X1 U1159 ( .A1(n111), .A2(n801), .B1(n3442), .B2(n820), .ZN(n6211) );
  OAI22_X1 U1160 ( .A1(n113), .A2(n801), .B1(n3442), .B2(n821), .ZN(n6212) );
  OAI22_X1 U1161 ( .A1(n115), .A2(n801), .B1(n3442), .B2(n822), .ZN(n6213) );
  OAI22_X1 U1162 ( .A1(n117), .A2(n801), .B1(n3442), .B2(n823), .ZN(n6214) );
  OAI22_X1 U1163 ( .A1(n119), .A2(n801), .B1(n3442), .B2(n824), .ZN(n6215) );
  OAI22_X1 U1164 ( .A1(n121), .A2(n801), .B1(n3442), .B2(n825), .ZN(n6216) );
  OAI22_X1 U1165 ( .A1(n123), .A2(n801), .B1(n3442), .B2(n826), .ZN(n6217) );
  OAI22_X1 U1166 ( .A1(n125), .A2(n801), .B1(n3442), .B2(n827), .ZN(n6218) );
  OAI22_X1 U1167 ( .A1(n127), .A2(n801), .B1(n3442), .B2(n828), .ZN(n6219) );
  OAI22_X1 U1168 ( .A1(n129), .A2(n801), .B1(n3442), .B2(n829), .ZN(n6220) );
  OAI22_X1 U1169 ( .A1(n131), .A2(n801), .B1(n3442), .B2(n830), .ZN(n6221) );
  OAI22_X1 U1170 ( .A1(n133), .A2(n801), .B1(n3442), .B2(n831), .ZN(n6222) );
  OAI22_X1 U1171 ( .A1(n135), .A2(n801), .B1(n3442), .B2(n832), .ZN(n6223) );
  OAI22_X1 U1172 ( .A1(n137), .A2(n801), .B1(n3442), .B2(n833), .ZN(n6224) );
  OAI22_X1 U1173 ( .A1(n139), .A2(n801), .B1(n3442), .B2(n834), .ZN(n6225) );
  OAI22_X1 U1176 ( .A1(n75), .A2(n835), .B1(n836), .B2(n837), .ZN(n6226) );
  OAI22_X1 U1177 ( .A1(n79), .A2(n835), .B1(n836), .B2(n838), .ZN(n6227) );
  OAI22_X1 U1178 ( .A1(n81), .A2(n835), .B1(n836), .B2(n839), .ZN(n6228) );
  OAI22_X1 U1179 ( .A1(n83), .A2(n835), .B1(n836), .B2(n840), .ZN(n6229) );
  OAI22_X1 U1180 ( .A1(n85), .A2(n835), .B1(n836), .B2(n841), .ZN(n6230) );
  OAI22_X1 U1181 ( .A1(n87), .A2(n835), .B1(n836), .B2(n842), .ZN(n6231) );
  OAI22_X1 U1182 ( .A1(n89), .A2(n835), .B1(n836), .B2(n843), .ZN(n6232) );
  OAI22_X1 U1183 ( .A1(n91), .A2(n835), .B1(n836), .B2(n844), .ZN(n6233) );
  OAI22_X1 U1184 ( .A1(n93), .A2(n835), .B1(n836), .B2(n845), .ZN(n6234) );
  OAI22_X1 U1185 ( .A1(n95), .A2(n835), .B1(n836), .B2(n846), .ZN(n6235) );
  OAI22_X1 U1186 ( .A1(n97), .A2(n835), .B1(n836), .B2(n847), .ZN(n6236) );
  OAI22_X1 U1187 ( .A1(n99), .A2(n835), .B1(n836), .B2(n848), .ZN(n6237) );
  OAI22_X1 U1188 ( .A1(n101), .A2(n835), .B1(n836), .B2(n849), .ZN(n6238) );
  OAI22_X1 U1189 ( .A1(n103), .A2(n835), .B1(n836), .B2(n850), .ZN(n6239) );
  OAI22_X1 U1190 ( .A1(n105), .A2(n835), .B1(n836), .B2(n851), .ZN(n6240) );
  OAI22_X1 U1191 ( .A1(n107), .A2(n835), .B1(n836), .B2(n852), .ZN(n6241) );
  OAI22_X1 U1192 ( .A1(n109), .A2(n835), .B1(n836), .B2(n853), .ZN(n6242) );
  OAI22_X1 U1193 ( .A1(n111), .A2(n835), .B1(n836), .B2(n854), .ZN(n6243) );
  OAI22_X1 U1194 ( .A1(n113), .A2(n835), .B1(n836), .B2(n855), .ZN(n6244) );
  OAI22_X1 U1195 ( .A1(n115), .A2(n835), .B1(n836), .B2(n856), .ZN(n6245) );
  OAI22_X1 U1196 ( .A1(n117), .A2(n835), .B1(n836), .B2(n857), .ZN(n6246) );
  OAI22_X1 U1197 ( .A1(n119), .A2(n835), .B1(n836), .B2(n858), .ZN(n6247) );
  OAI22_X1 U1198 ( .A1(n121), .A2(n835), .B1(n836), .B2(n859), .ZN(n6248) );
  OAI22_X1 U1199 ( .A1(n123), .A2(n835), .B1(n836), .B2(n860), .ZN(n6249) );
  OAI22_X1 U1200 ( .A1(n125), .A2(n835), .B1(n836), .B2(n861), .ZN(n6250) );
  OAI22_X1 U1201 ( .A1(n127), .A2(n835), .B1(n836), .B2(n862), .ZN(n6251) );
  OAI22_X1 U1202 ( .A1(n129), .A2(n835), .B1(n836), .B2(n863), .ZN(n6252) );
  OAI22_X1 U1203 ( .A1(n131), .A2(n835), .B1(n836), .B2(n864), .ZN(n6253) );
  OAI22_X1 U1204 ( .A1(n133), .A2(n835), .B1(n836), .B2(n865), .ZN(n6254) );
  OAI22_X1 U1205 ( .A1(n135), .A2(n835), .B1(n836), .B2(n866), .ZN(n6255) );
  OAI22_X1 U1206 ( .A1(n137), .A2(n835), .B1(n836), .B2(n867), .ZN(n6256) );
  OAI22_X1 U1207 ( .A1(n139), .A2(n835), .B1(n836), .B2(n868), .ZN(n6257) );
  INV_X1 U1211 ( .A(n869), .ZN(n6258) );
  AOI22_X1 U1212 ( .A1(Set_target[30]), .A2(n870), .B1(n1656), .B2(
        \pc_target[7][30] ), .ZN(n869) );
  INV_X1 U1213 ( .A(n872), .ZN(n6259) );
  AOI22_X1 U1214 ( .A1(Set_target[28]), .A2(n870), .B1(n1656), .B2(
        \pc_target[7][28] ), .ZN(n872) );
  INV_X1 U1215 ( .A(n873), .ZN(n6260) );
  AOI22_X1 U1216 ( .A1(Set_target[26]), .A2(n870), .B1(n1611), .B2(
        \pc_target[7][26] ), .ZN(n873) );
  INV_X1 U1217 ( .A(n874), .ZN(n6261) );
  AOI22_X1 U1218 ( .A1(Set_target[24]), .A2(n870), .B1(n1656), .B2(
        \pc_target[7][24] ), .ZN(n874) );
  INV_X1 U1219 ( .A(n875), .ZN(n6262) );
  AOI22_X1 U1220 ( .A1(Set_target[22]), .A2(n870), .B1(n1656), .B2(
        \pc_target[7][22] ), .ZN(n875) );
  INV_X1 U1221 ( .A(n876), .ZN(n6263) );
  AOI22_X1 U1222 ( .A1(Set_target[20]), .A2(n870), .B1(n1656), .B2(
        \pc_target[7][20] ), .ZN(n876) );
  INV_X1 U1223 ( .A(n877), .ZN(n6264) );
  AOI22_X1 U1224 ( .A1(Set_target[18]), .A2(n870), .B1(n1656), .B2(
        \pc_target[7][18] ), .ZN(n877) );
  INV_X1 U1225 ( .A(n878), .ZN(n6265) );
  AOI22_X1 U1226 ( .A1(Set_target[16]), .A2(n870), .B1(n1656), .B2(
        \pc_target[7][16] ), .ZN(n878) );
  INV_X1 U1227 ( .A(n879), .ZN(n6266) );
  AOI22_X1 U1228 ( .A1(Set_target[14]), .A2(n870), .B1(n1611), .B2(
        \pc_target[7][14] ), .ZN(n879) );
  INV_X1 U1229 ( .A(n880), .ZN(n6267) );
  AOI22_X1 U1230 ( .A1(Set_target[12]), .A2(n870), .B1(n1656), .B2(
        \pc_target[7][12] ), .ZN(n880) );
  INV_X1 U1231 ( .A(n881), .ZN(n6268) );
  AOI22_X1 U1232 ( .A1(Set_target[10]), .A2(n870), .B1(n1656), .B2(
        \pc_target[7][10] ), .ZN(n881) );
  INV_X1 U1233 ( .A(n882), .ZN(n6269) );
  AOI22_X1 U1234 ( .A1(Set_target[8]), .A2(n870), .B1(n1656), .B2(
        \pc_target[7][8] ), .ZN(n882) );
  INV_X1 U1235 ( .A(n883), .ZN(n6270) );
  AOI22_X1 U1236 ( .A1(Set_target[6]), .A2(n870), .B1(n1656), .B2(
        \pc_target[7][6] ), .ZN(n883) );
  INV_X1 U1237 ( .A(n884), .ZN(n6271) );
  AOI22_X1 U1238 ( .A1(Set_target[4]), .A2(n870), .B1(n1656), .B2(
        \pc_target[7][4] ), .ZN(n884) );
  INV_X1 U1239 ( .A(n885), .ZN(n6272) );
  AOI22_X1 U1240 ( .A1(Set_target[2]), .A2(n870), .B1(n1656), .B2(
        \pc_target[7][2] ), .ZN(n885) );
  INV_X1 U1241 ( .A(n886), .ZN(n6273) );
  AOI22_X1 U1242 ( .A1(Set_target[0]), .A2(n870), .B1(n1656), .B2(
        \pc_target[7][0] ), .ZN(n886) );
  INV_X1 U1243 ( .A(n887), .ZN(n6274) );
  AOI22_X1 U1244 ( .A1(Set_target[1]), .A2(n870), .B1(n1656), .B2(
        \pc_target[7][1] ), .ZN(n887) );
  INV_X1 U1245 ( .A(n888), .ZN(n6275) );
  AOI22_X1 U1246 ( .A1(Set_target[3]), .A2(n870), .B1(n1656), .B2(
        \pc_target[7][3] ), .ZN(n888) );
  INV_X1 U1247 ( .A(n889), .ZN(n6276) );
  AOI22_X1 U1248 ( .A1(Set_target[5]), .A2(n870), .B1(n1656), .B2(
        \pc_target[7][5] ), .ZN(n889) );
  INV_X1 U1249 ( .A(n890), .ZN(n6277) );
  AOI22_X1 U1250 ( .A1(Set_target[7]), .A2(n870), .B1(n1656), .B2(
        \pc_target[7][7] ), .ZN(n890) );
  INV_X1 U1251 ( .A(n891), .ZN(n6278) );
  AOI22_X1 U1252 ( .A1(Set_target[9]), .A2(n870), .B1(n1656), .B2(
        \pc_target[7][9] ), .ZN(n891) );
  INV_X1 U1253 ( .A(n892), .ZN(n6279) );
  AOI22_X1 U1254 ( .A1(Set_target[11]), .A2(n870), .B1(n1611), .B2(
        \pc_target[7][11] ), .ZN(n892) );
  INV_X1 U1255 ( .A(n893), .ZN(n6280) );
  AOI22_X1 U1256 ( .A1(Set_target[13]), .A2(n870), .B1(n1656), .B2(
        \pc_target[7][13] ), .ZN(n893) );
  INV_X1 U1257 ( .A(n894), .ZN(n6281) );
  AOI22_X1 U1258 ( .A1(Set_target[15]), .A2(n870), .B1(n1656), .B2(
        \pc_target[7][15] ), .ZN(n894) );
  INV_X1 U1259 ( .A(n895), .ZN(n6282) );
  AOI22_X1 U1260 ( .A1(Set_target[17]), .A2(n870), .B1(n1656), .B2(
        \pc_target[7][17] ), .ZN(n895) );
  INV_X1 U1261 ( .A(n896), .ZN(n6283) );
  AOI22_X1 U1262 ( .A1(Set_target[19]), .A2(n870), .B1(n1611), .B2(
        \pc_target[7][19] ), .ZN(n896) );
  INV_X1 U1263 ( .A(n897), .ZN(n6284) );
  AOI22_X1 U1264 ( .A1(Set_target[21]), .A2(n870), .B1(n1656), .B2(
        \pc_target[7][21] ), .ZN(n897) );
  INV_X1 U1265 ( .A(n898), .ZN(n6285) );
  AOI22_X1 U1266 ( .A1(Set_target[23]), .A2(n870), .B1(n1611), .B2(
        \pc_target[7][23] ), .ZN(n898) );
  INV_X1 U1267 ( .A(n899), .ZN(n6286) );
  AOI22_X1 U1268 ( .A1(Set_target[25]), .A2(n870), .B1(n1656), .B2(
        \pc_target[7][25] ), .ZN(n899) );
  INV_X1 U1269 ( .A(n900), .ZN(n6287) );
  AOI22_X1 U1270 ( .A1(Set_target[27]), .A2(n870), .B1(n1656), .B2(
        \pc_target[7][27] ), .ZN(n900) );
  INV_X1 U1271 ( .A(n901), .ZN(n6288) );
  AOI22_X1 U1272 ( .A1(Set_target[29]), .A2(n870), .B1(n1656), .B2(
        \pc_target[7][29] ), .ZN(n901) );
  INV_X1 U1273 ( .A(n902), .ZN(n6289) );
  AOI22_X1 U1274 ( .A1(Set_target[31]), .A2(n870), .B1(n1611), .B2(
        \pc_target[7][31] ), .ZN(n902) );
  INV_X1 U1277 ( .A(n904), .ZN(n6290) );
  AOI22_X1 U1278 ( .A1(Set_target[30]), .A2(n905), .B1(n906), .B2(
        \pc_target[6][30] ), .ZN(n904) );
  INV_X1 U1279 ( .A(n907), .ZN(n6291) );
  AOI22_X1 U1280 ( .A1(Set_target[28]), .A2(n905), .B1(n906), .B2(
        \pc_target[6][28] ), .ZN(n907) );
  INV_X1 U1281 ( .A(n908), .ZN(n6292) );
  AOI22_X1 U1282 ( .A1(Set_target[26]), .A2(n905), .B1(n906), .B2(
        \pc_target[6][26] ), .ZN(n908) );
  INV_X1 U1283 ( .A(n909), .ZN(n6293) );
  AOI22_X1 U1284 ( .A1(Set_target[24]), .A2(n905), .B1(n906), .B2(
        \pc_target[6][24] ), .ZN(n909) );
  INV_X1 U1285 ( .A(n910), .ZN(n6294) );
  AOI22_X1 U1286 ( .A1(Set_target[22]), .A2(n905), .B1(n906), .B2(
        \pc_target[6][22] ), .ZN(n910) );
  INV_X1 U1287 ( .A(n911), .ZN(n6295) );
  AOI22_X1 U1288 ( .A1(Set_target[20]), .A2(n905), .B1(n906), .B2(
        \pc_target[6][20] ), .ZN(n911) );
  INV_X1 U1289 ( .A(n912), .ZN(n6296) );
  AOI22_X1 U1290 ( .A1(Set_target[18]), .A2(n905), .B1(n906), .B2(
        \pc_target[6][18] ), .ZN(n912) );
  INV_X1 U1291 ( .A(n913), .ZN(n6297) );
  AOI22_X1 U1292 ( .A1(Set_target[16]), .A2(n905), .B1(n906), .B2(
        \pc_target[6][16] ), .ZN(n913) );
  INV_X1 U1293 ( .A(n914), .ZN(n6298) );
  AOI22_X1 U1294 ( .A1(Set_target[14]), .A2(n905), .B1(n906), .B2(
        \pc_target[6][14] ), .ZN(n914) );
  INV_X1 U1295 ( .A(n915), .ZN(n6299) );
  AOI22_X1 U1296 ( .A1(Set_target[12]), .A2(n905), .B1(n906), .B2(
        \pc_target[6][12] ), .ZN(n915) );
  INV_X1 U1297 ( .A(n916), .ZN(n6300) );
  AOI22_X1 U1298 ( .A1(Set_target[10]), .A2(n905), .B1(n906), .B2(
        \pc_target[6][10] ), .ZN(n916) );
  INV_X1 U1299 ( .A(n917), .ZN(n6301) );
  AOI22_X1 U1300 ( .A1(Set_target[8]), .A2(n905), .B1(n906), .B2(
        \pc_target[6][8] ), .ZN(n917) );
  INV_X1 U1301 ( .A(n918), .ZN(n6302) );
  AOI22_X1 U1302 ( .A1(Set_target[6]), .A2(n905), .B1(n906), .B2(
        \pc_target[6][6] ), .ZN(n918) );
  INV_X1 U1303 ( .A(n919), .ZN(n6303) );
  AOI22_X1 U1304 ( .A1(Set_target[4]), .A2(n905), .B1(n906), .B2(
        \pc_target[6][4] ), .ZN(n919) );
  INV_X1 U1305 ( .A(n920), .ZN(n6304) );
  AOI22_X1 U1306 ( .A1(Set_target[2]), .A2(n905), .B1(n906), .B2(
        \pc_target[6][2] ), .ZN(n920) );
  INV_X1 U1307 ( .A(n921), .ZN(n6305) );
  AOI22_X1 U1308 ( .A1(Set_target[0]), .A2(n905), .B1(n906), .B2(
        \pc_target[6][0] ), .ZN(n921) );
  INV_X1 U1309 ( .A(n922), .ZN(n6306) );
  AOI22_X1 U1310 ( .A1(Set_target[1]), .A2(n905), .B1(n906), .B2(
        \pc_target[6][1] ), .ZN(n922) );
  INV_X1 U1311 ( .A(n923), .ZN(n6307) );
  AOI22_X1 U1312 ( .A1(Set_target[3]), .A2(n905), .B1(n906), .B2(
        \pc_target[6][3] ), .ZN(n923) );
  INV_X1 U1313 ( .A(n924), .ZN(n6308) );
  AOI22_X1 U1314 ( .A1(Set_target[5]), .A2(n905), .B1(n906), .B2(
        \pc_target[6][5] ), .ZN(n924) );
  INV_X1 U1315 ( .A(n925), .ZN(n6309) );
  AOI22_X1 U1316 ( .A1(Set_target[7]), .A2(n905), .B1(n906), .B2(
        \pc_target[6][7] ), .ZN(n925) );
  INV_X1 U1317 ( .A(n926), .ZN(n6310) );
  AOI22_X1 U1318 ( .A1(Set_target[9]), .A2(n905), .B1(n906), .B2(
        \pc_target[6][9] ), .ZN(n926) );
  INV_X1 U1319 ( .A(n927), .ZN(n6311) );
  AOI22_X1 U1320 ( .A1(Set_target[11]), .A2(n905), .B1(n906), .B2(
        \pc_target[6][11] ), .ZN(n927) );
  INV_X1 U1321 ( .A(n928), .ZN(n6312) );
  AOI22_X1 U1322 ( .A1(Set_target[13]), .A2(n905), .B1(n906), .B2(
        \pc_target[6][13] ), .ZN(n928) );
  INV_X1 U1323 ( .A(n929), .ZN(n6313) );
  AOI22_X1 U1324 ( .A1(Set_target[15]), .A2(n905), .B1(n906), .B2(
        \pc_target[6][15] ), .ZN(n929) );
  INV_X1 U1325 ( .A(n930), .ZN(n6314) );
  AOI22_X1 U1326 ( .A1(Set_target[17]), .A2(n905), .B1(n906), .B2(
        \pc_target[6][17] ), .ZN(n930) );
  INV_X1 U1327 ( .A(n931), .ZN(n6315) );
  AOI22_X1 U1328 ( .A1(Set_target[19]), .A2(n905), .B1(n906), .B2(
        \pc_target[6][19] ), .ZN(n931) );
  INV_X1 U1329 ( .A(n932), .ZN(n6316) );
  AOI22_X1 U1330 ( .A1(Set_target[21]), .A2(n905), .B1(n906), .B2(
        \pc_target[6][21] ), .ZN(n932) );
  INV_X1 U1331 ( .A(n933), .ZN(n6317) );
  AOI22_X1 U1332 ( .A1(Set_target[23]), .A2(n905), .B1(n906), .B2(
        \pc_target[6][23] ), .ZN(n933) );
  INV_X1 U1333 ( .A(n934), .ZN(n6318) );
  AOI22_X1 U1334 ( .A1(Set_target[25]), .A2(n905), .B1(n906), .B2(
        \pc_target[6][25] ), .ZN(n934) );
  INV_X1 U1335 ( .A(n935), .ZN(n6319) );
  AOI22_X1 U1336 ( .A1(Set_target[27]), .A2(n905), .B1(n906), .B2(
        \pc_target[6][27] ), .ZN(n935) );
  INV_X1 U1337 ( .A(n936), .ZN(n6320) );
  AOI22_X1 U1338 ( .A1(Set_target[29]), .A2(n905), .B1(n906), .B2(
        \pc_target[6][29] ), .ZN(n936) );
  INV_X1 U1339 ( .A(n937), .ZN(n6321) );
  AOI22_X1 U1340 ( .A1(Set_target[31]), .A2(n905), .B1(n906), .B2(
        \pc_target[6][31] ), .ZN(n937) );
  OAI22_X1 U1343 ( .A1(n75), .A2(n938), .B1(n939), .B2(n940), .ZN(n6322) );
  OAI22_X1 U1344 ( .A1(n79), .A2(n938), .B1(n939), .B2(n941), .ZN(n6323) );
  OAI22_X1 U1345 ( .A1(n81), .A2(n938), .B1(n939), .B2(n942), .ZN(n6324) );
  OAI22_X1 U1346 ( .A1(n83), .A2(n938), .B1(n939), .B2(n943), .ZN(n6325) );
  OAI22_X1 U1347 ( .A1(n85), .A2(n938), .B1(n939), .B2(n944), .ZN(n6326) );
  OAI22_X1 U1348 ( .A1(n87), .A2(n938), .B1(n939), .B2(n945), .ZN(n6327) );
  OAI22_X1 U1349 ( .A1(n89), .A2(n938), .B1(n939), .B2(n946), .ZN(n6328) );
  OAI22_X1 U1350 ( .A1(n91), .A2(n938), .B1(n939), .B2(n947), .ZN(n6329) );
  OAI22_X1 U1351 ( .A1(n93), .A2(n938), .B1(n939), .B2(n948), .ZN(n6330) );
  OAI22_X1 U1352 ( .A1(n95), .A2(n938), .B1(n939), .B2(n949), .ZN(n6331) );
  OAI22_X1 U1353 ( .A1(n97), .A2(n938), .B1(n939), .B2(n950), .ZN(n6332) );
  OAI22_X1 U1354 ( .A1(n99), .A2(n938), .B1(n939), .B2(n951), .ZN(n6333) );
  OAI22_X1 U1355 ( .A1(n101), .A2(n938), .B1(n939), .B2(n952), .ZN(n6334) );
  OAI22_X1 U1356 ( .A1(n103), .A2(n938), .B1(n939), .B2(n953), .ZN(n6335) );
  OAI22_X1 U1357 ( .A1(n105), .A2(n938), .B1(n939), .B2(n954), .ZN(n6336) );
  OAI22_X1 U1358 ( .A1(n107), .A2(n938), .B1(n939), .B2(n955), .ZN(n6337) );
  OAI22_X1 U1359 ( .A1(n109), .A2(n938), .B1(n939), .B2(n956), .ZN(n6338) );
  OAI22_X1 U1360 ( .A1(n111), .A2(n938), .B1(n939), .B2(n957), .ZN(n6339) );
  OAI22_X1 U1361 ( .A1(n113), .A2(n938), .B1(n939), .B2(n958), .ZN(n6340) );
  OAI22_X1 U1362 ( .A1(n115), .A2(n938), .B1(n939), .B2(n959), .ZN(n6341) );
  OAI22_X1 U1363 ( .A1(n117), .A2(n938), .B1(n939), .B2(n960), .ZN(n6342) );
  OAI22_X1 U1364 ( .A1(n119), .A2(n938), .B1(n939), .B2(n961), .ZN(n6343) );
  OAI22_X1 U1365 ( .A1(n121), .A2(n938), .B1(n939), .B2(n962), .ZN(n6344) );
  OAI22_X1 U1366 ( .A1(n123), .A2(n938), .B1(n939), .B2(n963), .ZN(n6345) );
  OAI22_X1 U1367 ( .A1(n125), .A2(n938), .B1(n939), .B2(n964), .ZN(n6346) );
  OAI22_X1 U1368 ( .A1(n127), .A2(n938), .B1(n939), .B2(n965), .ZN(n6347) );
  OAI22_X1 U1369 ( .A1(n129), .A2(n938), .B1(n939), .B2(n966), .ZN(n6348) );
  OAI22_X1 U1370 ( .A1(n131), .A2(n938), .B1(n939), .B2(n967), .ZN(n6349) );
  OAI22_X1 U1371 ( .A1(n133), .A2(n938), .B1(n939), .B2(n968), .ZN(n6350) );
  OAI22_X1 U1372 ( .A1(n135), .A2(n938), .B1(n939), .B2(n969), .ZN(n6351) );
  OAI22_X1 U1373 ( .A1(n137), .A2(n938), .B1(n939), .B2(n970), .ZN(n6352) );
  OAI22_X1 U1374 ( .A1(n139), .A2(n938), .B1(n939), .B2(n971), .ZN(n6353) );
  OAI22_X1 U1377 ( .A1(n75), .A2(n972), .B1(n3443), .B2(n974), .ZN(n6354) );
  OAI22_X1 U1378 ( .A1(n79), .A2(n972), .B1(n3443), .B2(n975), .ZN(n6355) );
  OAI22_X1 U1379 ( .A1(n81), .A2(n972), .B1(n3443), .B2(n976), .ZN(n6356) );
  OAI22_X1 U1380 ( .A1(n83), .A2(n972), .B1(n3443), .B2(n977), .ZN(n6357) );
  OAI22_X1 U1381 ( .A1(n85), .A2(n972), .B1(n3443), .B2(n978), .ZN(n6358) );
  OAI22_X1 U1382 ( .A1(n87), .A2(n972), .B1(n3443), .B2(n979), .ZN(n6359) );
  OAI22_X1 U1383 ( .A1(n89), .A2(n972), .B1(n3443), .B2(n980), .ZN(n6360) );
  OAI22_X1 U1384 ( .A1(n91), .A2(n972), .B1(n3443), .B2(n981), .ZN(n6361) );
  OAI22_X1 U1385 ( .A1(n93), .A2(n972), .B1(n3443), .B2(n982), .ZN(n6362) );
  OAI22_X1 U1386 ( .A1(n95), .A2(n972), .B1(n3443), .B2(n983), .ZN(n6363) );
  OAI22_X1 U1387 ( .A1(n97), .A2(n972), .B1(n3443), .B2(n984), .ZN(n6364) );
  OAI22_X1 U1388 ( .A1(n99), .A2(n972), .B1(n3443), .B2(n985), .ZN(n6365) );
  OAI22_X1 U1389 ( .A1(n101), .A2(n972), .B1(n3443), .B2(n986), .ZN(n6366) );
  OAI22_X1 U1390 ( .A1(n103), .A2(n972), .B1(n3443), .B2(n987), .ZN(n6367) );
  OAI22_X1 U1391 ( .A1(n105), .A2(n972), .B1(n3443), .B2(n988), .ZN(n6368) );
  OAI22_X1 U1392 ( .A1(n107), .A2(n972), .B1(n3443), .B2(n989), .ZN(n6369) );
  OAI22_X1 U1393 ( .A1(n109), .A2(n972), .B1(n3443), .B2(n990), .ZN(n6370) );
  OAI22_X1 U1394 ( .A1(n111), .A2(n972), .B1(n3443), .B2(n991), .ZN(n6371) );
  OAI22_X1 U1395 ( .A1(n113), .A2(n972), .B1(n3443), .B2(n992), .ZN(n6372) );
  OAI22_X1 U1396 ( .A1(n115), .A2(n972), .B1(n3443), .B2(n993), .ZN(n6373) );
  OAI22_X1 U1397 ( .A1(n117), .A2(n972), .B1(n3443), .B2(n994), .ZN(n6374) );
  OAI22_X1 U1398 ( .A1(n119), .A2(n972), .B1(n3443), .B2(n995), .ZN(n6375) );
  OAI22_X1 U1399 ( .A1(n121), .A2(n972), .B1(n3443), .B2(n996), .ZN(n6376) );
  OAI22_X1 U1400 ( .A1(n123), .A2(n972), .B1(n3443), .B2(n997), .ZN(n6377) );
  OAI22_X1 U1401 ( .A1(n125), .A2(n972), .B1(n3443), .B2(n998), .ZN(n6378) );
  OAI22_X1 U1402 ( .A1(n127), .A2(n972), .B1(n3443), .B2(n999), .ZN(n6379) );
  OAI22_X1 U1403 ( .A1(n129), .A2(n972), .B1(n3443), .B2(n1000), .ZN(n6380) );
  OAI22_X1 U1404 ( .A1(n131), .A2(n972), .B1(n3443), .B2(n1001), .ZN(n6381) );
  OAI22_X1 U1405 ( .A1(n133), .A2(n972), .B1(n3443), .B2(n1002), .ZN(n6382) );
  OAI22_X1 U1406 ( .A1(n135), .A2(n972), .B1(n3443), .B2(n1003), .ZN(n6383) );
  OAI22_X1 U1407 ( .A1(n137), .A2(n972), .B1(n3443), .B2(n1004), .ZN(n6384) );
  OAI22_X1 U1408 ( .A1(n139), .A2(n972), .B1(n3443), .B2(n1005), .ZN(n6385) );
  INV_X1 U1412 ( .A(n1006), .ZN(n6386) );
  AOI22_X1 U1413 ( .A1(Set_target[30]), .A2(n1007), .B1(n1008), .B2(
        \pc_target[3][30] ), .ZN(n1006) );
  INV_X1 U1414 ( .A(n1009), .ZN(n6387) );
  AOI22_X1 U1415 ( .A1(Set_target[28]), .A2(n1007), .B1(n1008), .B2(
        \pc_target[3][28] ), .ZN(n1009) );
  INV_X1 U1416 ( .A(n1010), .ZN(n6388) );
  AOI22_X1 U1417 ( .A1(Set_target[26]), .A2(n1007), .B1(n1008), .B2(
        \pc_target[3][26] ), .ZN(n1010) );
  INV_X1 U1418 ( .A(n1011), .ZN(n6389) );
  AOI22_X1 U1419 ( .A1(Set_target[24]), .A2(n1007), .B1(n1008), .B2(
        \pc_target[3][24] ), .ZN(n1011) );
  INV_X1 U1420 ( .A(n1012), .ZN(n6390) );
  AOI22_X1 U1421 ( .A1(Set_target[22]), .A2(n1007), .B1(n1008), .B2(
        \pc_target[3][22] ), .ZN(n1012) );
  INV_X1 U1422 ( .A(n1013), .ZN(n6391) );
  AOI22_X1 U1423 ( .A1(Set_target[20]), .A2(n1007), .B1(n1008), .B2(
        \pc_target[3][20] ), .ZN(n1013) );
  INV_X1 U1424 ( .A(n1014), .ZN(n6392) );
  AOI22_X1 U1425 ( .A1(Set_target[18]), .A2(n1007), .B1(n1008), .B2(
        \pc_target[3][18] ), .ZN(n1014) );
  INV_X1 U1426 ( .A(n1015), .ZN(n6393) );
  AOI22_X1 U1427 ( .A1(Set_target[16]), .A2(n1007), .B1(n1008), .B2(
        \pc_target[3][16] ), .ZN(n1015) );
  INV_X1 U1428 ( .A(n1016), .ZN(n6394) );
  AOI22_X1 U1429 ( .A1(Set_target[14]), .A2(n1007), .B1(n1008), .B2(
        \pc_target[3][14] ), .ZN(n1016) );
  INV_X1 U1430 ( .A(n1017), .ZN(n6395) );
  AOI22_X1 U1431 ( .A1(Set_target[12]), .A2(n1007), .B1(n1008), .B2(
        \pc_target[3][12] ), .ZN(n1017) );
  INV_X1 U1432 ( .A(n1018), .ZN(n6396) );
  AOI22_X1 U1433 ( .A1(Set_target[10]), .A2(n1007), .B1(n1008), .B2(
        \pc_target[3][10] ), .ZN(n1018) );
  INV_X1 U1434 ( .A(n1019), .ZN(n6397) );
  AOI22_X1 U1435 ( .A1(Set_target[8]), .A2(n1007), .B1(n1008), .B2(
        \pc_target[3][8] ), .ZN(n1019) );
  INV_X1 U1436 ( .A(n1020), .ZN(n6398) );
  AOI22_X1 U1437 ( .A1(Set_target[6]), .A2(n1007), .B1(n1008), .B2(
        \pc_target[3][6] ), .ZN(n1020) );
  INV_X1 U1438 ( .A(n1021), .ZN(n6399) );
  AOI22_X1 U1439 ( .A1(Set_target[4]), .A2(n1007), .B1(n1008), .B2(
        \pc_target[3][4] ), .ZN(n1021) );
  INV_X1 U1440 ( .A(n1022), .ZN(n6400) );
  AOI22_X1 U1441 ( .A1(Set_target[2]), .A2(n1007), .B1(n1008), .B2(
        \pc_target[3][2] ), .ZN(n1022) );
  INV_X1 U1442 ( .A(n1023), .ZN(n6401) );
  AOI22_X1 U1443 ( .A1(Set_target[0]), .A2(n1007), .B1(n1008), .B2(
        \pc_target[3][0] ), .ZN(n1023) );
  INV_X1 U1444 ( .A(n1024), .ZN(n6402) );
  AOI22_X1 U1445 ( .A1(Set_target[1]), .A2(n1007), .B1(n1008), .B2(
        \pc_target[3][1] ), .ZN(n1024) );
  INV_X1 U1446 ( .A(n1025), .ZN(n6403) );
  AOI22_X1 U1447 ( .A1(Set_target[3]), .A2(n1007), .B1(n1008), .B2(
        \pc_target[3][3] ), .ZN(n1025) );
  INV_X1 U1448 ( .A(n1026), .ZN(n6404) );
  AOI22_X1 U1449 ( .A1(Set_target[5]), .A2(n1007), .B1(n1008), .B2(
        \pc_target[3][5] ), .ZN(n1026) );
  INV_X1 U1450 ( .A(n1027), .ZN(n6405) );
  AOI22_X1 U1451 ( .A1(Set_target[7]), .A2(n1007), .B1(n1008), .B2(
        \pc_target[3][7] ), .ZN(n1027) );
  INV_X1 U1452 ( .A(n1028), .ZN(n6406) );
  AOI22_X1 U1453 ( .A1(Set_target[9]), .A2(n1007), .B1(n1008), .B2(
        \pc_target[3][9] ), .ZN(n1028) );
  INV_X1 U1454 ( .A(n1029), .ZN(n6407) );
  AOI22_X1 U1455 ( .A1(Set_target[11]), .A2(n1007), .B1(n1008), .B2(
        \pc_target[3][11] ), .ZN(n1029) );
  INV_X1 U1456 ( .A(n1030), .ZN(n6408) );
  AOI22_X1 U1457 ( .A1(Set_target[13]), .A2(n1007), .B1(n1008), .B2(
        \pc_target[3][13] ), .ZN(n1030) );
  INV_X1 U1458 ( .A(n1031), .ZN(n6409) );
  AOI22_X1 U1459 ( .A1(Set_target[15]), .A2(n1007), .B1(n1008), .B2(
        \pc_target[3][15] ), .ZN(n1031) );
  INV_X1 U1460 ( .A(n1032), .ZN(n6410) );
  AOI22_X1 U1461 ( .A1(Set_target[17]), .A2(n1007), .B1(n1008), .B2(
        \pc_target[3][17] ), .ZN(n1032) );
  INV_X1 U1462 ( .A(n1033), .ZN(n6411) );
  AOI22_X1 U1463 ( .A1(Set_target[19]), .A2(n1007), .B1(n1008), .B2(
        \pc_target[3][19] ), .ZN(n1033) );
  INV_X1 U1464 ( .A(n1034), .ZN(n6412) );
  AOI22_X1 U1465 ( .A1(Set_target[21]), .A2(n1007), .B1(n1008), .B2(
        \pc_target[3][21] ), .ZN(n1034) );
  INV_X1 U1466 ( .A(n1035), .ZN(n6413) );
  AOI22_X1 U1467 ( .A1(Set_target[23]), .A2(n1007), .B1(n1008), .B2(
        \pc_target[3][23] ), .ZN(n1035) );
  INV_X1 U1468 ( .A(n1036), .ZN(n6414) );
  AOI22_X1 U1469 ( .A1(Set_target[25]), .A2(n1007), .B1(n1008), .B2(
        \pc_target[3][25] ), .ZN(n1036) );
  INV_X1 U1470 ( .A(n1037), .ZN(n6415) );
  AOI22_X1 U1471 ( .A1(Set_target[27]), .A2(n1007), .B1(n1008), .B2(
        \pc_target[3][27] ), .ZN(n1037) );
  INV_X1 U1472 ( .A(n1038), .ZN(n6416) );
  AOI22_X1 U1473 ( .A1(Set_target[29]), .A2(n1007), .B1(n1008), .B2(
        \pc_target[3][29] ), .ZN(n1038) );
  INV_X1 U1474 ( .A(n1039), .ZN(n6417) );
  AOI22_X1 U1475 ( .A1(Set_target[31]), .A2(n1007), .B1(n1008), .B2(
        \pc_target[3][31] ), .ZN(n1039) );
  INV_X1 U1478 ( .A(n1041), .ZN(n6418) );
  AOI22_X1 U1479 ( .A1(Set_target[30]), .A2(n1042), .B1(n1043), .B2(
        \pc_target[2][30] ), .ZN(n1041) );
  INV_X1 U1480 ( .A(n1044), .ZN(n6419) );
  AOI22_X1 U1481 ( .A1(Set_target[28]), .A2(n1042), .B1(n1043), .B2(
        \pc_target[2][28] ), .ZN(n1044) );
  INV_X1 U1482 ( .A(n1045), .ZN(n6420) );
  AOI22_X1 U1483 ( .A1(Set_target[26]), .A2(n1042), .B1(n1043), .B2(
        \pc_target[2][26] ), .ZN(n1045) );
  INV_X1 U1484 ( .A(n1046), .ZN(n6421) );
  AOI22_X1 U1485 ( .A1(Set_target[24]), .A2(n1042), .B1(n1043), .B2(
        \pc_target[2][24] ), .ZN(n1046) );
  INV_X1 U1486 ( .A(n1047), .ZN(n6422) );
  AOI22_X1 U1487 ( .A1(Set_target[22]), .A2(n1042), .B1(n1043), .B2(
        \pc_target[2][22] ), .ZN(n1047) );
  INV_X1 U1488 ( .A(n1048), .ZN(n6423) );
  AOI22_X1 U1489 ( .A1(Set_target[20]), .A2(n1042), .B1(n1043), .B2(
        \pc_target[2][20] ), .ZN(n1048) );
  INV_X1 U1490 ( .A(n1049), .ZN(n6424) );
  AOI22_X1 U1491 ( .A1(Set_target[18]), .A2(n1042), .B1(n1043), .B2(
        \pc_target[2][18] ), .ZN(n1049) );
  INV_X1 U1492 ( .A(n1050), .ZN(n6425) );
  AOI22_X1 U1493 ( .A1(Set_target[16]), .A2(n1042), .B1(n1043), .B2(
        \pc_target[2][16] ), .ZN(n1050) );
  INV_X1 U1494 ( .A(n1051), .ZN(n6426) );
  AOI22_X1 U1495 ( .A1(Set_target[14]), .A2(n1042), .B1(n1043), .B2(
        \pc_target[2][14] ), .ZN(n1051) );
  INV_X1 U1496 ( .A(n1052), .ZN(n6427) );
  AOI22_X1 U1497 ( .A1(Set_target[12]), .A2(n1042), .B1(n1043), .B2(
        \pc_target[2][12] ), .ZN(n1052) );
  INV_X1 U1498 ( .A(n1053), .ZN(n6428) );
  AOI22_X1 U1499 ( .A1(Set_target[10]), .A2(n1042), .B1(n1043), .B2(
        \pc_target[2][10] ), .ZN(n1053) );
  INV_X1 U1500 ( .A(n1054), .ZN(n6429) );
  AOI22_X1 U1501 ( .A1(Set_target[8]), .A2(n1042), .B1(n1043), .B2(
        \pc_target[2][8] ), .ZN(n1054) );
  INV_X1 U1502 ( .A(n1055), .ZN(n6430) );
  AOI22_X1 U1503 ( .A1(Set_target[6]), .A2(n1042), .B1(n1043), .B2(
        \pc_target[2][6] ), .ZN(n1055) );
  INV_X1 U1504 ( .A(n1056), .ZN(n6431) );
  AOI22_X1 U1505 ( .A1(Set_target[4]), .A2(n1042), .B1(n1043), .B2(
        \pc_target[2][4] ), .ZN(n1056) );
  INV_X1 U1506 ( .A(n1057), .ZN(n6432) );
  AOI22_X1 U1507 ( .A1(Set_target[2]), .A2(n1042), .B1(n1043), .B2(
        \pc_target[2][2] ), .ZN(n1057) );
  INV_X1 U1508 ( .A(n1058), .ZN(n6433) );
  AOI22_X1 U1509 ( .A1(Set_target[0]), .A2(n1042), .B1(n1043), .B2(
        \pc_target[2][0] ), .ZN(n1058) );
  INV_X1 U1510 ( .A(n1059), .ZN(n6434) );
  AOI22_X1 U1511 ( .A1(Set_target[1]), .A2(n1042), .B1(n1043), .B2(
        \pc_target[2][1] ), .ZN(n1059) );
  INV_X1 U1512 ( .A(n1060), .ZN(n6435) );
  AOI22_X1 U1513 ( .A1(Set_target[3]), .A2(n1042), .B1(n1043), .B2(
        \pc_target[2][3] ), .ZN(n1060) );
  INV_X1 U1514 ( .A(n1061), .ZN(n6436) );
  AOI22_X1 U1515 ( .A1(Set_target[5]), .A2(n1042), .B1(n1043), .B2(
        \pc_target[2][5] ), .ZN(n1061) );
  INV_X1 U1516 ( .A(n1062), .ZN(n6437) );
  AOI22_X1 U1517 ( .A1(Set_target[7]), .A2(n1042), .B1(n1043), .B2(
        \pc_target[2][7] ), .ZN(n1062) );
  INV_X1 U1518 ( .A(n1063), .ZN(n6438) );
  AOI22_X1 U1519 ( .A1(Set_target[9]), .A2(n1042), .B1(n1043), .B2(
        \pc_target[2][9] ), .ZN(n1063) );
  INV_X1 U1520 ( .A(n1064), .ZN(n6439) );
  AOI22_X1 U1521 ( .A1(Set_target[11]), .A2(n1042), .B1(n1043), .B2(
        \pc_target[2][11] ), .ZN(n1064) );
  INV_X1 U1522 ( .A(n1065), .ZN(n6440) );
  AOI22_X1 U1523 ( .A1(Set_target[13]), .A2(n1042), .B1(n1043), .B2(
        \pc_target[2][13] ), .ZN(n1065) );
  INV_X1 U1524 ( .A(n1066), .ZN(n6441) );
  AOI22_X1 U1525 ( .A1(Set_target[15]), .A2(n1042), .B1(n1043), .B2(
        \pc_target[2][15] ), .ZN(n1066) );
  INV_X1 U1526 ( .A(n1067), .ZN(n6442) );
  AOI22_X1 U1527 ( .A1(Set_target[17]), .A2(n1042), .B1(n1043), .B2(
        \pc_target[2][17] ), .ZN(n1067) );
  INV_X1 U1528 ( .A(n1068), .ZN(n6443) );
  AOI22_X1 U1529 ( .A1(Set_target[19]), .A2(n1042), .B1(n1043), .B2(
        \pc_target[2][19] ), .ZN(n1068) );
  INV_X1 U1530 ( .A(n1069), .ZN(n6444) );
  AOI22_X1 U1531 ( .A1(Set_target[21]), .A2(n1042), .B1(n1043), .B2(
        \pc_target[2][21] ), .ZN(n1069) );
  INV_X1 U1532 ( .A(n1070), .ZN(n6445) );
  AOI22_X1 U1533 ( .A1(Set_target[23]), .A2(n1042), .B1(n1043), .B2(
        \pc_target[2][23] ), .ZN(n1070) );
  INV_X1 U1534 ( .A(n1071), .ZN(n6446) );
  AOI22_X1 U1535 ( .A1(Set_target[25]), .A2(n1042), .B1(n1043), .B2(
        \pc_target[2][25] ), .ZN(n1071) );
  INV_X1 U1536 ( .A(n1072), .ZN(n6447) );
  AOI22_X1 U1537 ( .A1(Set_target[27]), .A2(n1042), .B1(n1043), .B2(
        \pc_target[2][27] ), .ZN(n1072) );
  INV_X1 U1538 ( .A(n1073), .ZN(n6448) );
  AOI22_X1 U1539 ( .A1(Set_target[29]), .A2(n1042), .B1(n1043), .B2(
        \pc_target[2][29] ), .ZN(n1073) );
  INV_X1 U1540 ( .A(n1074), .ZN(n6449) );
  AOI22_X1 U1541 ( .A1(Set_target[31]), .A2(n1042), .B1(n1043), .B2(
        \pc_target[2][31] ), .ZN(n1074) );
  OAI22_X1 U1544 ( .A1(n75), .A2(n1075), .B1(n1076), .B2(n1077), .ZN(n6450) );
  OAI22_X1 U1545 ( .A1(n79), .A2(n1075), .B1(n1076), .B2(n1078), .ZN(n6451) );
  OAI22_X1 U1546 ( .A1(n81), .A2(n1075), .B1(n1076), .B2(n1079), .ZN(n6452) );
  OAI22_X1 U1547 ( .A1(n83), .A2(n1075), .B1(n1076), .B2(n1080), .ZN(n6453) );
  OAI22_X1 U1548 ( .A1(n85), .A2(n1075), .B1(n1076), .B2(n1081), .ZN(n6454) );
  OAI22_X1 U1549 ( .A1(n87), .A2(n1075), .B1(n1076), .B2(n1082), .ZN(n6455) );
  OAI22_X1 U1550 ( .A1(n89), .A2(n1075), .B1(n1076), .B2(n1083), .ZN(n6456) );
  OAI22_X1 U1551 ( .A1(n91), .A2(n1075), .B1(n1076), .B2(n1084), .ZN(n6457) );
  OAI22_X1 U1552 ( .A1(n93), .A2(n1075), .B1(n1076), .B2(n1085), .ZN(n6458) );
  OAI22_X1 U1553 ( .A1(n95), .A2(n1075), .B1(n1076), .B2(n1086), .ZN(n6459) );
  OAI22_X1 U1554 ( .A1(n97), .A2(n1075), .B1(n1076), .B2(n1087), .ZN(n6460) );
  OAI22_X1 U1555 ( .A1(n99), .A2(n1075), .B1(n1076), .B2(n1088), .ZN(n6461) );
  OAI22_X1 U1556 ( .A1(n101), .A2(n1075), .B1(n1076), .B2(n1089), .ZN(n6462)
         );
  OAI22_X1 U1557 ( .A1(n103), .A2(n1075), .B1(n1076), .B2(n1090), .ZN(n6463)
         );
  OAI22_X1 U1558 ( .A1(n105), .A2(n1075), .B1(n1076), .B2(n1091), .ZN(n6464)
         );
  OAI22_X1 U1559 ( .A1(n107), .A2(n1075), .B1(n1076), .B2(n1092), .ZN(n6465)
         );
  OAI22_X1 U1560 ( .A1(n109), .A2(n1075), .B1(n1076), .B2(n1093), .ZN(n6466)
         );
  OAI22_X1 U1561 ( .A1(n111), .A2(n1075), .B1(n1076), .B2(n1094), .ZN(n6467)
         );
  OAI22_X1 U1562 ( .A1(n113), .A2(n1075), .B1(n1076), .B2(n1095), .ZN(n6468)
         );
  OAI22_X1 U1563 ( .A1(n115), .A2(n1075), .B1(n1076), .B2(n1096), .ZN(n6469)
         );
  OAI22_X1 U1564 ( .A1(n117), .A2(n1075), .B1(n1076), .B2(n1097), .ZN(n6470)
         );
  OAI22_X1 U1565 ( .A1(n119), .A2(n1075), .B1(n1076), .B2(n1098), .ZN(n6471)
         );
  OAI22_X1 U1566 ( .A1(n121), .A2(n1075), .B1(n1076), .B2(n1099), .ZN(n6472)
         );
  OAI22_X1 U1567 ( .A1(n123), .A2(n1075), .B1(n1076), .B2(n1100), .ZN(n6473)
         );
  OAI22_X1 U1568 ( .A1(n125), .A2(n1075), .B1(n1076), .B2(n1101), .ZN(n6474)
         );
  OAI22_X1 U1569 ( .A1(n127), .A2(n1075), .B1(n1076), .B2(n1102), .ZN(n6475)
         );
  OAI22_X1 U1570 ( .A1(n129), .A2(n1075), .B1(n1076), .B2(n1103), .ZN(n6476)
         );
  OAI22_X1 U1571 ( .A1(n131), .A2(n1075), .B1(n1076), .B2(n1104), .ZN(n6477)
         );
  OAI22_X1 U1572 ( .A1(n133), .A2(n1075), .B1(n1076), .B2(n1105), .ZN(n6478)
         );
  OAI22_X1 U1573 ( .A1(n135), .A2(n1075), .B1(n1076), .B2(n1106), .ZN(n6479)
         );
  OAI22_X1 U1574 ( .A1(n137), .A2(n1075), .B1(n1076), .B2(n1107), .ZN(n6480)
         );
  OAI22_X1 U1575 ( .A1(n139), .A2(n1075), .B1(n1076), .B2(n1108), .ZN(n6481)
         );
  OAI22_X1 U1578 ( .A1(n75), .A2(n1109), .B1(n1110), .B2(n1111), .ZN(n6482) );
  OAI22_X1 U1580 ( .A1(n79), .A2(n1109), .B1(n1110), .B2(n1112), .ZN(n6483) );
  OAI22_X1 U1582 ( .A1(n81), .A2(n1109), .B1(n1110), .B2(n1113), .ZN(n6484) );
  OAI22_X1 U1584 ( .A1(n83), .A2(n1109), .B1(n1110), .B2(n1114), .ZN(n6485) );
  OAI22_X1 U1586 ( .A1(n85), .A2(n1109), .B1(n1110), .B2(n1115), .ZN(n6486) );
  OAI22_X1 U1588 ( .A1(n87), .A2(n1109), .B1(n1110), .B2(n1116), .ZN(n6487) );
  OAI22_X1 U1590 ( .A1(n89), .A2(n1109), .B1(n1110), .B2(n1117), .ZN(n6488) );
  OAI22_X1 U1592 ( .A1(n91), .A2(n1109), .B1(n1110), .B2(n1118), .ZN(n6489) );
  OAI22_X1 U1594 ( .A1(n93), .A2(n1109), .B1(n1110), .B2(n1119), .ZN(n6490) );
  OAI22_X1 U1596 ( .A1(n95), .A2(n1109), .B1(n1110), .B2(n1120), .ZN(n6491) );
  OAI22_X1 U1598 ( .A1(n97), .A2(n1109), .B1(n1110), .B2(n1121), .ZN(n6492) );
  INV_X1 U1599 ( .A(Set_target[10]), .ZN(n97) );
  OAI22_X1 U1600 ( .A1(n99), .A2(n1109), .B1(n1110), .B2(n1122), .ZN(n6493) );
  INV_X1 U1601 ( .A(Set_target[8]), .ZN(n99) );
  OAI22_X1 U1602 ( .A1(n101), .A2(n1109), .B1(n1110), .B2(n1123), .ZN(n6494)
         );
  INV_X1 U1603 ( .A(Set_target[6]), .ZN(n101) );
  OAI22_X1 U1604 ( .A1(n103), .A2(n1109), .B1(n1110), .B2(n1124), .ZN(n6495)
         );
  INV_X1 U1605 ( .A(Set_target[4]), .ZN(n103) );
  OAI22_X1 U1606 ( .A1(n105), .A2(n1109), .B1(n1110), .B2(n1125), .ZN(n6496)
         );
  INV_X1 U1607 ( .A(Set_target[2]), .ZN(n105) );
  OAI22_X1 U1608 ( .A1(n107), .A2(n1109), .B1(n1110), .B2(n1126), .ZN(n6497)
         );
  INV_X1 U1609 ( .A(Set_target[0]), .ZN(n107) );
  OAI22_X1 U1610 ( .A1(n109), .A2(n1109), .B1(n1110), .B2(n1127), .ZN(n6498)
         );
  INV_X1 U1611 ( .A(Set_target[1]), .ZN(n109) );
  OAI22_X1 U1612 ( .A1(n111), .A2(n1109), .B1(n1110), .B2(n1128), .ZN(n6499)
         );
  INV_X1 U1613 ( .A(Set_target[3]), .ZN(n111) );
  OAI22_X1 U1614 ( .A1(n113), .A2(n1109), .B1(n1110), .B2(n1129), .ZN(n6500)
         );
  INV_X1 U1615 ( .A(Set_target[5]), .ZN(n113) );
  OAI22_X1 U1616 ( .A1(n115), .A2(n1109), .B1(n1110), .B2(n1130), .ZN(n6501)
         );
  INV_X1 U1617 ( .A(Set_target[7]), .ZN(n115) );
  OAI22_X1 U1618 ( .A1(n117), .A2(n1109), .B1(n1110), .B2(n1131), .ZN(n6502)
         );
  INV_X1 U1619 ( .A(Set_target[9]), .ZN(n117) );
  OAI22_X1 U1620 ( .A1(n119), .A2(n1109), .B1(n1110), .B2(n1132), .ZN(n6503)
         );
  OAI22_X1 U1622 ( .A1(n121), .A2(n1109), .B1(n1110), .B2(n1133), .ZN(n6504)
         );
  OAI22_X1 U1624 ( .A1(n123), .A2(n1109), .B1(n1110), .B2(n1134), .ZN(n6505)
         );
  OAI22_X1 U1626 ( .A1(n125), .A2(n1109), .B1(n1110), .B2(n1135), .ZN(n6506)
         );
  OAI22_X1 U1628 ( .A1(n127), .A2(n1109), .B1(n1110), .B2(n1136), .ZN(n6507)
         );
  OAI22_X1 U1630 ( .A1(n129), .A2(n1109), .B1(n1110), .B2(n1137), .ZN(n6508)
         );
  OAI22_X1 U1632 ( .A1(n131), .A2(n1109), .B1(n1110), .B2(n1138), .ZN(n6509)
         );
  OAI22_X1 U1634 ( .A1(n133), .A2(n1109), .B1(n1110), .B2(n1139), .ZN(n6510)
         );
  OAI22_X1 U1636 ( .A1(n135), .A2(n1109), .B1(n1110), .B2(n1140), .ZN(n6511)
         );
  OAI22_X1 U1638 ( .A1(n137), .A2(n1109), .B1(n1110), .B2(n1141), .ZN(n6512)
         );
  OAI22_X1 U1640 ( .A1(n139), .A2(n1109), .B1(n1110), .B2(n1142), .ZN(n6513)
         );
  INV_X1 U1646 ( .A(Set_target[31]), .ZN(n139) );
  OAI22_X1 U1647 ( .A1(n3808), .A2(n1146), .B1(n1147), .B2(n1148), .ZN(n6514)
         );
  OAI22_X1 U1649 ( .A1(n3808), .A2(n1149), .B1(n1148), .B2(n1150), .ZN(n6515)
         );
  OAI22_X1 U1651 ( .A1(n3809), .A2(n1151), .B1(n1148), .B2(n1152), .ZN(n6516)
         );
  OAI22_X1 U1653 ( .A1(n3809), .A2(n1153), .B1(n1148), .B2(n1154), .ZN(n6517)
         );
  OAI22_X1 U1655 ( .A1(n3808), .A2(n1155), .B1(n1148), .B2(n1156), .ZN(n6518)
         );
  OAI22_X1 U1657 ( .A1(n3808), .A2(n1157), .B1(n1148), .B2(n1158), .ZN(n6519)
         );
  OAI22_X1 U1659 ( .A1(n3809), .A2(n1159), .B1(n1148), .B2(n1160), .ZN(n6520)
         );
  OAI22_X1 U1661 ( .A1(n3809), .A2(n1161), .B1(n1148), .B2(n1162), .ZN(n6521)
         );
  OAI22_X1 U1663 ( .A1(n3809), .A2(n1163), .B1(n1148), .B2(n1164), .ZN(n6522)
         );
  OAI22_X1 U1665 ( .A1(n3808), .A2(n1165), .B1(n1148), .B2(n1166), .ZN(n6523)
         );
  OAI22_X1 U1667 ( .A1(n3809), .A2(n1167), .B1(n1148), .B2(n1168), .ZN(n6524)
         );
  OAI22_X1 U1669 ( .A1(n3809), .A2(n1169), .B1(n1148), .B2(n1170), .ZN(n6525)
         );
  OAI22_X1 U1671 ( .A1(n3809), .A2(n1171), .B1(n1148), .B2(n1172), .ZN(n6526)
         );
  INV_X1 U1673 ( .A(n1173), .ZN(n6527) );
  AOI22_X1 U1674 ( .A1(n1148), .A2(\pc_lut[31][4] ), .B1(n3521), .B2(n3809), 
        .ZN(n1173) );
  INV_X1 U1675 ( .A(n1174), .ZN(n6528) );
  AOI22_X1 U1676 ( .A1(n1148), .A2(\pc_lut[31][2] ), .B1(n3521), .B2(n3807), 
        .ZN(n1174) );
  INV_X1 U1677 ( .A(n1175), .ZN(n6529) );
  AOI22_X1 U1678 ( .A1(n1148), .A2(\pc_lut[31][0] ), .B1(n3521), .B2(n3807), 
        .ZN(n1175) );
  INV_X1 U1679 ( .A(n1176), .ZN(n6530) );
  AOI22_X1 U1680 ( .A1(n1148), .A2(\pc_lut[31][1] ), .B1(n3521), .B2(n3807), 
        .ZN(n1176) );
  INV_X1 U1681 ( .A(n1177), .ZN(n6531) );
  AOI22_X1 U1682 ( .A1(n1148), .A2(\pc_lut[31][3] ), .B1(n3521), .B2(n3807), 
        .ZN(n1177) );
  OAI22_X1 U1683 ( .A1(n3808), .A2(n1178), .B1(n1148), .B2(n1179), .ZN(n6532)
         );
  OAI22_X1 U1685 ( .A1(n3809), .A2(n1180), .B1(n1148), .B2(n1181), .ZN(n6533)
         );
  OAI22_X1 U1687 ( .A1(n3809), .A2(n1182), .B1(n1148), .B2(n1183), .ZN(n6534)
         );
  OAI22_X1 U1689 ( .A1(n3808), .A2(n1184), .B1(n1148), .B2(n1185), .ZN(n6535)
         );
  OAI22_X1 U1691 ( .A1(n3809), .A2(n1186), .B1(n1148), .B2(n1187), .ZN(n6536)
         );
  OAI22_X1 U1693 ( .A1(n3808), .A2(n1188), .B1(n1148), .B2(n1189), .ZN(n6537)
         );
  OAI22_X1 U1695 ( .A1(n3809), .A2(n1190), .B1(n1148), .B2(n1191), .ZN(n6538)
         );
  OAI22_X1 U1697 ( .A1(n3808), .A2(n1192), .B1(n1148), .B2(n1193), .ZN(n6539)
         );
  OAI22_X1 U1699 ( .A1(n3809), .A2(n1194), .B1(n1148), .B2(n1195), .ZN(n6540)
         );
  OAI22_X1 U1701 ( .A1(n3808), .A2(n1196), .B1(n1148), .B2(n1197), .ZN(n6541)
         );
  OAI22_X1 U1703 ( .A1(n3808), .A2(n1198), .B1(n1148), .B2(n1199), .ZN(n6542)
         );
  OAI22_X1 U1705 ( .A1(n3808), .A2(n1200), .B1(n1148), .B2(n1201), .ZN(n6543)
         );
  OAI22_X1 U1707 ( .A1(n3808), .A2(n1202), .B1(n1148), .B2(n1203), .ZN(n6544)
         );
  OAI22_X1 U1709 ( .A1(n3808), .A2(n1204), .B1(n1148), .B2(n1205), .ZN(n6545)
         );
  OAI22_X1 U1713 ( .A1(n3805), .A2(n1208), .B1(n1147), .B2(n1209), .ZN(n6546)
         );
  OAI22_X1 U1715 ( .A1(n3805), .A2(n1210), .B1(n1150), .B2(n1209), .ZN(n6547)
         );
  OAI22_X1 U1717 ( .A1(n3805), .A2(n1211), .B1(n1152), .B2(n1209), .ZN(n6548)
         );
  OAI22_X1 U1719 ( .A1(n3805), .A2(n1212), .B1(n1154), .B2(n1209), .ZN(n6549)
         );
  OAI22_X1 U1721 ( .A1(n3805), .A2(n1213), .B1(n1156), .B2(n1209), .ZN(n6550)
         );
  OAI22_X1 U1723 ( .A1(n3805), .A2(n1214), .B1(n1158), .B2(n1209), .ZN(n6551)
         );
  OAI22_X1 U1725 ( .A1(n3805), .A2(n1215), .B1(n1160), .B2(n1209), .ZN(n6552)
         );
  OAI22_X1 U1727 ( .A1(n3805), .A2(n1216), .B1(n1162), .B2(n1209), .ZN(n6553)
         );
  OAI22_X1 U1729 ( .A1(n3805), .A2(n1217), .B1(n1164), .B2(n1209), .ZN(n6554)
         );
  OAI22_X1 U1731 ( .A1(n3805), .A2(n1218), .B1(n1166), .B2(n1209), .ZN(n6555)
         );
  OAI22_X1 U1733 ( .A1(n3805), .A2(n1219), .B1(n1168), .B2(n1209), .ZN(n6556)
         );
  OAI22_X1 U1735 ( .A1(n3805), .A2(n1220), .B1(n1170), .B2(n1209), .ZN(n6557)
         );
  OAI22_X1 U1737 ( .A1(n3805), .A2(n1221), .B1(n1172), .B2(n1209), .ZN(n6558)
         );
  INV_X1 U1739 ( .A(n1222), .ZN(n6559) );
  AOI22_X1 U1740 ( .A1(n1209), .A2(\pc_lut[30][4] ), .B1(n3521), .B2(n3805), 
        .ZN(n1222) );
  INV_X1 U1741 ( .A(n1223), .ZN(n6560) );
  AOI22_X1 U1742 ( .A1(n1209), .A2(\pc_lut[30][2] ), .B1(n3521), .B2(n3805), 
        .ZN(n1223) );
  INV_X1 U1744 ( .A(n1224), .ZN(n6562) );
  AOI22_X1 U1745 ( .A1(n1209), .A2(\pc_lut[30][1] ), .B1(n3521), .B2(n3805), 
        .ZN(n1224) );
  INV_X1 U1746 ( .A(n1225), .ZN(n6563) );
  AOI22_X1 U1747 ( .A1(n1209), .A2(\pc_lut[30][3] ), .B1(n3521), .B2(n3805), 
        .ZN(n1225) );
  OAI22_X1 U1748 ( .A1(n3805), .A2(n1226), .B1(n1179), .B2(n1209), .ZN(n6564)
         );
  OAI22_X1 U1750 ( .A1(n3805), .A2(n1227), .B1(n1181), .B2(n1209), .ZN(n6565)
         );
  OAI22_X1 U1752 ( .A1(n3805), .A2(n1228), .B1(n1183), .B2(n1209), .ZN(n6566)
         );
  OAI22_X1 U1754 ( .A1(n3805), .A2(n1229), .B1(n1185), .B2(n1209), .ZN(n6567)
         );
  OAI22_X1 U1756 ( .A1(n3805), .A2(n1230), .B1(n1187), .B2(n1209), .ZN(n6568)
         );
  OAI22_X1 U1758 ( .A1(n3805), .A2(n1231), .B1(n1189), .B2(n1209), .ZN(n6569)
         );
  OAI22_X1 U1760 ( .A1(n3805), .A2(n1232), .B1(n1191), .B2(n1209), .ZN(n6570)
         );
  OAI22_X1 U1762 ( .A1(n3805), .A2(n1233), .B1(n1193), .B2(n1209), .ZN(n6571)
         );
  OAI22_X1 U1764 ( .A1(n3805), .A2(n1234), .B1(n1195), .B2(n1209), .ZN(n6572)
         );
  OAI22_X1 U1766 ( .A1(n3805), .A2(n1235), .B1(n1197), .B2(n1209), .ZN(n6573)
         );
  OAI22_X1 U1768 ( .A1(n3805), .A2(n1236), .B1(n1199), .B2(n1209), .ZN(n6574)
         );
  OAI22_X1 U1770 ( .A1(n3805), .A2(n1237), .B1(n1201), .B2(n1209), .ZN(n6575)
         );
  OAI22_X1 U1772 ( .A1(n3805), .A2(n1238), .B1(n1203), .B2(n1209), .ZN(n6576)
         );
  OAI22_X1 U1774 ( .A1(n3805), .A2(n1239), .B1(n1205), .B2(n1209), .ZN(n6577)
         );
  OAI22_X1 U1778 ( .A1(n3536), .A2(n1241), .B1(n1147), .B2(n1242), .ZN(n6578)
         );
  OAI22_X1 U1779 ( .A1(n3536), .A2(n1243), .B1(n1150), .B2(n1242), .ZN(n6579)
         );
  OAI22_X1 U1780 ( .A1(n3536), .A2(n1244), .B1(n1152), .B2(n1242), .ZN(n6580)
         );
  OAI22_X1 U1781 ( .A1(n3536), .A2(n1245), .B1(n1154), .B2(n1242), .ZN(n6581)
         );
  OAI22_X1 U1782 ( .A1(n3536), .A2(n1246), .B1(n1156), .B2(n1242), .ZN(n6582)
         );
  OAI22_X1 U1783 ( .A1(n3536), .A2(n1247), .B1(n1158), .B2(n1242), .ZN(n6583)
         );
  OAI22_X1 U1784 ( .A1(n3536), .A2(n1248), .B1(n1160), .B2(n1242), .ZN(n6584)
         );
  OAI22_X1 U1785 ( .A1(n3536), .A2(n1249), .B1(n1162), .B2(n1242), .ZN(n6585)
         );
  OAI22_X1 U1786 ( .A1(n3536), .A2(n1250), .B1(n1164), .B2(n1242), .ZN(n6586)
         );
  OAI22_X1 U1787 ( .A1(n3536), .A2(n1251), .B1(n1166), .B2(n1242), .ZN(n6587)
         );
  OAI22_X1 U1788 ( .A1(n3536), .A2(n1252), .B1(n1168), .B2(n1242), .ZN(n6588)
         );
  OAI22_X1 U1789 ( .A1(n3536), .A2(n1253), .B1(n1170), .B2(n1242), .ZN(n6589)
         );
  OAI22_X1 U1790 ( .A1(n3536), .A2(n1254), .B1(n1172), .B2(n1242), .ZN(n6590)
         );
  OAI22_X1 U1791 ( .A1(n3536), .A2(n1255), .B1(n1496), .B2(n1242), .ZN(n6591)
         );
  OAI22_X1 U1792 ( .A1(n3536), .A2(n1257), .B1(n1496), .B2(n1242), .ZN(n6592)
         );
  OAI22_X1 U1793 ( .A1(n3536), .A2(n1258), .B1(n1496), .B2(n1242), .ZN(n6593)
         );
  OAI22_X1 U1795 ( .A1(n3536), .A2(n1260), .B1(n1496), .B2(n1242), .ZN(n6595)
         );
  OAI22_X1 U1796 ( .A1(n3536), .A2(n1261), .B1(n1179), .B2(n1242), .ZN(n6596)
         );
  OAI22_X1 U1797 ( .A1(n3536), .A2(n1262), .B1(n1181), .B2(n1242), .ZN(n6597)
         );
  OAI22_X1 U1798 ( .A1(n3536), .A2(n1263), .B1(n1183), .B2(n1242), .ZN(n6598)
         );
  OAI22_X1 U1799 ( .A1(n3536), .A2(n1264), .B1(n1185), .B2(n1242), .ZN(n6599)
         );
  OAI22_X1 U1800 ( .A1(n3536), .A2(n1265), .B1(n1187), .B2(n1242), .ZN(n6600)
         );
  OAI22_X1 U1801 ( .A1(n3536), .A2(n1266), .B1(n1189), .B2(n1242), .ZN(n6601)
         );
  OAI22_X1 U1802 ( .A1(n3536), .A2(n1267), .B1(n1191), .B2(n1242), .ZN(n6602)
         );
  OAI22_X1 U1803 ( .A1(n3536), .A2(n1268), .B1(n1193), .B2(n1242), .ZN(n6603)
         );
  OAI22_X1 U1804 ( .A1(n3536), .A2(n1269), .B1(n1195), .B2(n1242), .ZN(n6604)
         );
  OAI22_X1 U1805 ( .A1(n3536), .A2(n1270), .B1(n1197), .B2(n1242), .ZN(n6605)
         );
  OAI22_X1 U1806 ( .A1(n3536), .A2(n1271), .B1(n1199), .B2(n1242), .ZN(n6606)
         );
  OAI22_X1 U1807 ( .A1(n3536), .A2(n1272), .B1(n1201), .B2(n1242), .ZN(n6607)
         );
  OAI22_X1 U1808 ( .A1(n3536), .A2(n1273), .B1(n1203), .B2(n1242), .ZN(n6608)
         );
  OAI22_X1 U1809 ( .A1(n3536), .A2(n1274), .B1(n1205), .B2(n1242), .ZN(n6609)
         );
  OAI22_X1 U1812 ( .A1(n3534), .A2(n1276), .B1(n1147), .B2(n1277), .ZN(n6610)
         );
  OAI22_X1 U1813 ( .A1(n3534), .A2(n1278), .B1(n1150), .B2(n1277), .ZN(n6611)
         );
  OAI22_X1 U1814 ( .A1(n3534), .A2(n1279), .B1(n1152), .B2(n1277), .ZN(n6612)
         );
  OAI22_X1 U1815 ( .A1(n3534), .A2(n1280), .B1(n1154), .B2(n1277), .ZN(n6613)
         );
  OAI22_X1 U1816 ( .A1(n3534), .A2(n1281), .B1(n1156), .B2(n1277), .ZN(n6614)
         );
  OAI22_X1 U1817 ( .A1(n3534), .A2(n1282), .B1(n1158), .B2(n1277), .ZN(n6615)
         );
  OAI22_X1 U1818 ( .A1(n3534), .A2(n1283), .B1(n1160), .B2(n1277), .ZN(n6616)
         );
  OAI22_X1 U1819 ( .A1(n3534), .A2(n1284), .B1(n1162), .B2(n1277), .ZN(n6617)
         );
  OAI22_X1 U1820 ( .A1(n3534), .A2(n1285), .B1(n1164), .B2(n1277), .ZN(n6618)
         );
  OAI22_X1 U1821 ( .A1(n3534), .A2(n1286), .B1(n1166), .B2(n1277), .ZN(n6619)
         );
  OAI22_X1 U1822 ( .A1(n3534), .A2(n1287), .B1(n1168), .B2(n1277), .ZN(n6620)
         );
  OAI22_X1 U1823 ( .A1(n3534), .A2(n1288), .B1(n1170), .B2(n1277), .ZN(n6621)
         );
  OAI22_X1 U1824 ( .A1(n3534), .A2(n1289), .B1(n1172), .B2(n1277), .ZN(n6622)
         );
  OAI22_X1 U1825 ( .A1(n3534), .A2(n1290), .B1(n1496), .B2(n1277), .ZN(n6623)
         );
  OAI22_X1 U1826 ( .A1(n3534), .A2(n1291), .B1(n1496), .B2(n1277), .ZN(n6624)
         );
  OAI22_X1 U1829 ( .A1(n3534), .A2(n1294), .B1(n1496), .B2(n1277), .ZN(n6627)
         );
  OAI22_X1 U1830 ( .A1(n3534), .A2(n1295), .B1(n1179), .B2(n1277), .ZN(n6628)
         );
  OAI22_X1 U1831 ( .A1(n3534), .A2(n1296), .B1(n1181), .B2(n1277), .ZN(n6629)
         );
  OAI22_X1 U1832 ( .A1(n3534), .A2(n1297), .B1(n1183), .B2(n1277), .ZN(n6630)
         );
  OAI22_X1 U1833 ( .A1(n3534), .A2(n1298), .B1(n1185), .B2(n1277), .ZN(n6631)
         );
  OAI22_X1 U1834 ( .A1(n3534), .A2(n1299), .B1(n1187), .B2(n1277), .ZN(n6632)
         );
  OAI22_X1 U1835 ( .A1(n3534), .A2(n1300), .B1(n1189), .B2(n1277), .ZN(n6633)
         );
  OAI22_X1 U1836 ( .A1(n3534), .A2(n1301), .B1(n1191), .B2(n1277), .ZN(n6634)
         );
  OAI22_X1 U1837 ( .A1(n3534), .A2(n1302), .B1(n1193), .B2(n1277), .ZN(n6635)
         );
  OAI22_X1 U1838 ( .A1(n3534), .A2(n1303), .B1(n1195), .B2(n1277), .ZN(n6636)
         );
  OAI22_X1 U1839 ( .A1(n3534), .A2(n1304), .B1(n1197), .B2(n1277), .ZN(n6637)
         );
  OAI22_X1 U1840 ( .A1(n3534), .A2(n1305), .B1(n1199), .B2(n1277), .ZN(n6638)
         );
  OAI22_X1 U1841 ( .A1(n3534), .A2(n1306), .B1(n1201), .B2(n1277), .ZN(n6639)
         );
  OAI22_X1 U1842 ( .A1(n3534), .A2(n1307), .B1(n1203), .B2(n1277), .ZN(n6640)
         );
  OAI22_X1 U1843 ( .A1(n3534), .A2(n1308), .B1(n1205), .B2(n1277), .ZN(n6641)
         );
  OAI22_X1 U1847 ( .A1(n3803), .A2(n1311), .B1(n1147), .B2(n1312), .ZN(n6642)
         );
  OAI22_X1 U1849 ( .A1(n3803), .A2(n1313), .B1(n1150), .B2(n1312), .ZN(n6643)
         );
  OAI22_X1 U1851 ( .A1(n3804), .A2(n1314), .B1(n1152), .B2(n1312), .ZN(n6644)
         );
  OAI22_X1 U1853 ( .A1(n3804), .A2(n1315), .B1(n1154), .B2(n1312), .ZN(n6645)
         );
  OAI22_X1 U1855 ( .A1(n3803), .A2(n1316), .B1(n1156), .B2(n1312), .ZN(n6646)
         );
  OAI22_X1 U1857 ( .A1(n3803), .A2(n1317), .B1(n1158), .B2(n1312), .ZN(n6647)
         );
  OAI22_X1 U1859 ( .A1(n3804), .A2(n1318), .B1(n1160), .B2(n1312), .ZN(n6648)
         );
  OAI22_X1 U1861 ( .A1(n3803), .A2(n1319), .B1(n1162), .B2(n1312), .ZN(n6649)
         );
  OAI22_X1 U1863 ( .A1(n3804), .A2(n1320), .B1(n1164), .B2(n1312), .ZN(n6650)
         );
  OAI22_X1 U1865 ( .A1(n3804), .A2(n1321), .B1(n1166), .B2(n1312), .ZN(n6651)
         );
  OAI22_X1 U1867 ( .A1(n3804), .A2(n1322), .B1(n1168), .B2(n1312), .ZN(n6652)
         );
  OAI22_X1 U1869 ( .A1(n3804), .A2(n1323), .B1(n1170), .B2(n1312), .ZN(n6653)
         );
  OAI22_X1 U1871 ( .A1(n3803), .A2(n1324), .B1(n1172), .B2(n1312), .ZN(n6654)
         );
  INV_X1 U1873 ( .A(n1325), .ZN(n6655) );
  AOI22_X1 U1874 ( .A1(n1312), .A2(\pc_lut[27][4] ), .B1(n3521), .B2(n3804), 
        .ZN(n1325) );
  INV_X1 U1876 ( .A(n1326), .ZN(n6657) );
  AOI22_X1 U1877 ( .A1(n1312), .A2(\pc_lut[27][0] ), .B1(n3521), .B2(n3802), 
        .ZN(n1326) );
  INV_X1 U1878 ( .A(n1327), .ZN(n6658) );
  AOI22_X1 U1879 ( .A1(n1312), .A2(\pc_lut[27][1] ), .B1(n3521), .B2(n3802), 
        .ZN(n1327) );
  INV_X1 U1880 ( .A(n1328), .ZN(n6659) );
  AOI22_X1 U1881 ( .A1(n1312), .A2(\pc_lut[27][3] ), .B1(n3521), .B2(n3802), 
        .ZN(n1328) );
  OAI22_X1 U1882 ( .A1(n3803), .A2(n1329), .B1(n1179), .B2(n1312), .ZN(n6660)
         );
  OAI22_X1 U1884 ( .A1(n3803), .A2(n1330), .B1(n1181), .B2(n1312), .ZN(n6661)
         );
  OAI22_X1 U1886 ( .A1(n3804), .A2(n1331), .B1(n1183), .B2(n1312), .ZN(n6662)
         );
  OAI22_X1 U1888 ( .A1(n3803), .A2(n1332), .B1(n1185), .B2(n1312), .ZN(n6663)
         );
  OAI22_X1 U1890 ( .A1(n3804), .A2(n1333), .B1(n1187), .B2(n1312), .ZN(n6664)
         );
  OAI22_X1 U1892 ( .A1(n3803), .A2(n1334), .B1(n1189), .B2(n1312), .ZN(n6665)
         );
  OAI22_X1 U1894 ( .A1(n3804), .A2(n1335), .B1(n1191), .B2(n1312), .ZN(n6666)
         );
  OAI22_X1 U1896 ( .A1(n3803), .A2(n1336), .B1(n1193), .B2(n1312), .ZN(n6667)
         );
  OAI22_X1 U1898 ( .A1(n3804), .A2(n1337), .B1(n1195), .B2(n1312), .ZN(n6668)
         );
  OAI22_X1 U1900 ( .A1(n3803), .A2(n1338), .B1(n1197), .B2(n1312), .ZN(n6669)
         );
  OAI22_X1 U1902 ( .A1(n3804), .A2(n1339), .B1(n1199), .B2(n1312), .ZN(n6670)
         );
  OAI22_X1 U1904 ( .A1(n3803), .A2(n1340), .B1(n1201), .B2(n1312), .ZN(n6671)
         );
  OAI22_X1 U1906 ( .A1(n3804), .A2(n1341), .B1(n1203), .B2(n1312), .ZN(n6672)
         );
  OAI22_X1 U1908 ( .A1(n3803), .A2(n1342), .B1(n1205), .B2(n1312), .ZN(n6673)
         );
  OAI22_X1 U1912 ( .A1(n3538), .A2(n1345), .B1(n1147), .B2(n1346), .ZN(n6674)
         );
  OAI22_X1 U1914 ( .A1(n3538), .A2(n1347), .B1(n1150), .B2(n1346), .ZN(n6675)
         );
  OAI22_X1 U1916 ( .A1(n3538), .A2(n1348), .B1(n1152), .B2(n1346), .ZN(n6676)
         );
  OAI22_X1 U1918 ( .A1(n3538), .A2(n1349), .B1(n1154), .B2(n1346), .ZN(n6677)
         );
  OAI22_X1 U1920 ( .A1(n3538), .A2(n1350), .B1(n1156), .B2(n1346), .ZN(n6678)
         );
  OAI22_X1 U1922 ( .A1(n3538), .A2(n1351), .B1(n1158), .B2(n1346), .ZN(n6679)
         );
  OAI22_X1 U1924 ( .A1(n3538), .A2(n1352), .B1(n1160), .B2(n1346), .ZN(n6680)
         );
  OAI22_X1 U1926 ( .A1(n3538), .A2(n1353), .B1(n1162), .B2(n1346), .ZN(n6681)
         );
  OAI22_X1 U1928 ( .A1(n3538), .A2(n1354), .B1(n1164), .B2(n1346), .ZN(n6682)
         );
  OAI22_X1 U1930 ( .A1(n3538), .A2(n1355), .B1(n1166), .B2(n1346), .ZN(n6683)
         );
  OAI22_X1 U1932 ( .A1(n3538), .A2(n1356), .B1(n1168), .B2(n1346), .ZN(n6684)
         );
  OAI22_X1 U1934 ( .A1(n3538), .A2(n1357), .B1(n1170), .B2(n1346), .ZN(n6685)
         );
  OAI22_X1 U1936 ( .A1(n3538), .A2(n1358), .B1(n1172), .B2(n1346), .ZN(n6686)
         );
  INV_X1 U1938 ( .A(n1359), .ZN(n6687) );
  AOI22_X1 U1939 ( .A1(n1346), .A2(\pc_lut[26][4] ), .B1(n3521), .B2(n3538), 
        .ZN(n1359) );
  INV_X1 U1942 ( .A(n1360), .ZN(n6690) );
  AOI22_X1 U1943 ( .A1(n1346), .A2(\pc_lut[26][1] ), .B1(n3521), .B2(n3538), 
        .ZN(n1360) );
  INV_X1 U1944 ( .A(n1361), .ZN(n6691) );
  AOI22_X1 U1945 ( .A1(n1346), .A2(\pc_lut[26][3] ), .B1(n3521), .B2(n3538), 
        .ZN(n1361) );
  OAI22_X1 U1946 ( .A1(n3538), .A2(n1362), .B1(n1179), .B2(n1346), .ZN(n6692)
         );
  OAI22_X1 U1948 ( .A1(n3538), .A2(n1363), .B1(n1181), .B2(n1346), .ZN(n6693)
         );
  OAI22_X1 U1950 ( .A1(n3538), .A2(n1364), .B1(n1183), .B2(n1346), .ZN(n6694)
         );
  OAI22_X1 U1952 ( .A1(n3538), .A2(n1365), .B1(n1185), .B2(n1346), .ZN(n6695)
         );
  OAI22_X1 U1954 ( .A1(n3538), .A2(n1366), .B1(n1187), .B2(n1346), .ZN(n6696)
         );
  OAI22_X1 U1956 ( .A1(n3538), .A2(n1367), .B1(n1189), .B2(n1346), .ZN(n6697)
         );
  OAI22_X1 U1958 ( .A1(n3538), .A2(n1368), .B1(n1191), .B2(n1346), .ZN(n6698)
         );
  OAI22_X1 U1960 ( .A1(n3538), .A2(n1369), .B1(n1193), .B2(n1346), .ZN(n6699)
         );
  OAI22_X1 U1962 ( .A1(n3538), .A2(n1370), .B1(n1195), .B2(n1346), .ZN(n6700)
         );
  OAI22_X1 U1964 ( .A1(n3538), .A2(n1371), .B1(n1197), .B2(n1346), .ZN(n6701)
         );
  OAI22_X1 U1966 ( .A1(n3538), .A2(n1372), .B1(n1199), .B2(n1346), .ZN(n6702)
         );
  OAI22_X1 U1968 ( .A1(n3538), .A2(n1373), .B1(n1201), .B2(n1346), .ZN(n6703)
         );
  OAI22_X1 U1970 ( .A1(n3538), .A2(n1374), .B1(n1203), .B2(n1346), .ZN(n6704)
         );
  OAI22_X1 U1972 ( .A1(n3538), .A2(n1375), .B1(n1205), .B2(n1346), .ZN(n6705)
         );
  OAI22_X1 U1976 ( .A1(n1376), .A2(n1377), .B1(n1147), .B2(n1378), .ZN(n6706)
         );
  OAI22_X1 U1977 ( .A1(n1376), .A2(n1379), .B1(n1150), .B2(n1378), .ZN(n6707)
         );
  OAI22_X1 U1978 ( .A1(n1376), .A2(n1380), .B1(n1152), .B2(n1378), .ZN(n6708)
         );
  OAI22_X1 U1979 ( .A1(n1376), .A2(n1381), .B1(n1154), .B2(n1378), .ZN(n6709)
         );
  OAI22_X1 U1980 ( .A1(n1376), .A2(n1382), .B1(n1156), .B2(n1378), .ZN(n6710)
         );
  OAI22_X1 U1981 ( .A1(n1376), .A2(n1383), .B1(n1158), .B2(n1378), .ZN(n6711)
         );
  OAI22_X1 U1982 ( .A1(n1376), .A2(n1384), .B1(n1160), .B2(n1378), .ZN(n6712)
         );
  OAI22_X1 U1983 ( .A1(n1376), .A2(n1385), .B1(n1162), .B2(n1378), .ZN(n6713)
         );
  OAI22_X1 U1984 ( .A1(n1376), .A2(n1386), .B1(n1164), .B2(n1378), .ZN(n6714)
         );
  OAI22_X1 U1985 ( .A1(n1376), .A2(n1387), .B1(n1166), .B2(n1378), .ZN(n6715)
         );
  OAI22_X1 U1986 ( .A1(n1376), .A2(n1388), .B1(n1168), .B2(n1378), .ZN(n6716)
         );
  OAI22_X1 U1987 ( .A1(n1376), .A2(n1389), .B1(n1170), .B2(n1378), .ZN(n6717)
         );
  OAI22_X1 U1988 ( .A1(n1376), .A2(n1390), .B1(n1172), .B2(n1378), .ZN(n6718)
         );
  OAI22_X1 U1989 ( .A1(n1376), .A2(n1391), .B1(n3529), .B2(n1378), .ZN(n6719)
         );
  OAI22_X1 U1991 ( .A1(n1376), .A2(n1393), .B1(n3529), .B2(n1378), .ZN(n6721)
         );
  OAI22_X1 U1993 ( .A1(n1376), .A2(n1395), .B1(n3529), .B2(n1378), .ZN(n6723)
         );
  OAI22_X1 U1994 ( .A1(n1376), .A2(n1396), .B1(n1179), .B2(n1378), .ZN(n6724)
         );
  OAI22_X1 U1995 ( .A1(n1376), .A2(n1397), .B1(n1181), .B2(n1378), .ZN(n6725)
         );
  OAI22_X1 U1996 ( .A1(n1376), .A2(n1398), .B1(n1183), .B2(n1378), .ZN(n6726)
         );
  OAI22_X1 U1997 ( .A1(n1376), .A2(n1399), .B1(n1185), .B2(n1378), .ZN(n6727)
         );
  OAI22_X1 U1998 ( .A1(n1376), .A2(n1400), .B1(n1187), .B2(n1378), .ZN(n6728)
         );
  OAI22_X1 U1999 ( .A1(n1376), .A2(n1401), .B1(n1189), .B2(n1378), .ZN(n6729)
         );
  OAI22_X1 U2000 ( .A1(n1376), .A2(n1402), .B1(n1191), .B2(n1378), .ZN(n6730)
         );
  OAI22_X1 U2001 ( .A1(n1376), .A2(n1403), .B1(n1193), .B2(n1378), .ZN(n6731)
         );
  OAI22_X1 U2002 ( .A1(n1376), .A2(n1404), .B1(n1195), .B2(n1378), .ZN(n6732)
         );
  OAI22_X1 U2003 ( .A1(n1376), .A2(n1405), .B1(n1197), .B2(n1378), .ZN(n6733)
         );
  OAI22_X1 U2004 ( .A1(n1376), .A2(n1406), .B1(n1199), .B2(n1378), .ZN(n6734)
         );
  OAI22_X1 U2005 ( .A1(n1376), .A2(n1407), .B1(n1201), .B2(n1378), .ZN(n6735)
         );
  OAI22_X1 U2006 ( .A1(n1376), .A2(n1408), .B1(n1203), .B2(n1378), .ZN(n6736)
         );
  OAI22_X1 U2007 ( .A1(n1376), .A2(n1409), .B1(n1205), .B2(n1378), .ZN(n6737)
         );
  OAI22_X1 U2010 ( .A1(n1410), .A2(n1411), .B1(n1147), .B2(n1412), .ZN(n6738)
         );
  OAI22_X1 U2011 ( .A1(n1410), .A2(n1413), .B1(n1150), .B2(n1412), .ZN(n6739)
         );
  OAI22_X1 U2012 ( .A1(n1410), .A2(n1414), .B1(n1152), .B2(n1412), .ZN(n6740)
         );
  OAI22_X1 U2013 ( .A1(n1410), .A2(n1415), .B1(n1154), .B2(n1412), .ZN(n6741)
         );
  OAI22_X1 U2014 ( .A1(n1410), .A2(n1416), .B1(n1156), .B2(n1412), .ZN(n6742)
         );
  OAI22_X1 U2015 ( .A1(n1410), .A2(n1417), .B1(n1158), .B2(n1412), .ZN(n6743)
         );
  OAI22_X1 U2016 ( .A1(n1410), .A2(n1418), .B1(n1160), .B2(n1412), .ZN(n6744)
         );
  OAI22_X1 U2017 ( .A1(n1410), .A2(n1419), .B1(n1162), .B2(n1412), .ZN(n6745)
         );
  OAI22_X1 U2018 ( .A1(n1410), .A2(n1420), .B1(n1164), .B2(n1412), .ZN(n6746)
         );
  OAI22_X1 U2019 ( .A1(n1410), .A2(n1421), .B1(n1166), .B2(n1412), .ZN(n6747)
         );
  OAI22_X1 U2020 ( .A1(n1410), .A2(n1422), .B1(n1168), .B2(n1412), .ZN(n6748)
         );
  OAI22_X1 U2021 ( .A1(n1410), .A2(n1423), .B1(n1170), .B2(n1412), .ZN(n6749)
         );
  OAI22_X1 U2022 ( .A1(n1410), .A2(n1424), .B1(n1172), .B2(n1412), .ZN(n6750)
         );
  OAI22_X1 U2023 ( .A1(n1410), .A2(n1425), .B1(n1496), .B2(n1412), .ZN(n6751)
         );
  OAI22_X1 U2027 ( .A1(n1410), .A2(n1429), .B1(n1496), .B2(n1412), .ZN(n6755)
         );
  OAI22_X1 U2028 ( .A1(n1410), .A2(n1430), .B1(n1179), .B2(n1412), .ZN(n6756)
         );
  OAI22_X1 U2029 ( .A1(n1410), .A2(n1431), .B1(n1181), .B2(n1412), .ZN(n6757)
         );
  OAI22_X1 U2030 ( .A1(n1410), .A2(n1432), .B1(n1183), .B2(n1412), .ZN(n6758)
         );
  OAI22_X1 U2031 ( .A1(n1410), .A2(n1433), .B1(n1185), .B2(n1412), .ZN(n6759)
         );
  OAI22_X1 U2032 ( .A1(n1410), .A2(n1434), .B1(n1187), .B2(n1412), .ZN(n6760)
         );
  OAI22_X1 U2033 ( .A1(n1410), .A2(n1435), .B1(n1189), .B2(n1412), .ZN(n6761)
         );
  OAI22_X1 U2034 ( .A1(n1410), .A2(n1436), .B1(n1191), .B2(n1412), .ZN(n6762)
         );
  OAI22_X1 U2035 ( .A1(n1410), .A2(n1437), .B1(n1193), .B2(n1412), .ZN(n6763)
         );
  OAI22_X1 U2036 ( .A1(n1410), .A2(n1438), .B1(n1195), .B2(n1412), .ZN(n6764)
         );
  OAI22_X1 U2037 ( .A1(n1410), .A2(n1439), .B1(n1197), .B2(n1412), .ZN(n6765)
         );
  OAI22_X1 U2038 ( .A1(n1410), .A2(n1440), .B1(n1199), .B2(n1412), .ZN(n6766)
         );
  OAI22_X1 U2039 ( .A1(n1410), .A2(n1441), .B1(n1201), .B2(n1412), .ZN(n6767)
         );
  OAI22_X1 U2040 ( .A1(n1410), .A2(n1442), .B1(n1203), .B2(n1412), .ZN(n6768)
         );
  OAI22_X1 U2041 ( .A1(n1410), .A2(n1443), .B1(n1205), .B2(n1412), .ZN(n6769)
         );
  OAI22_X1 U2045 ( .A1(n1444), .A2(n1445), .B1(n1147), .B2(n1427), .ZN(n6770)
         );
  OAI22_X1 U2046 ( .A1(n1444), .A2(n1447), .B1(n1150), .B2(n1428), .ZN(n6771)
         );
  OAI22_X1 U2047 ( .A1(n1444), .A2(n1448), .B1(n1152), .B2(n1428), .ZN(n6772)
         );
  OAI22_X1 U2048 ( .A1(n1444), .A2(n1449), .B1(n1154), .B2(n1428), .ZN(n6773)
         );
  OAI22_X1 U2049 ( .A1(n1444), .A2(n1450), .B1(n1156), .B2(n1428), .ZN(n6774)
         );
  OAI22_X1 U2050 ( .A1(n1444), .A2(n1451), .B1(n1158), .B2(n1427), .ZN(n6775)
         );
  OAI22_X1 U2051 ( .A1(n1444), .A2(n1452), .B1(n1160), .B2(n1428), .ZN(n6776)
         );
  OAI22_X1 U2052 ( .A1(n1444), .A2(n1453), .B1(n1162), .B2(n1427), .ZN(n6777)
         );
  OAI22_X1 U2053 ( .A1(n1444), .A2(n1454), .B1(n1164), .B2(n1428), .ZN(n6778)
         );
  OAI22_X1 U2054 ( .A1(n1444), .A2(n1455), .B1(n1166), .B2(n1427), .ZN(n6779)
         );
  OAI22_X1 U2055 ( .A1(n1444), .A2(n1456), .B1(n1168), .B2(n1428), .ZN(n6780)
         );
  OAI22_X1 U2056 ( .A1(n1444), .A2(n1457), .B1(n1170), .B2(n1428), .ZN(n6781)
         );
  OAI22_X1 U2057 ( .A1(n1444), .A2(n1458), .B1(n1172), .B2(n1428), .ZN(n6782)
         );
  OAI22_X1 U2058 ( .A1(n1444), .A2(n1459), .B1(n3529), .B2(n1428), .ZN(n6783)
         );
  OAI22_X1 U2059 ( .A1(n1444), .A2(n1460), .B1(n3529), .B2(n1428), .ZN(n6784)
         );
  OAI22_X1 U2060 ( .A1(n1444), .A2(n1461), .B1(n3529), .B2(n1428), .ZN(n6785)
         );
  OAI22_X1 U2061 ( .A1(n1444), .A2(n1462), .B1(n3529), .B2(n1428), .ZN(n6786)
         );
  OAI22_X1 U2063 ( .A1(n1444), .A2(n1464), .B1(n1179), .B2(n1428), .ZN(n6788)
         );
  OAI22_X1 U2064 ( .A1(n1444), .A2(n1465), .B1(n1181), .B2(n1428), .ZN(n6789)
         );
  OAI22_X1 U2065 ( .A1(n1444), .A2(n1466), .B1(n1183), .B2(n1428), .ZN(n6790)
         );
  OAI22_X1 U2066 ( .A1(n1444), .A2(n1467), .B1(n1185), .B2(n1428), .ZN(n6791)
         );
  OAI22_X1 U2067 ( .A1(n1444), .A2(n1468), .B1(n1187), .B2(n1428), .ZN(n6792)
         );
  OAI22_X1 U2068 ( .A1(n1444), .A2(n1469), .B1(n1189), .B2(n1428), .ZN(n6793)
         );
  OAI22_X1 U2069 ( .A1(n1444), .A2(n1470), .B1(n1191), .B2(n1428), .ZN(n6794)
         );
  OAI22_X1 U2070 ( .A1(n1444), .A2(n1471), .B1(n1193), .B2(n1428), .ZN(n6795)
         );
  OAI22_X1 U2071 ( .A1(n1444), .A2(n1472), .B1(n1195), .B2(n1427), .ZN(n6796)
         );
  OAI22_X1 U2072 ( .A1(n1444), .A2(n1473), .B1(n1197), .B2(n1428), .ZN(n6797)
         );
  OAI22_X1 U2073 ( .A1(n1444), .A2(n1474), .B1(n1199), .B2(n1428), .ZN(n6798)
         );
  OAI22_X1 U2074 ( .A1(n1444), .A2(n1475), .B1(n1201), .B2(n1428), .ZN(n6799)
         );
  OAI22_X1 U2075 ( .A1(n1444), .A2(n1476), .B1(n1203), .B2(n1428), .ZN(n6800)
         );
  OAI22_X1 U2076 ( .A1(n1444), .A2(n1477), .B1(n1205), .B2(n1428), .ZN(n6801)
         );
  OAI22_X1 U2079 ( .A1(n1479), .A2(n1480), .B1(n1147), .B2(n1394), .ZN(n6802)
         );
  OAI22_X1 U2080 ( .A1(n1479), .A2(n1482), .B1(n1150), .B2(n1394), .ZN(n6803)
         );
  OAI22_X1 U2081 ( .A1(n1479), .A2(n1483), .B1(n1152), .B2(n1392), .ZN(n6804)
         );
  OAI22_X1 U2082 ( .A1(n1479), .A2(n1484), .B1(n1154), .B2(n1394), .ZN(n6805)
         );
  OAI22_X1 U2083 ( .A1(n1479), .A2(n1485), .B1(n1156), .B2(n1394), .ZN(n6806)
         );
  OAI22_X1 U2084 ( .A1(n1479), .A2(n1486), .B1(n1158), .B2(n1392), .ZN(n6807)
         );
  OAI22_X1 U2085 ( .A1(n1479), .A2(n1487), .B1(n1160), .B2(n1394), .ZN(n6808)
         );
  OAI22_X1 U2086 ( .A1(n1479), .A2(n1488), .B1(n1162), .B2(n1392), .ZN(n6809)
         );
  OAI22_X1 U2087 ( .A1(n1479), .A2(n1489), .B1(n1164), .B2(n1394), .ZN(n6810)
         );
  OAI22_X1 U2088 ( .A1(n1479), .A2(n1490), .B1(n1166), .B2(n1394), .ZN(n6811)
         );
  OAI22_X1 U2089 ( .A1(n1479), .A2(n1491), .B1(n1168), .B2(n1394), .ZN(n6812)
         );
  OAI22_X1 U2090 ( .A1(n1479), .A2(n1492), .B1(n1170), .B2(n1394), .ZN(n6813)
         );
  OAI22_X1 U2091 ( .A1(n1479), .A2(n1493), .B1(n1172), .B2(n1394), .ZN(n6814)
         );
  OAI22_X1 U2092 ( .A1(n1479), .A2(n1494), .B1(n3529), .B2(n1394), .ZN(n6815)
         );
  OAI22_X1 U2093 ( .A1(n1479), .A2(n1495), .B1(n3529), .B2(n1394), .ZN(n6816)
         );
  OAI22_X1 U2095 ( .A1(n1479), .A2(n1497), .B1(n3529), .B2(n1392), .ZN(n6818)
         );
  OAI22_X1 U2097 ( .A1(n1479), .A2(n1499), .B1(n1179), .B2(n1394), .ZN(n6820)
         );
  OAI22_X1 U2098 ( .A1(n1479), .A2(n1500), .B1(n1181), .B2(n1394), .ZN(n6821)
         );
  OAI22_X1 U2099 ( .A1(n1479), .A2(n1501), .B1(n1183), .B2(n1394), .ZN(n6822)
         );
  OAI22_X1 U2100 ( .A1(n1479), .A2(n1502), .B1(n1185), .B2(n1394), .ZN(n6823)
         );
  OAI22_X1 U2101 ( .A1(n1479), .A2(n1503), .B1(n1187), .B2(n1394), .ZN(n6824)
         );
  OAI22_X1 U2102 ( .A1(n1479), .A2(n1504), .B1(n1189), .B2(n1394), .ZN(n6825)
         );
  OAI22_X1 U2103 ( .A1(n1479), .A2(n1505), .B1(n1191), .B2(n1394), .ZN(n6826)
         );
  OAI22_X1 U2104 ( .A1(n1479), .A2(n1506), .B1(n1193), .B2(n1394), .ZN(n6827)
         );
  OAI22_X1 U2105 ( .A1(n1479), .A2(n1507), .B1(n1195), .B2(n1394), .ZN(n6828)
         );
  OAI22_X1 U2106 ( .A1(n1479), .A2(n1508), .B1(n1197), .B2(n1394), .ZN(n6829)
         );
  OAI22_X1 U2107 ( .A1(n1479), .A2(n1509), .B1(n1199), .B2(n1394), .ZN(n6830)
         );
  OAI22_X1 U2108 ( .A1(n1479), .A2(n1510), .B1(n1201), .B2(n1394), .ZN(n6831)
         );
  OAI22_X1 U2109 ( .A1(n1479), .A2(n1511), .B1(n1203), .B2(n1394), .ZN(n6832)
         );
  OAI22_X1 U2110 ( .A1(n1479), .A2(n1512), .B1(n1205), .B2(n1394), .ZN(n6833)
         );
  OAI22_X1 U2113 ( .A1(n3810), .A2(n1514), .B1(n1147), .B2(n1515), .ZN(n6834)
         );
  OAI22_X1 U2115 ( .A1(n3810), .A2(n1516), .B1(n1150), .B2(n1515), .ZN(n6835)
         );
  OAI22_X1 U2117 ( .A1(n3810), .A2(n1517), .B1(n1152), .B2(n1515), .ZN(n6836)
         );
  OAI22_X1 U2119 ( .A1(n3810), .A2(n1518), .B1(n1154), .B2(n1515), .ZN(n6837)
         );
  OAI22_X1 U2121 ( .A1(n3810), .A2(n1519), .B1(n1156), .B2(n1515), .ZN(n6838)
         );
  OAI22_X1 U2123 ( .A1(n3810), .A2(n1520), .B1(n1158), .B2(n1515), .ZN(n6839)
         );
  OAI22_X1 U2125 ( .A1(n3810), .A2(n1521), .B1(n1160), .B2(n1515), .ZN(n6840)
         );
  OAI22_X1 U2127 ( .A1(n3810), .A2(n1522), .B1(n1162), .B2(n1515), .ZN(n6841)
         );
  OAI22_X1 U2129 ( .A1(n3810), .A2(n1523), .B1(n1164), .B2(n1515), .ZN(n6842)
         );
  OAI22_X1 U2131 ( .A1(n3810), .A2(n1524), .B1(n1166), .B2(n1515), .ZN(n6843)
         );
  OAI22_X1 U2133 ( .A1(n3810), .A2(n1525), .B1(n1168), .B2(n1515), .ZN(n6844)
         );
  OAI22_X1 U2135 ( .A1(n3810), .A2(n1526), .B1(n1170), .B2(n1515), .ZN(n6845)
         );
  OAI22_X1 U2137 ( .A1(n3810), .A2(n1527), .B1(n1172), .B2(n1515), .ZN(n6846)
         );
  INV_X1 U2139 ( .A(n1528), .ZN(n6847) );
  AOI22_X1 U2140 ( .A1(n1515), .A2(\pc_lut[21][4] ), .B1(n3521), .B2(n3810), 
        .ZN(n1528) );
  INV_X1 U2141 ( .A(n1529), .ZN(n6848) );
  AOI22_X1 U2142 ( .A1(n1515), .A2(\pc_lut[21][2] ), .B1(n3521), .B2(n3810), 
        .ZN(n1529) );
  INV_X1 U2143 ( .A(n1530), .ZN(n6849) );
  AOI22_X1 U2144 ( .A1(n1515), .A2(\pc_lut[21][0] ), .B1(n3521), .B2(n3810), 
        .ZN(n1530) );
  OAI22_X1 U2147 ( .A1(n3810), .A2(n1531), .B1(n1179), .B2(n1515), .ZN(n6852)
         );
  OAI22_X1 U2149 ( .A1(n3810), .A2(n1532), .B1(n1181), .B2(n1515), .ZN(n6853)
         );
  OAI22_X1 U2151 ( .A1(n3810), .A2(n1533), .B1(n1183), .B2(n1515), .ZN(n6854)
         );
  OAI22_X1 U2153 ( .A1(n3810), .A2(n1534), .B1(n1185), .B2(n1515), .ZN(n6855)
         );
  OAI22_X1 U2155 ( .A1(n3810), .A2(n1535), .B1(n1187), .B2(n1515), .ZN(n6856)
         );
  OAI22_X1 U2157 ( .A1(n3810), .A2(n1536), .B1(n1189), .B2(n1515), .ZN(n6857)
         );
  OAI22_X1 U2159 ( .A1(n3810), .A2(n1537), .B1(n1191), .B2(n1515), .ZN(n6858)
         );
  OAI22_X1 U2161 ( .A1(n3810), .A2(n1538), .B1(n1193), .B2(n1515), .ZN(n6859)
         );
  OAI22_X1 U2163 ( .A1(n3810), .A2(n1539), .B1(n1195), .B2(n1515), .ZN(n6860)
         );
  OAI22_X1 U2165 ( .A1(n3810), .A2(n1540), .B1(n1197), .B2(n1515), .ZN(n6861)
         );
  OAI22_X1 U2167 ( .A1(n3810), .A2(n1541), .B1(n1199), .B2(n1515), .ZN(n6862)
         );
  OAI22_X1 U2169 ( .A1(n3810), .A2(n1542), .B1(n1201), .B2(n1515), .ZN(n6863)
         );
  OAI22_X1 U2171 ( .A1(n3810), .A2(n1543), .B1(n1203), .B2(n1515), .ZN(n6864)
         );
  OAI22_X1 U2173 ( .A1(n3810), .A2(n1544), .B1(n1205), .B2(n1515), .ZN(n6865)
         );
  OAI22_X1 U2177 ( .A1(n3800), .A2(n1546), .B1(n1147), .B2(n1547), .ZN(n6866)
         );
  OAI22_X1 U2179 ( .A1(n3800), .A2(n1548), .B1(n1150), .B2(n1547), .ZN(n6867)
         );
  OAI22_X1 U2181 ( .A1(n3800), .A2(n1549), .B1(n1152), .B2(n1547), .ZN(n6868)
         );
  OAI22_X1 U2183 ( .A1(n3800), .A2(n1550), .B1(n1154), .B2(n1547), .ZN(n6869)
         );
  OAI22_X1 U2185 ( .A1(n3800), .A2(n1551), .B1(n1156), .B2(n1547), .ZN(n6870)
         );
  OAI22_X1 U2187 ( .A1(n3800), .A2(n1552), .B1(n1158), .B2(n1547), .ZN(n6871)
         );
  OAI22_X1 U2189 ( .A1(n3800), .A2(n1553), .B1(n1160), .B2(n1547), .ZN(n6872)
         );
  OAI22_X1 U2191 ( .A1(n3800), .A2(n1554), .B1(n1162), .B2(n1547), .ZN(n6873)
         );
  OAI22_X1 U2193 ( .A1(n3800), .A2(n1555), .B1(n1164), .B2(n1547), .ZN(n6874)
         );
  OAI22_X1 U2195 ( .A1(n3800), .A2(n1556), .B1(n1166), .B2(n1547), .ZN(n6875)
         );
  OAI22_X1 U2197 ( .A1(n3800), .A2(n1557), .B1(n1168), .B2(n1547), .ZN(n6876)
         );
  OAI22_X1 U2199 ( .A1(n3800), .A2(n1558), .B1(n1170), .B2(n1547), .ZN(n6877)
         );
  OAI22_X1 U2201 ( .A1(n3800), .A2(n1559), .B1(n1172), .B2(n1547), .ZN(n6878)
         );
  INV_X1 U2203 ( .A(n1560), .ZN(n6879) );
  AOI22_X1 U2204 ( .A1(n1547), .A2(\pc_lut[20][4] ), .B1(n3521), .B2(n3800), 
        .ZN(n1560) );
  INV_X1 U2205 ( .A(n1561), .ZN(n6880) );
  AOI22_X1 U2206 ( .A1(n1547), .A2(\pc_lut[20][2] ), .B1(n3521), .B2(n3800), 
        .ZN(n1561) );
  OAI22_X1 U2210 ( .A1(n3800), .A2(n1562), .B1(n1179), .B2(n1547), .ZN(n6884)
         );
  OAI22_X1 U2212 ( .A1(n3800), .A2(n1563), .B1(n1181), .B2(n1547), .ZN(n6885)
         );
  OAI22_X1 U2214 ( .A1(n3800), .A2(n1564), .B1(n1183), .B2(n1547), .ZN(n6886)
         );
  OAI22_X1 U2216 ( .A1(n3800), .A2(n1565), .B1(n1185), .B2(n1547), .ZN(n6887)
         );
  OAI22_X1 U2218 ( .A1(n3800), .A2(n1566), .B1(n1187), .B2(n1547), .ZN(n6888)
         );
  OAI22_X1 U2220 ( .A1(n3800), .A2(n1567), .B1(n1189), .B2(n1547), .ZN(n6889)
         );
  OAI22_X1 U2222 ( .A1(n3800), .A2(n1568), .B1(n1191), .B2(n1547), .ZN(n6890)
         );
  OAI22_X1 U2224 ( .A1(n3800), .A2(n1569), .B1(n1193), .B2(n1547), .ZN(n6891)
         );
  OAI22_X1 U2226 ( .A1(n3800), .A2(n1570), .B1(n1195), .B2(n1547), .ZN(n6892)
         );
  OAI22_X1 U2228 ( .A1(n3800), .A2(n1571), .B1(n1197), .B2(n1547), .ZN(n6893)
         );
  OAI22_X1 U2230 ( .A1(n3800), .A2(n1572), .B1(n1199), .B2(n1547), .ZN(n6894)
         );
  OAI22_X1 U2232 ( .A1(n3800), .A2(n1573), .B1(n1201), .B2(n1547), .ZN(n6895)
         );
  OAI22_X1 U2234 ( .A1(n3800), .A2(n1574), .B1(n1203), .B2(n1547), .ZN(n6896)
         );
  OAI22_X1 U2236 ( .A1(n3800), .A2(n1575), .B1(n1205), .B2(n1547), .ZN(n6897)
         );
  AND2_X1 U2240 ( .A1(n1309), .A2(n454), .ZN(n1478) );
  OAI22_X1 U2241 ( .A1(n1576), .A2(n1577), .B1(n1147), .B2(n3532), .ZN(n6898)
         );
  OAI22_X1 U2243 ( .A1(n1576), .A2(n1579), .B1(n1150), .B2(n3532), .ZN(n6899)
         );
  OAI22_X1 U2245 ( .A1(n1576), .A2(n1580), .B1(n1152), .B2(n3532), .ZN(n6900)
         );
  OAI22_X1 U2247 ( .A1(n1576), .A2(n1581), .B1(n1154), .B2(n3532), .ZN(n6901)
         );
  OAI22_X1 U2249 ( .A1(n1576), .A2(n1582), .B1(n1156), .B2(n3533), .ZN(n6902)
         );
  OAI22_X1 U2251 ( .A1(n1576), .A2(n1583), .B1(n1158), .B2(n3533), .ZN(n6903)
         );
  OAI22_X1 U2253 ( .A1(n1576), .A2(n1584), .B1(n1160), .B2(n3532), .ZN(n6904)
         );
  OAI22_X1 U2255 ( .A1(n1576), .A2(n1585), .B1(n1162), .B2(n3533), .ZN(n6905)
         );
  OAI22_X1 U2257 ( .A1(n1576), .A2(n1586), .B1(n1164), .B2(n3533), .ZN(n6906)
         );
  OAI22_X1 U2259 ( .A1(n1576), .A2(n1587), .B1(n1166), .B2(n3533), .ZN(n6907)
         );
  OAI22_X1 U2261 ( .A1(n1576), .A2(n1588), .B1(n1168), .B2(n3532), .ZN(n6908)
         );
  OAI22_X1 U2263 ( .A1(n1576), .A2(n1589), .B1(n1170), .B2(n3532), .ZN(n6909)
         );
  OAI22_X1 U2265 ( .A1(n1576), .A2(n1590), .B1(n1172), .B2(n3532), .ZN(n6910)
         );
  INV_X1 U2267 ( .A(n1591), .ZN(n6911) );
  AOI22_X1 U2268 ( .A1(n3533), .A2(\pc_lut[19][4] ), .B1(n3521), .B2(n1576), 
        .ZN(n1591) );
  INV_X1 U2270 ( .A(n1592), .ZN(n6913) );
  AOI22_X1 U2271 ( .A1(n3532), .A2(\pc_lut[19][0] ), .B1(n3521), .B2(n1576), 
        .ZN(n1592) );
  INV_X1 U2272 ( .A(n1593), .ZN(n6914) );
  AOI22_X1 U2273 ( .A1(n3533), .A2(\pc_lut[19][1] ), .B1(n3521), .B2(n1576), 
        .ZN(n1593) );
  OAI22_X1 U2275 ( .A1(n1576), .A2(n1594), .B1(n1179), .B2(n3532), .ZN(n6916)
         );
  OAI22_X1 U2277 ( .A1(n1576), .A2(n1595), .B1(n1181), .B2(n3533), .ZN(n6917)
         );
  OAI22_X1 U2279 ( .A1(n1576), .A2(n1596), .B1(n1183), .B2(n3532), .ZN(n6918)
         );
  OAI22_X1 U2281 ( .A1(n1576), .A2(n1597), .B1(n1185), .B2(n3533), .ZN(n6919)
         );
  OAI22_X1 U2283 ( .A1(n1576), .A2(n1598), .B1(n1187), .B2(n3532), .ZN(n6920)
         );
  OAI22_X1 U2285 ( .A1(n1576), .A2(n1599), .B1(n1189), .B2(n3533), .ZN(n6921)
         );
  OAI22_X1 U2287 ( .A1(n1576), .A2(n1600), .B1(n1191), .B2(n3533), .ZN(n6922)
         );
  OAI22_X1 U2289 ( .A1(n1576), .A2(n1601), .B1(n1193), .B2(n3533), .ZN(n6923)
         );
  OAI22_X1 U2291 ( .A1(n1576), .A2(n1602), .B1(n1195), .B2(n3532), .ZN(n6924)
         );
  OAI22_X1 U2293 ( .A1(n1576), .A2(n1603), .B1(n1197), .B2(n3533), .ZN(n6925)
         );
  OAI22_X1 U2295 ( .A1(n1576), .A2(n1604), .B1(n1199), .B2(n3532), .ZN(n6926)
         );
  OAI22_X1 U2297 ( .A1(n1576), .A2(n1605), .B1(n1201), .B2(n3533), .ZN(n6927)
         );
  OAI22_X1 U2299 ( .A1(n1576), .A2(n1606), .B1(n1203), .B2(n3532), .ZN(n6928)
         );
  OAI22_X1 U2301 ( .A1(n1576), .A2(n1607), .B1(n1205), .B2(n3533), .ZN(n6929)
         );
  NAND2_X1 U2304 ( .A1(n1608), .A2(n38), .ZN(n1578) );
  OAI22_X1 U2305 ( .A1(n1609), .A2(n1610), .B1(n1147), .B2(n558), .ZN(n6930)
         );
  OAI22_X1 U2307 ( .A1(n1609), .A2(n1612), .B1(n1150), .B2(n768), .ZN(n6931)
         );
  OAI22_X1 U2309 ( .A1(n1609), .A2(n1613), .B1(n1152), .B2(n768), .ZN(n6932)
         );
  OAI22_X1 U2311 ( .A1(n1609), .A2(n1614), .B1(n1154), .B2(n768), .ZN(n6933)
         );
  OAI22_X1 U2313 ( .A1(n1609), .A2(n1615), .B1(n1156), .B2(n768), .ZN(n6934)
         );
  OAI22_X1 U2315 ( .A1(n1609), .A2(n1616), .B1(n1158), .B2(n768), .ZN(n6935)
         );
  OAI22_X1 U2317 ( .A1(n1609), .A2(n1617), .B1(n1160), .B2(n768), .ZN(n6936)
         );
  OAI22_X1 U2319 ( .A1(n1609), .A2(n1618), .B1(n1162), .B2(n768), .ZN(n6937)
         );
  OAI22_X1 U2321 ( .A1(n1609), .A2(n1619), .B1(n1164), .B2(n768), .ZN(n6938)
         );
  OAI22_X1 U2323 ( .A1(n1609), .A2(n1620), .B1(n1166), .B2(n768), .ZN(n6939)
         );
  OAI22_X1 U2325 ( .A1(n1609), .A2(n1621), .B1(n1168), .B2(n768), .ZN(n6940)
         );
  OAI22_X1 U2327 ( .A1(n1609), .A2(n1622), .B1(n1170), .B2(n768), .ZN(n6941)
         );
  OAI22_X1 U2329 ( .A1(n1609), .A2(n1623), .B1(n1172), .B2(n768), .ZN(n6942)
         );
  INV_X1 U2331 ( .A(n1624), .ZN(n6943) );
  AOI22_X1 U2332 ( .A1(n558), .A2(\pc_lut[18][4] ), .B1(n3521), .B2(n1609), 
        .ZN(n1624) );
  INV_X1 U2335 ( .A(n1625), .ZN(n6946) );
  AOI22_X1 U2336 ( .A1(n558), .A2(\pc_lut[18][1] ), .B1(n3521), .B2(n1609), 
        .ZN(n1625) );
  OAI22_X1 U2338 ( .A1(n1609), .A2(n1626), .B1(n1179), .B2(n768), .ZN(n6948)
         );
  OAI22_X1 U2340 ( .A1(n1609), .A2(n1627), .B1(n1181), .B2(n768), .ZN(n6949)
         );
  OAI22_X1 U2342 ( .A1(n1609), .A2(n1628), .B1(n1183), .B2(n768), .ZN(n6950)
         );
  OAI22_X1 U2344 ( .A1(n1609), .A2(n1629), .B1(n1185), .B2(n768), .ZN(n6951)
         );
  OAI22_X1 U2346 ( .A1(n1609), .A2(n1630), .B1(n1187), .B2(n768), .ZN(n6952)
         );
  OAI22_X1 U2348 ( .A1(n1609), .A2(n1631), .B1(n1189), .B2(n768), .ZN(n6953)
         );
  OAI22_X1 U2350 ( .A1(n1609), .A2(n1632), .B1(n1191), .B2(n768), .ZN(n6954)
         );
  OAI22_X1 U2352 ( .A1(n1609), .A2(n1633), .B1(n1193), .B2(n768), .ZN(n6955)
         );
  OAI22_X1 U2354 ( .A1(n1609), .A2(n1634), .B1(n1195), .B2(n768), .ZN(n6956)
         );
  OAI22_X1 U2356 ( .A1(n1609), .A2(n1635), .B1(n1197), .B2(n768), .ZN(n6957)
         );
  OAI22_X1 U2358 ( .A1(n1609), .A2(n1636), .B1(n1199), .B2(n768), .ZN(n6958)
         );
  OAI22_X1 U2360 ( .A1(n1609), .A2(n1637), .B1(n1201), .B2(n768), .ZN(n6959)
         );
  OAI22_X1 U2362 ( .A1(n1609), .A2(n1638), .B1(n1203), .B2(n768), .ZN(n6960)
         );
  OAI22_X1 U2364 ( .A1(n1609), .A2(n1639), .B1(n1205), .B2(n768), .ZN(n6961)
         );
  OAI22_X1 U2368 ( .A1(n1640), .A2(n1641), .B1(n1147), .B2(n1642), .ZN(n6962)
         );
  OAI22_X1 U2369 ( .A1(n1640), .A2(n1643), .B1(n1150), .B2(n1642), .ZN(n6963)
         );
  OAI22_X1 U2370 ( .A1(n1640), .A2(n1644), .B1(n1152), .B2(n1642), .ZN(n6964)
         );
  OAI22_X1 U2371 ( .A1(n1640), .A2(n1645), .B1(n1154), .B2(n1642), .ZN(n6965)
         );
  OAI22_X1 U2372 ( .A1(n1640), .A2(n1646), .B1(n1156), .B2(n1642), .ZN(n6966)
         );
  OAI22_X1 U2373 ( .A1(n1640), .A2(n1647), .B1(n1158), .B2(n1642), .ZN(n6967)
         );
  OAI22_X1 U2374 ( .A1(n1640), .A2(n1648), .B1(n1160), .B2(n1642), .ZN(n6968)
         );
  OAI22_X1 U2375 ( .A1(n1640), .A2(n1649), .B1(n1162), .B2(n1642), .ZN(n6969)
         );
  OAI22_X1 U2376 ( .A1(n1640), .A2(n1650), .B1(n1164), .B2(n1642), .ZN(n6970)
         );
  OAI22_X1 U2377 ( .A1(n1640), .A2(n1651), .B1(n1166), .B2(n1642), .ZN(n6971)
         );
  OAI22_X1 U2378 ( .A1(n1640), .A2(n1652), .B1(n1168), .B2(n1642), .ZN(n6972)
         );
  OAI22_X1 U2379 ( .A1(n1640), .A2(n1653), .B1(n1170), .B2(n1642), .ZN(n6973)
         );
  OAI22_X1 U2380 ( .A1(n1640), .A2(n1654), .B1(n1172), .B2(n1642), .ZN(n6974)
         );
  OAI22_X1 U2381 ( .A1(n1640), .A2(n1655), .B1(n1496), .B2(n1642), .ZN(n6975)
         );
  OAI22_X1 U2383 ( .A1(n1640), .A2(n1657), .B1(n1496), .B2(n1642), .ZN(n6977)
         );
  OAI22_X1 U2386 ( .A1(n1640), .A2(n1660), .B1(n1179), .B2(n1642), .ZN(n6980)
         );
  OAI22_X1 U2387 ( .A1(n1640), .A2(n1661), .B1(n1181), .B2(n1642), .ZN(n6981)
         );
  OAI22_X1 U2388 ( .A1(n1640), .A2(n1662), .B1(n1183), .B2(n1642), .ZN(n6982)
         );
  OAI22_X1 U2389 ( .A1(n1640), .A2(n1663), .B1(n1185), .B2(n1642), .ZN(n6983)
         );
  OAI22_X1 U2390 ( .A1(n1640), .A2(n1664), .B1(n1187), .B2(n1642), .ZN(n6984)
         );
  OAI22_X1 U2391 ( .A1(n1640), .A2(n1665), .B1(n1189), .B2(n1642), .ZN(n6985)
         );
  OAI22_X1 U2392 ( .A1(n1640), .A2(n1666), .B1(n1191), .B2(n1642), .ZN(n6986)
         );
  OAI22_X1 U2393 ( .A1(n1640), .A2(n1667), .B1(n1193), .B2(n1642), .ZN(n6987)
         );
  OAI22_X1 U2394 ( .A1(n1640), .A2(n1668), .B1(n1195), .B2(n1642), .ZN(n6988)
         );
  OAI22_X1 U2395 ( .A1(n1640), .A2(n1669), .B1(n1197), .B2(n1642), .ZN(n6989)
         );
  OAI22_X1 U2396 ( .A1(n1640), .A2(n1670), .B1(n1199), .B2(n1642), .ZN(n6990)
         );
  OAI22_X1 U2397 ( .A1(n1640), .A2(n1671), .B1(n1201), .B2(n1642), .ZN(n6991)
         );
  OAI22_X1 U2398 ( .A1(n1640), .A2(n1672), .B1(n1203), .B2(n1642), .ZN(n6992)
         );
  OAI22_X1 U2399 ( .A1(n1640), .A2(n1673), .B1(n1205), .B2(n1642), .ZN(n6993)
         );
  OAI22_X1 U2402 ( .A1(n1674), .A2(n1675), .B1(n1147), .B2(n1676), .ZN(n6994)
         );
  OAI22_X1 U2403 ( .A1(n1674), .A2(n1677), .B1(n1150), .B2(n1676), .ZN(n6995)
         );
  OAI22_X1 U2404 ( .A1(n1674), .A2(n1678), .B1(n1152), .B2(n1676), .ZN(n6996)
         );
  OAI22_X1 U2405 ( .A1(n1674), .A2(n1679), .B1(n1154), .B2(n1676), .ZN(n6997)
         );
  OAI22_X1 U2406 ( .A1(n1674), .A2(n1680), .B1(n1156), .B2(n1676), .ZN(n6998)
         );
  OAI22_X1 U2407 ( .A1(n1674), .A2(n1681), .B1(n1158), .B2(n1676), .ZN(n6999)
         );
  OAI22_X1 U2408 ( .A1(n1674), .A2(n1682), .B1(n1160), .B2(n1676), .ZN(n7000)
         );
  OAI22_X1 U2409 ( .A1(n1674), .A2(n1683), .B1(n1162), .B2(n1676), .ZN(n7001)
         );
  OAI22_X1 U2410 ( .A1(n1674), .A2(n1684), .B1(n1164), .B2(n1676), .ZN(n7002)
         );
  OAI22_X1 U2411 ( .A1(n1674), .A2(n1685), .B1(n1166), .B2(n1676), .ZN(n7003)
         );
  OAI22_X1 U2412 ( .A1(n1674), .A2(n1686), .B1(n1168), .B2(n1676), .ZN(n7004)
         );
  OAI22_X1 U2413 ( .A1(n1674), .A2(n1687), .B1(n1170), .B2(n1676), .ZN(n7005)
         );
  OAI22_X1 U2414 ( .A1(n1674), .A2(n1688), .B1(n1172), .B2(n1676), .ZN(n7006)
         );
  OAI22_X1 U2415 ( .A1(n1674), .A2(n1689), .B1(n1496), .B2(n1676), .ZN(n7007)
         );
  OAI22_X1 U2420 ( .A1(n1674), .A2(n1694), .B1(n1179), .B2(n1676), .ZN(n7012)
         );
  OAI22_X1 U2421 ( .A1(n1674), .A2(n1695), .B1(n1181), .B2(n1676), .ZN(n7013)
         );
  OAI22_X1 U2422 ( .A1(n1674), .A2(n1696), .B1(n1183), .B2(n1676), .ZN(n7014)
         );
  OAI22_X1 U2423 ( .A1(n1674), .A2(n1697), .B1(n1185), .B2(n1676), .ZN(n7015)
         );
  OAI22_X1 U2424 ( .A1(n1674), .A2(n1698), .B1(n1187), .B2(n1676), .ZN(n7016)
         );
  OAI22_X1 U2425 ( .A1(n1674), .A2(n1699), .B1(n1189), .B2(n1676), .ZN(n7017)
         );
  OAI22_X1 U2426 ( .A1(n1674), .A2(n1700), .B1(n1191), .B2(n1676), .ZN(n7018)
         );
  OAI22_X1 U2427 ( .A1(n1674), .A2(n1701), .B1(n1193), .B2(n1676), .ZN(n7019)
         );
  OAI22_X1 U2428 ( .A1(n1674), .A2(n1702), .B1(n1195), .B2(n1676), .ZN(n7020)
         );
  OAI22_X1 U2429 ( .A1(n1674), .A2(n1703), .B1(n1197), .B2(n1676), .ZN(n7021)
         );
  OAI22_X1 U2430 ( .A1(n1674), .A2(n1704), .B1(n1199), .B2(n1676), .ZN(n7022)
         );
  OAI22_X1 U2431 ( .A1(n1674), .A2(n1705), .B1(n1201), .B2(n1676), .ZN(n7023)
         );
  OAI22_X1 U2432 ( .A1(n1674), .A2(n1706), .B1(n1203), .B2(n1676), .ZN(n7024)
         );
  OAI22_X1 U2433 ( .A1(n1674), .A2(n1707), .B1(n1205), .B2(n1676), .ZN(n7025)
         );
  NOR2_X1 U2437 ( .A1(n3793), .A2(n1143), .ZN(n1309) );
  INV_X1 U2438 ( .A(PC_write[4]), .ZN(n1143) );
  OAI22_X1 U2439 ( .A1(n3537), .A2(n1710), .B1(n1147), .B2(n1711), .ZN(n7026)
         );
  OAI22_X1 U2441 ( .A1(n3537), .A2(n1712), .B1(n1150), .B2(n1711), .ZN(n7027)
         );
  OAI22_X1 U2443 ( .A1(n3537), .A2(n1713), .B1(n1152), .B2(n1711), .ZN(n7028)
         );
  OAI22_X1 U2445 ( .A1(n3537), .A2(n1714), .B1(n1154), .B2(n1711), .ZN(n7029)
         );
  OAI22_X1 U2447 ( .A1(n3537), .A2(n1715), .B1(n1156), .B2(n1711), .ZN(n7030)
         );
  OAI22_X1 U2449 ( .A1(n3537), .A2(n1716), .B1(n1158), .B2(n1711), .ZN(n7031)
         );
  OAI22_X1 U2451 ( .A1(n3537), .A2(n1717), .B1(n1160), .B2(n1711), .ZN(n7032)
         );
  OAI22_X1 U2453 ( .A1(n3537), .A2(n1718), .B1(n1162), .B2(n1711), .ZN(n7033)
         );
  OAI22_X1 U2455 ( .A1(n3537), .A2(n1719), .B1(n1164), .B2(n1711), .ZN(n7034)
         );
  OAI22_X1 U2457 ( .A1(n3537), .A2(n1720), .B1(n1166), .B2(n1711), .ZN(n7035)
         );
  OAI22_X1 U2459 ( .A1(n3537), .A2(n1721), .B1(n1168), .B2(n1711), .ZN(n7036)
         );
  OAI22_X1 U2461 ( .A1(n3537), .A2(n1722), .B1(n1170), .B2(n1711), .ZN(n7037)
         );
  OAI22_X1 U2463 ( .A1(n3537), .A2(n1723), .B1(n1172), .B2(n1711), .ZN(n7038)
         );
  INV_X1 U2466 ( .A(n1724), .ZN(n7040) );
  AOI22_X1 U2467 ( .A1(n1711), .A2(\pc_lut[15][2] ), .B1(n3521), .B2(n3537), 
        .ZN(n1724) );
  INV_X1 U2468 ( .A(n1725), .ZN(n7041) );
  AOI22_X1 U2469 ( .A1(n1711), .A2(\pc_lut[15][0] ), .B1(n3521), .B2(n3537), 
        .ZN(n1725) );
  INV_X1 U2470 ( .A(n1726), .ZN(n7042) );
  AOI22_X1 U2471 ( .A1(n1711), .A2(\pc_lut[15][1] ), .B1(n3521), .B2(n3537), 
        .ZN(n1726) );
  INV_X1 U2472 ( .A(n1727), .ZN(n7043) );
  AOI22_X1 U2473 ( .A1(n1711), .A2(\pc_lut[15][3] ), .B1(n3521), .B2(n3537), 
        .ZN(n1727) );
  OAI22_X1 U2474 ( .A1(n3537), .A2(n1728), .B1(n1179), .B2(n1711), .ZN(n7044)
         );
  OAI22_X1 U2476 ( .A1(n3537), .A2(n1729), .B1(n1181), .B2(n1711), .ZN(n7045)
         );
  OAI22_X1 U2478 ( .A1(n3537), .A2(n1730), .B1(n1183), .B2(n1711), .ZN(n7046)
         );
  OAI22_X1 U2480 ( .A1(n3537), .A2(n1731), .B1(n1185), .B2(n1711), .ZN(n7047)
         );
  OAI22_X1 U2482 ( .A1(n3537), .A2(n1732), .B1(n1187), .B2(n1711), .ZN(n7048)
         );
  OAI22_X1 U2484 ( .A1(n3537), .A2(n1733), .B1(n1189), .B2(n1711), .ZN(n7049)
         );
  OAI22_X1 U2486 ( .A1(n3537), .A2(n1734), .B1(n1191), .B2(n1711), .ZN(n7050)
         );
  OAI22_X1 U2488 ( .A1(n3537), .A2(n1735), .B1(n1193), .B2(n1711), .ZN(n7051)
         );
  OAI22_X1 U2490 ( .A1(n3537), .A2(n1736), .B1(n1195), .B2(n1711), .ZN(n7052)
         );
  OAI22_X1 U2492 ( .A1(n3537), .A2(n1737), .B1(n1197), .B2(n1711), .ZN(n7053)
         );
  OAI22_X1 U2494 ( .A1(n3537), .A2(n1738), .B1(n1199), .B2(n1711), .ZN(n7054)
         );
  OAI22_X1 U2496 ( .A1(n3537), .A2(n1739), .B1(n1201), .B2(n1711), .ZN(n7055)
         );
  OAI22_X1 U2498 ( .A1(n3537), .A2(n1740), .B1(n1203), .B2(n1711), .ZN(n7056)
         );
  OAI22_X1 U2500 ( .A1(n3537), .A2(n1741), .B1(n1205), .B2(n1711), .ZN(n7057)
         );
  OAI22_X1 U2504 ( .A1(n3535), .A2(n1744), .B1(n1147), .B2(n1745), .ZN(n7058)
         );
  OAI22_X1 U2506 ( .A1(n3535), .A2(n1746), .B1(n1150), .B2(n1745), .ZN(n7059)
         );
  OAI22_X1 U2508 ( .A1(n3535), .A2(n1747), .B1(n1152), .B2(n1745), .ZN(n7060)
         );
  OAI22_X1 U2510 ( .A1(n3535), .A2(n1748), .B1(n1154), .B2(n1745), .ZN(n7061)
         );
  OAI22_X1 U2512 ( .A1(n3535), .A2(n1749), .B1(n1156), .B2(n1745), .ZN(n7062)
         );
  OAI22_X1 U2514 ( .A1(n3535), .A2(n1750), .B1(n1158), .B2(n1745), .ZN(n7063)
         );
  OAI22_X1 U2516 ( .A1(n3535), .A2(n1751), .B1(n1160), .B2(n1745), .ZN(n7064)
         );
  OAI22_X1 U2518 ( .A1(n3535), .A2(n1752), .B1(n1162), .B2(n1745), .ZN(n7065)
         );
  OAI22_X1 U2520 ( .A1(n3535), .A2(n1753), .B1(n1164), .B2(n1745), .ZN(n7066)
         );
  OAI22_X1 U2522 ( .A1(n3535), .A2(n1754), .B1(n1166), .B2(n1745), .ZN(n7067)
         );
  OAI22_X1 U2524 ( .A1(n3535), .A2(n1755), .B1(n1168), .B2(n1745), .ZN(n7068)
         );
  OAI22_X1 U2526 ( .A1(n3535), .A2(n1756), .B1(n1170), .B2(n1745), .ZN(n7069)
         );
  OAI22_X1 U2528 ( .A1(n3535), .A2(n1757), .B1(n1172), .B2(n1745), .ZN(n7070)
         );
  INV_X1 U2531 ( .A(n1758), .ZN(n7072) );
  AOI22_X1 U2532 ( .A1(n1745), .A2(\pc_lut[14][2] ), .B1(n3521), .B2(n3535), 
        .ZN(n1758) );
  INV_X1 U2534 ( .A(n1759), .ZN(n7074) );
  AOI22_X1 U2535 ( .A1(n1745), .A2(\pc_lut[14][1] ), .B1(n3521), .B2(n3535), 
        .ZN(n1759) );
  INV_X1 U2536 ( .A(n1760), .ZN(n7075) );
  AOI22_X1 U2537 ( .A1(n1745), .A2(\pc_lut[14][3] ), .B1(n3521), .B2(n3535), 
        .ZN(n1760) );
  OAI22_X1 U2538 ( .A1(n3535), .A2(n1761), .B1(n1179), .B2(n1745), .ZN(n7076)
         );
  OAI22_X1 U2540 ( .A1(n3535), .A2(n1762), .B1(n1181), .B2(n1745), .ZN(n7077)
         );
  OAI22_X1 U2542 ( .A1(n3535), .A2(n1763), .B1(n1183), .B2(n1745), .ZN(n7078)
         );
  OAI22_X1 U2544 ( .A1(n3535), .A2(n1764), .B1(n1185), .B2(n1745), .ZN(n7079)
         );
  OAI22_X1 U2546 ( .A1(n3535), .A2(n1765), .B1(n1187), .B2(n1745), .ZN(n7080)
         );
  OAI22_X1 U2548 ( .A1(n3535), .A2(n1766), .B1(n1189), .B2(n1745), .ZN(n7081)
         );
  OAI22_X1 U2550 ( .A1(n3535), .A2(n1767), .B1(n1191), .B2(n1745), .ZN(n7082)
         );
  OAI22_X1 U2552 ( .A1(n3535), .A2(n1768), .B1(n1193), .B2(n1745), .ZN(n7083)
         );
  OAI22_X1 U2554 ( .A1(n3535), .A2(n1769), .B1(n1195), .B2(n1745), .ZN(n7084)
         );
  OAI22_X1 U2556 ( .A1(n3535), .A2(n1770), .B1(n1197), .B2(n1745), .ZN(n7085)
         );
  OAI22_X1 U2558 ( .A1(n3535), .A2(n1771), .B1(n1199), .B2(n1745), .ZN(n7086)
         );
  OAI22_X1 U2560 ( .A1(n3535), .A2(n1772), .B1(n1201), .B2(n1745), .ZN(n7087)
         );
  OAI22_X1 U2562 ( .A1(n3535), .A2(n1773), .B1(n1203), .B2(n1745), .ZN(n7088)
         );
  OAI22_X1 U2564 ( .A1(n3535), .A2(n1774), .B1(n1205), .B2(n1745), .ZN(n7089)
         );
  OAI22_X1 U2568 ( .A1(n1775), .A2(n1776), .B1(n1147), .B2(n1777), .ZN(n7090)
         );
  OAI22_X1 U2569 ( .A1(n1775), .A2(n1778), .B1(n1150), .B2(n1777), .ZN(n7091)
         );
  OAI22_X1 U2570 ( .A1(n1775), .A2(n1779), .B1(n1152), .B2(n1777), .ZN(n7092)
         );
  OAI22_X1 U2571 ( .A1(n1775), .A2(n1780), .B1(n1154), .B2(n1777), .ZN(n7093)
         );
  OAI22_X1 U2572 ( .A1(n1775), .A2(n1781), .B1(n1156), .B2(n1777), .ZN(n7094)
         );
  OAI22_X1 U2573 ( .A1(n1775), .A2(n1782), .B1(n1158), .B2(n1777), .ZN(n7095)
         );
  OAI22_X1 U2574 ( .A1(n1775), .A2(n1783), .B1(n1160), .B2(n1777), .ZN(n7096)
         );
  OAI22_X1 U2575 ( .A1(n1775), .A2(n1784), .B1(n1162), .B2(n1777), .ZN(n7097)
         );
  OAI22_X1 U2576 ( .A1(n1775), .A2(n1785), .B1(n1164), .B2(n1777), .ZN(n7098)
         );
  OAI22_X1 U2577 ( .A1(n1775), .A2(n1786), .B1(n1166), .B2(n1777), .ZN(n7099)
         );
  OAI22_X1 U2578 ( .A1(n1775), .A2(n1787), .B1(n1168), .B2(n1777), .ZN(n7100)
         );
  OAI22_X1 U2579 ( .A1(n1775), .A2(n1788), .B1(n1170), .B2(n1777), .ZN(n7101)
         );
  OAI22_X1 U2580 ( .A1(n1775), .A2(n1789), .B1(n1172), .B2(n1777), .ZN(n7102)
         );
  OAI22_X1 U2582 ( .A1(n1775), .A2(n1791), .B1(n3529), .B2(n1777), .ZN(n7104)
         );
  OAI22_X1 U2583 ( .A1(n1775), .A2(n1792), .B1(n3529), .B2(n1777), .ZN(n7105)
         );
  OAI22_X1 U2585 ( .A1(n1775), .A2(n1794), .B1(n3529), .B2(n1777), .ZN(n7107)
         );
  OAI22_X1 U2586 ( .A1(n1775), .A2(n1795), .B1(n1179), .B2(n1777), .ZN(n7108)
         );
  OAI22_X1 U2587 ( .A1(n1775), .A2(n1796), .B1(n1181), .B2(n1777), .ZN(n7109)
         );
  OAI22_X1 U2588 ( .A1(n1775), .A2(n1797), .B1(n1183), .B2(n1777), .ZN(n7110)
         );
  OAI22_X1 U2589 ( .A1(n1775), .A2(n1798), .B1(n1185), .B2(n1777), .ZN(n7111)
         );
  OAI22_X1 U2590 ( .A1(n1775), .A2(n1799), .B1(n1187), .B2(n1777), .ZN(n7112)
         );
  OAI22_X1 U2591 ( .A1(n1775), .A2(n1800), .B1(n1189), .B2(n1777), .ZN(n7113)
         );
  OAI22_X1 U2592 ( .A1(n1775), .A2(n1801), .B1(n1191), .B2(n1777), .ZN(n7114)
         );
  OAI22_X1 U2593 ( .A1(n1775), .A2(n1802), .B1(n1193), .B2(n1777), .ZN(n7115)
         );
  OAI22_X1 U2594 ( .A1(n1775), .A2(n1803), .B1(n1195), .B2(n1777), .ZN(n7116)
         );
  OAI22_X1 U2595 ( .A1(n1775), .A2(n1804), .B1(n1197), .B2(n1777), .ZN(n7117)
         );
  OAI22_X1 U2596 ( .A1(n1775), .A2(n1805), .B1(n1199), .B2(n1777), .ZN(n7118)
         );
  OAI22_X1 U2597 ( .A1(n1775), .A2(n1806), .B1(n1201), .B2(n1777), .ZN(n7119)
         );
  OAI22_X1 U2598 ( .A1(n1775), .A2(n1807), .B1(n1203), .B2(n1777), .ZN(n7120)
         );
  OAI22_X1 U2599 ( .A1(n1775), .A2(n1808), .B1(n1205), .B2(n1777), .ZN(n7121)
         );
  OAI22_X1 U2602 ( .A1(n1809), .A2(n1810), .B1(n1147), .B2(n1811), .ZN(n7122)
         );
  OAI22_X1 U2603 ( .A1(n1809), .A2(n1812), .B1(n1150), .B2(n1811), .ZN(n7123)
         );
  OAI22_X1 U2604 ( .A1(n1809), .A2(n1813), .B1(n1152), .B2(n1811), .ZN(n7124)
         );
  OAI22_X1 U2605 ( .A1(n1809), .A2(n1814), .B1(n1154), .B2(n1811), .ZN(n7125)
         );
  OAI22_X1 U2606 ( .A1(n1809), .A2(n1815), .B1(n1156), .B2(n1811), .ZN(n7126)
         );
  OAI22_X1 U2607 ( .A1(n1809), .A2(n1816), .B1(n1158), .B2(n1811), .ZN(n7127)
         );
  OAI22_X1 U2608 ( .A1(n1809), .A2(n1817), .B1(n1160), .B2(n1811), .ZN(n7128)
         );
  OAI22_X1 U2609 ( .A1(n1809), .A2(n1818), .B1(n1162), .B2(n1811), .ZN(n7129)
         );
  OAI22_X1 U2610 ( .A1(n1809), .A2(n1819), .B1(n1164), .B2(n1811), .ZN(n7130)
         );
  OAI22_X1 U2611 ( .A1(n1809), .A2(n1820), .B1(n1166), .B2(n1811), .ZN(n7131)
         );
  OAI22_X1 U2612 ( .A1(n1809), .A2(n1821), .B1(n1168), .B2(n1811), .ZN(n7132)
         );
  OAI22_X1 U2613 ( .A1(n1809), .A2(n1822), .B1(n1170), .B2(n1811), .ZN(n7133)
         );
  OAI22_X1 U2614 ( .A1(n1809), .A2(n1823), .B1(n1172), .B2(n1811), .ZN(n7134)
         );
  OAI22_X1 U2616 ( .A1(n1809), .A2(n1825), .B1(n1496), .B2(n1811), .ZN(n7136)
         );
  OAI22_X1 U2619 ( .A1(n1809), .A2(n1828), .B1(n1496), .B2(n1811), .ZN(n7139)
         );
  OAI22_X1 U2620 ( .A1(n1809), .A2(n1829), .B1(n1179), .B2(n1811), .ZN(n7140)
         );
  OAI22_X1 U2621 ( .A1(n1809), .A2(n1830), .B1(n1181), .B2(n1811), .ZN(n7141)
         );
  OAI22_X1 U2622 ( .A1(n1809), .A2(n1831), .B1(n1183), .B2(n1811), .ZN(n7142)
         );
  OAI22_X1 U2623 ( .A1(n1809), .A2(n1832), .B1(n1185), .B2(n1811), .ZN(n7143)
         );
  OAI22_X1 U2624 ( .A1(n1809), .A2(n1833), .B1(n1187), .B2(n1811), .ZN(n7144)
         );
  OAI22_X1 U2625 ( .A1(n1809), .A2(n1834), .B1(n1189), .B2(n1811), .ZN(n7145)
         );
  OAI22_X1 U2626 ( .A1(n1809), .A2(n1835), .B1(n1191), .B2(n1811), .ZN(n7146)
         );
  OAI22_X1 U2627 ( .A1(n1809), .A2(n1836), .B1(n1193), .B2(n1811), .ZN(n7147)
         );
  OAI22_X1 U2628 ( .A1(n1809), .A2(n1837), .B1(n1195), .B2(n1811), .ZN(n7148)
         );
  OAI22_X1 U2629 ( .A1(n1809), .A2(n1838), .B1(n1197), .B2(n1811), .ZN(n7149)
         );
  OAI22_X1 U2630 ( .A1(n1809), .A2(n1839), .B1(n1199), .B2(n1811), .ZN(n7150)
         );
  OAI22_X1 U2631 ( .A1(n1809), .A2(n1840), .B1(n1201), .B2(n1811), .ZN(n7151)
         );
  OAI22_X1 U2632 ( .A1(n1809), .A2(n1841), .B1(n1203), .B2(n1811), .ZN(n7152)
         );
  OAI22_X1 U2633 ( .A1(n1809), .A2(n1842), .B1(n1205), .B2(n1811), .ZN(n7153)
         );
  NOR2_X1 U2637 ( .A1(n1844), .A2(n1845), .ZN(n178) );
  OAI22_X1 U2638 ( .A1(n1846), .A2(n1847), .B1(n1147), .B2(n3527), .ZN(n7154)
         );
  OAI22_X1 U2640 ( .A1(n1846), .A2(n1849), .B1(n1150), .B2(n3527), .ZN(n7155)
         );
  OAI22_X1 U2642 ( .A1(n1846), .A2(n1850), .B1(n1152), .B2(n3527), .ZN(n7156)
         );
  OAI22_X1 U2644 ( .A1(n1846), .A2(n1851), .B1(n1154), .B2(n3527), .ZN(n7157)
         );
  OAI22_X1 U2646 ( .A1(n1846), .A2(n1852), .B1(n1156), .B2(n3527), .ZN(n7158)
         );
  OAI22_X1 U2648 ( .A1(n1846), .A2(n1853), .B1(n1158), .B2(n3527), .ZN(n7159)
         );
  OAI22_X1 U2650 ( .A1(n1846), .A2(n1854), .B1(n1160), .B2(n3527), .ZN(n7160)
         );
  OAI22_X1 U2652 ( .A1(n1846), .A2(n1855), .B1(n1162), .B2(n3527), .ZN(n7161)
         );
  OAI22_X1 U2654 ( .A1(n1846), .A2(n1856), .B1(n1164), .B2(n3527), .ZN(n7162)
         );
  OAI22_X1 U2656 ( .A1(n1846), .A2(n1857), .B1(n1166), .B2(n3527), .ZN(n7163)
         );
  OAI22_X1 U2658 ( .A1(n1846), .A2(n1858), .B1(n1168), .B2(n3527), .ZN(n7164)
         );
  OAI22_X1 U2660 ( .A1(n1846), .A2(n1859), .B1(n1170), .B2(n3527), .ZN(n7165)
         );
  OAI22_X1 U2662 ( .A1(n1846), .A2(n1860), .B1(n1172), .B2(n3527), .ZN(n7166)
         );
  INV_X1 U2666 ( .A(n1861), .ZN(n7169) );
  AOI22_X1 U2667 ( .A1(n3527), .A2(\pc_lut[11][0] ), .B1(n3521), .B2(n1846), 
        .ZN(n1861) );
  INV_X1 U2668 ( .A(n1862), .ZN(n7170) );
  AOI22_X1 U2669 ( .A1(n3527), .A2(\pc_lut[11][1] ), .B1(n3521), .B2(n1846), 
        .ZN(n1862) );
  INV_X1 U2670 ( .A(n1863), .ZN(n7171) );
  AOI22_X1 U2671 ( .A1(n3527), .A2(\pc_lut[11][3] ), .B1(n3521), .B2(n1846), 
        .ZN(n1863) );
  OAI22_X1 U2672 ( .A1(n1846), .A2(n1864), .B1(n1179), .B2(n3527), .ZN(n7172)
         );
  OAI22_X1 U2674 ( .A1(n1846), .A2(n1865), .B1(n1181), .B2(n3527), .ZN(n7173)
         );
  OAI22_X1 U2676 ( .A1(n1846), .A2(n1866), .B1(n1183), .B2(n3527), .ZN(n7174)
         );
  OAI22_X1 U2678 ( .A1(n1846), .A2(n1867), .B1(n1185), .B2(n3527), .ZN(n7175)
         );
  OAI22_X1 U2680 ( .A1(n1846), .A2(n1868), .B1(n1187), .B2(n3527), .ZN(n7176)
         );
  OAI22_X1 U2682 ( .A1(n1846), .A2(n1869), .B1(n1189), .B2(n3527), .ZN(n7177)
         );
  OAI22_X1 U2684 ( .A1(n1846), .A2(n1870), .B1(n1191), .B2(n3527), .ZN(n7178)
         );
  OAI22_X1 U2686 ( .A1(n1846), .A2(n1871), .B1(n1193), .B2(n3527), .ZN(n7179)
         );
  OAI22_X1 U2688 ( .A1(n1846), .A2(n1872), .B1(n1195), .B2(n3527), .ZN(n7180)
         );
  OAI22_X1 U2690 ( .A1(n1846), .A2(n1873), .B1(n1197), .B2(n3527), .ZN(n7181)
         );
  OAI22_X1 U2692 ( .A1(n1846), .A2(n1874), .B1(n1199), .B2(n3527), .ZN(n7182)
         );
  OAI22_X1 U2694 ( .A1(n1846), .A2(n1875), .B1(n1201), .B2(n3527), .ZN(n7183)
         );
  OAI22_X1 U2696 ( .A1(n1846), .A2(n1876), .B1(n1203), .B2(n3527), .ZN(n7184)
         );
  OAI22_X1 U2698 ( .A1(n1846), .A2(n1877), .B1(n1205), .B2(n3527), .ZN(n7185)
         );
  NAND2_X1 U2701 ( .A1(n1878), .A2(n38), .ZN(n1848) );
  OAI22_X1 U2702 ( .A1(n1879), .A2(n1880), .B1(n1147), .B2(n1256), .ZN(n7186)
         );
  OAI22_X1 U2704 ( .A1(n1879), .A2(n1882), .B1(n1150), .B2(n1259), .ZN(n7187)
         );
  OAI22_X1 U2706 ( .A1(n1879), .A2(n1883), .B1(n1152), .B2(n1259), .ZN(n7188)
         );
  OAI22_X1 U2708 ( .A1(n1879), .A2(n1884), .B1(n1154), .B2(n1259), .ZN(n7189)
         );
  OAI22_X1 U2710 ( .A1(n1879), .A2(n1885), .B1(n1156), .B2(n1259), .ZN(n7190)
         );
  OAI22_X1 U2712 ( .A1(n1879), .A2(n1886), .B1(n1158), .B2(n1259), .ZN(n7191)
         );
  OAI22_X1 U2714 ( .A1(n1879), .A2(n1887), .B1(n1160), .B2(n1259), .ZN(n7192)
         );
  OAI22_X1 U2716 ( .A1(n1879), .A2(n1888), .B1(n1162), .B2(n1259), .ZN(n7193)
         );
  OAI22_X1 U2718 ( .A1(n1879), .A2(n1889), .B1(n1164), .B2(n1259), .ZN(n7194)
         );
  OAI22_X1 U2720 ( .A1(n1879), .A2(n1890), .B1(n1166), .B2(n1259), .ZN(n7195)
         );
  OAI22_X1 U2722 ( .A1(n1879), .A2(n1891), .B1(n1168), .B2(n1259), .ZN(n7196)
         );
  OAI22_X1 U2724 ( .A1(n1879), .A2(n1892), .B1(n1170), .B2(n1259), .ZN(n7197)
         );
  OAI22_X1 U2726 ( .A1(n1879), .A2(n1893), .B1(n1172), .B2(n1259), .ZN(n7198)
         );
  INV_X1 U2731 ( .A(n1894), .ZN(n7202) );
  AOI22_X1 U2732 ( .A1(n1256), .A2(\pc_lut[10][1] ), .B1(n3521), .B2(n1879), 
        .ZN(n1894) );
  INV_X1 U2733 ( .A(n1895), .ZN(n7203) );
  AOI22_X1 U2734 ( .A1(n1256), .A2(\pc_lut[10][3] ), .B1(n3521), .B2(n1879), 
        .ZN(n1895) );
  OAI22_X1 U2735 ( .A1(n1879), .A2(n1896), .B1(n1179), .B2(n1259), .ZN(n7204)
         );
  OAI22_X1 U2737 ( .A1(n1879), .A2(n1897), .B1(n1181), .B2(n1259), .ZN(n7205)
         );
  OAI22_X1 U2739 ( .A1(n1879), .A2(n1898), .B1(n1183), .B2(n1259), .ZN(n7206)
         );
  OAI22_X1 U2741 ( .A1(n1879), .A2(n1899), .B1(n1185), .B2(n1259), .ZN(n7207)
         );
  OAI22_X1 U2743 ( .A1(n1879), .A2(n1900), .B1(n1187), .B2(n1259), .ZN(n7208)
         );
  OAI22_X1 U2745 ( .A1(n1879), .A2(n1901), .B1(n1189), .B2(n1259), .ZN(n7209)
         );
  OAI22_X1 U2747 ( .A1(n1879), .A2(n1902), .B1(n1191), .B2(n1259), .ZN(n7210)
         );
  OAI22_X1 U2749 ( .A1(n1879), .A2(n1903), .B1(n1193), .B2(n1259), .ZN(n7211)
         );
  OAI22_X1 U2751 ( .A1(n1879), .A2(n1904), .B1(n1195), .B2(n1259), .ZN(n7212)
         );
  OAI22_X1 U2753 ( .A1(n1879), .A2(n1905), .B1(n1197), .B2(n1259), .ZN(n7213)
         );
  OAI22_X1 U2755 ( .A1(n1879), .A2(n1906), .B1(n1199), .B2(n1259), .ZN(n7214)
         );
  OAI22_X1 U2757 ( .A1(n1879), .A2(n1907), .B1(n1201), .B2(n1259), .ZN(n7215)
         );
  OAI22_X1 U2759 ( .A1(n1879), .A2(n1908), .B1(n1203), .B2(n1259), .ZN(n7216)
         );
  OAI22_X1 U2761 ( .A1(n1879), .A2(n1909), .B1(n1205), .B2(n1259), .ZN(n7217)
         );
  OAI22_X1 U2765 ( .A1(n1910), .A2(n1911), .B1(n1147), .B2(n1912), .ZN(n7218)
         );
  OAI22_X1 U2766 ( .A1(n1910), .A2(n1913), .B1(n1150), .B2(n1912), .ZN(n7219)
         );
  OAI22_X1 U2767 ( .A1(n1910), .A2(n1914), .B1(n1152), .B2(n1912), .ZN(n7220)
         );
  OAI22_X1 U2768 ( .A1(n1910), .A2(n1915), .B1(n1154), .B2(n1912), .ZN(n7221)
         );
  OAI22_X1 U2769 ( .A1(n1910), .A2(n1916), .B1(n1156), .B2(n1912), .ZN(n7222)
         );
  OAI22_X1 U2770 ( .A1(n1910), .A2(n1917), .B1(n1158), .B2(n1912), .ZN(n7223)
         );
  OAI22_X1 U2771 ( .A1(n1910), .A2(n1918), .B1(n1160), .B2(n1912), .ZN(n7224)
         );
  OAI22_X1 U2772 ( .A1(n1910), .A2(n1919), .B1(n1162), .B2(n1912), .ZN(n7225)
         );
  OAI22_X1 U2773 ( .A1(n1910), .A2(n1920), .B1(n1164), .B2(n1912), .ZN(n7226)
         );
  OAI22_X1 U2774 ( .A1(n1910), .A2(n1921), .B1(n1166), .B2(n1912), .ZN(n7227)
         );
  OAI22_X1 U2775 ( .A1(n1910), .A2(n1922), .B1(n1168), .B2(n1912), .ZN(n7228)
         );
  OAI22_X1 U2776 ( .A1(n1910), .A2(n1923), .B1(n1170), .B2(n1912), .ZN(n7229)
         );
  OAI22_X1 U2777 ( .A1(n1910), .A2(n1924), .B1(n1172), .B2(n1912), .ZN(n7230)
         );
  OAI22_X1 U2780 ( .A1(n1910), .A2(n1927), .B1(n1496), .B2(n1912), .ZN(n7233)
         );
  OAI22_X1 U2782 ( .A1(n1910), .A2(n1929), .B1(n1496), .B2(n1912), .ZN(n7235)
         );
  OAI22_X1 U2783 ( .A1(n1910), .A2(n1930), .B1(n1179), .B2(n1912), .ZN(n7236)
         );
  OAI22_X1 U2784 ( .A1(n1910), .A2(n1931), .B1(n1181), .B2(n1912), .ZN(n7237)
         );
  OAI22_X1 U2785 ( .A1(n1910), .A2(n1932), .B1(n1183), .B2(n1912), .ZN(n7238)
         );
  OAI22_X1 U2786 ( .A1(n1910), .A2(n1933), .B1(n1185), .B2(n1912), .ZN(n7239)
         );
  OAI22_X1 U2787 ( .A1(n1910), .A2(n1934), .B1(n1187), .B2(n1912), .ZN(n7240)
         );
  OAI22_X1 U2788 ( .A1(n1910), .A2(n1935), .B1(n1189), .B2(n1912), .ZN(n7241)
         );
  OAI22_X1 U2789 ( .A1(n1910), .A2(n1936), .B1(n1191), .B2(n1912), .ZN(n7242)
         );
  OAI22_X1 U2790 ( .A1(n1910), .A2(n1937), .B1(n1193), .B2(n1912), .ZN(n7243)
         );
  OAI22_X1 U2791 ( .A1(n1910), .A2(n1938), .B1(n1195), .B2(n1912), .ZN(n7244)
         );
  OAI22_X1 U2792 ( .A1(n1910), .A2(n1939), .B1(n1197), .B2(n1912), .ZN(n7245)
         );
  OAI22_X1 U2793 ( .A1(n1910), .A2(n1940), .B1(n1199), .B2(n1912), .ZN(n7246)
         );
  OAI22_X1 U2794 ( .A1(n1910), .A2(n1941), .B1(n1201), .B2(n1912), .ZN(n7247)
         );
  OAI22_X1 U2795 ( .A1(n1910), .A2(n1942), .B1(n1203), .B2(n1912), .ZN(n7248)
         );
  OAI22_X1 U2796 ( .A1(n1910), .A2(n1943), .B1(n1205), .B2(n1912), .ZN(n7249)
         );
  OAI22_X1 U2799 ( .A1(n1944), .A2(n1945), .B1(n1147), .B2(n1946), .ZN(n7250)
         );
  OAI22_X1 U2800 ( .A1(n1944), .A2(n1947), .B1(n1150), .B2(n1946), .ZN(n7251)
         );
  OAI22_X1 U2801 ( .A1(n1944), .A2(n1948), .B1(n1152), .B2(n1946), .ZN(n7252)
         );
  OAI22_X1 U2802 ( .A1(n1944), .A2(n1949), .B1(n1154), .B2(n1946), .ZN(n7253)
         );
  OAI22_X1 U2803 ( .A1(n1944), .A2(n1950), .B1(n1156), .B2(n1946), .ZN(n7254)
         );
  OAI22_X1 U2804 ( .A1(n1944), .A2(n1951), .B1(n1158), .B2(n1946), .ZN(n7255)
         );
  OAI22_X1 U2805 ( .A1(n1944), .A2(n1952), .B1(n1160), .B2(n1946), .ZN(n7256)
         );
  OAI22_X1 U2806 ( .A1(n1944), .A2(n1953), .B1(n1162), .B2(n1946), .ZN(n7257)
         );
  OAI22_X1 U2807 ( .A1(n1944), .A2(n1954), .B1(n1164), .B2(n1946), .ZN(n7258)
         );
  OAI22_X1 U2808 ( .A1(n1944), .A2(n1955), .B1(n1166), .B2(n1946), .ZN(n7259)
         );
  OAI22_X1 U2809 ( .A1(n1944), .A2(n1956), .B1(n1168), .B2(n1946), .ZN(n7260)
         );
  OAI22_X1 U2810 ( .A1(n1944), .A2(n1957), .B1(n1170), .B2(n1946), .ZN(n7261)
         );
  OAI22_X1 U2811 ( .A1(n1944), .A2(n1958), .B1(n1172), .B2(n1946), .ZN(n7262)
         );
  OAI22_X1 U2816 ( .A1(n1944), .A2(n1963), .B1(n1496), .B2(n1946), .ZN(n7267)
         );
  OAI22_X1 U2817 ( .A1(n1944), .A2(n1964), .B1(n1179), .B2(n1946), .ZN(n7268)
         );
  OAI22_X1 U2818 ( .A1(n1944), .A2(n1965), .B1(n1181), .B2(n1946), .ZN(n7269)
         );
  OAI22_X1 U2819 ( .A1(n1944), .A2(n1966), .B1(n1183), .B2(n1946), .ZN(n7270)
         );
  OAI22_X1 U2820 ( .A1(n1944), .A2(n1967), .B1(n1185), .B2(n1946), .ZN(n7271)
         );
  OAI22_X1 U2821 ( .A1(n1944), .A2(n1968), .B1(n1187), .B2(n1946), .ZN(n7272)
         );
  OAI22_X1 U2822 ( .A1(n1944), .A2(n1969), .B1(n1189), .B2(n1946), .ZN(n7273)
         );
  OAI22_X1 U2823 ( .A1(n1944), .A2(n1970), .B1(n1191), .B2(n1946), .ZN(n7274)
         );
  OAI22_X1 U2824 ( .A1(n1944), .A2(n1971), .B1(n1193), .B2(n1946), .ZN(n7275)
         );
  OAI22_X1 U2825 ( .A1(n1944), .A2(n1972), .B1(n1195), .B2(n1946), .ZN(n7276)
         );
  OAI22_X1 U2826 ( .A1(n1944), .A2(n1973), .B1(n1197), .B2(n1946), .ZN(n7277)
         );
  OAI22_X1 U2827 ( .A1(n1944), .A2(n1974), .B1(n1199), .B2(n1946), .ZN(n7278)
         );
  OAI22_X1 U2828 ( .A1(n1944), .A2(n1975), .B1(n1201), .B2(n1946), .ZN(n7279)
         );
  OAI22_X1 U2829 ( .A1(n1944), .A2(n1976), .B1(n1203), .B2(n1946), .ZN(n7280)
         );
  OAI22_X1 U2830 ( .A1(n1944), .A2(n1977), .B1(n1205), .B2(n1946), .ZN(n7281)
         );
  AND2_X1 U2833 ( .A1(n3794), .A2(n316), .ZN(n1878) );
  NOR2_X1 U2834 ( .A1(n1844), .A2(PC_write[2]), .ZN(n316) );
  INV_X1 U2835 ( .A(PC_write[3]), .ZN(n1844) );
  OAI22_X1 U2836 ( .A1(n1978), .A2(n1979), .B1(n1147), .B2(n3524), .ZN(n7282)
         );
  OAI22_X1 U2838 ( .A1(n1978), .A2(n1981), .B1(n1150), .B2(n3524), .ZN(n7283)
         );
  OAI22_X1 U2840 ( .A1(n1978), .A2(n1982), .B1(n1152), .B2(n3524), .ZN(n7284)
         );
  OAI22_X1 U2842 ( .A1(n1978), .A2(n1983), .B1(n1154), .B2(n3524), .ZN(n7285)
         );
  OAI22_X1 U2844 ( .A1(n1978), .A2(n1984), .B1(n1156), .B2(n3524), .ZN(n7286)
         );
  OAI22_X1 U2846 ( .A1(n1978), .A2(n1985), .B1(n1158), .B2(n3524), .ZN(n7287)
         );
  OAI22_X1 U2848 ( .A1(n1978), .A2(n1986), .B1(n1160), .B2(n3524), .ZN(n7288)
         );
  OAI22_X1 U2850 ( .A1(n1978), .A2(n1987), .B1(n1162), .B2(n3524), .ZN(n7289)
         );
  OAI22_X1 U2852 ( .A1(n1978), .A2(n1988), .B1(n1164), .B2(n3524), .ZN(n7290)
         );
  OAI22_X1 U2854 ( .A1(n1978), .A2(n1989), .B1(n1166), .B2(n3524), .ZN(n7291)
         );
  OAI22_X1 U2856 ( .A1(n1978), .A2(n1990), .B1(n1168), .B2(n3524), .ZN(n7292)
         );
  OAI22_X1 U2858 ( .A1(n1978), .A2(n1991), .B1(n1170), .B2(n3524), .ZN(n7293)
         );
  OAI22_X1 U2860 ( .A1(n1978), .A2(n1992), .B1(n1172), .B2(n3524), .ZN(n7294)
         );
  INV_X1 U2863 ( .A(n1993), .ZN(n7296) );
  AOI22_X1 U2864 ( .A1(n3524), .A2(\pc_lut[7][2] ), .B1(n3521), .B2(n1978), 
        .ZN(n1993) );
  INV_X1 U2865 ( .A(n1994), .ZN(n7297) );
  AOI22_X1 U2866 ( .A1(n3524), .A2(\pc_lut[7][0] ), .B1(n3521), .B2(n1978), 
        .ZN(n1994) );
  INV_X1 U2867 ( .A(n1995), .ZN(n7298) );
  AOI22_X1 U2868 ( .A1(n3524), .A2(\pc_lut[7][1] ), .B1(n3521), .B2(n1978), 
        .ZN(n1995) );
  OAI22_X1 U2870 ( .A1(n1978), .A2(n1996), .B1(n1179), .B2(n3524), .ZN(n7300)
         );
  OAI22_X1 U2872 ( .A1(n1978), .A2(n1997), .B1(n1181), .B2(n3524), .ZN(n7301)
         );
  OAI22_X1 U2874 ( .A1(n1978), .A2(n1998), .B1(n1183), .B2(n3524), .ZN(n7302)
         );
  OAI22_X1 U2876 ( .A1(n1978), .A2(n1999), .B1(n1185), .B2(n3524), .ZN(n7303)
         );
  OAI22_X1 U2878 ( .A1(n1978), .A2(n2000), .B1(n1187), .B2(n3524), .ZN(n7304)
         );
  OAI22_X1 U2880 ( .A1(n1978), .A2(n2001), .B1(n1189), .B2(n3524), .ZN(n7305)
         );
  OAI22_X1 U2882 ( .A1(n1978), .A2(n2002), .B1(n1191), .B2(n3524), .ZN(n7306)
         );
  OAI22_X1 U2884 ( .A1(n1978), .A2(n2003), .B1(n1193), .B2(n3524), .ZN(n7307)
         );
  OAI22_X1 U2886 ( .A1(n1978), .A2(n2004), .B1(n1195), .B2(n3524), .ZN(n7308)
         );
  OAI22_X1 U2888 ( .A1(n1978), .A2(n2005), .B1(n1197), .B2(n3524), .ZN(n7309)
         );
  OAI22_X1 U2890 ( .A1(n1978), .A2(n2006), .B1(n1199), .B2(n3524), .ZN(n7310)
         );
  OAI22_X1 U2892 ( .A1(n1978), .A2(n2007), .B1(n1201), .B2(n3524), .ZN(n7311)
         );
  OAI22_X1 U2894 ( .A1(n1978), .A2(n2008), .B1(n1203), .B2(n3524), .ZN(n7312)
         );
  OAI22_X1 U2896 ( .A1(n1978), .A2(n2009), .B1(n1205), .B2(n3524), .ZN(n7313)
         );
  NAND2_X1 U2899 ( .A1(n2010), .A2(n38), .ZN(n1980) );
  OAI22_X1 U2900 ( .A1(n2011), .A2(n2012), .B1(n1147), .B2(n1292), .ZN(n7314)
         );
  OAI22_X1 U2902 ( .A1(n2011), .A2(n2014), .B1(n1150), .B2(n1293), .ZN(n7315)
         );
  OAI22_X1 U2904 ( .A1(n2011), .A2(n2015), .B1(n1152), .B2(n1293), .ZN(n7316)
         );
  OAI22_X1 U2906 ( .A1(n2011), .A2(n2016), .B1(n1154), .B2(n1293), .ZN(n7317)
         );
  OAI22_X1 U2908 ( .A1(n2011), .A2(n2017), .B1(n1156), .B2(n1293), .ZN(n7318)
         );
  OAI22_X1 U2910 ( .A1(n2011), .A2(n2018), .B1(n1158), .B2(n1293), .ZN(n7319)
         );
  OAI22_X1 U2912 ( .A1(n2011), .A2(n2019), .B1(n1160), .B2(n1293), .ZN(n7320)
         );
  OAI22_X1 U2914 ( .A1(n2011), .A2(n2020), .B1(n1162), .B2(n1293), .ZN(n7321)
         );
  OAI22_X1 U2916 ( .A1(n2011), .A2(n2021), .B1(n1164), .B2(n1293), .ZN(n7322)
         );
  OAI22_X1 U2918 ( .A1(n2011), .A2(n2022), .B1(n1166), .B2(n1293), .ZN(n7323)
         );
  OAI22_X1 U2920 ( .A1(n2011), .A2(n2023), .B1(n1168), .B2(n1293), .ZN(n7324)
         );
  OAI22_X1 U2922 ( .A1(n2011), .A2(n2024), .B1(n1170), .B2(n1293), .ZN(n7325)
         );
  OAI22_X1 U2924 ( .A1(n2011), .A2(n2025), .B1(n1172), .B2(n1293), .ZN(n7326)
         );
  INV_X1 U2927 ( .A(n2026), .ZN(n7328) );
  AOI22_X1 U2928 ( .A1(n1292), .A2(\pc_lut[6][2] ), .B1(n3521), .B2(n2011), 
        .ZN(n2026) );
  INV_X1 U2930 ( .A(n2027), .ZN(n7330) );
  AOI22_X1 U2931 ( .A1(n1292), .A2(\pc_lut[6][1] ), .B1(n3521), .B2(n2011), 
        .ZN(n2027) );
  OAI22_X1 U2933 ( .A1(n2011), .A2(n2028), .B1(n1179), .B2(n1293), .ZN(n7332)
         );
  OAI22_X1 U2935 ( .A1(n2011), .A2(n2029), .B1(n1181), .B2(n1293), .ZN(n7333)
         );
  OAI22_X1 U2937 ( .A1(n2011), .A2(n2030), .B1(n1183), .B2(n1293), .ZN(n7334)
         );
  OAI22_X1 U2939 ( .A1(n2011), .A2(n2031), .B1(n1185), .B2(n1293), .ZN(n7335)
         );
  OAI22_X1 U2941 ( .A1(n2011), .A2(n2032), .B1(n1187), .B2(n1293), .ZN(n7336)
         );
  OAI22_X1 U2943 ( .A1(n2011), .A2(n2033), .B1(n1189), .B2(n1293), .ZN(n7337)
         );
  OAI22_X1 U2945 ( .A1(n2011), .A2(n2034), .B1(n1191), .B2(n1293), .ZN(n7338)
         );
  OAI22_X1 U2947 ( .A1(n2011), .A2(n2035), .B1(n1193), .B2(n1293), .ZN(n7339)
         );
  OAI22_X1 U2949 ( .A1(n2011), .A2(n2036), .B1(n1195), .B2(n1293), .ZN(n7340)
         );
  OAI22_X1 U2951 ( .A1(n2011), .A2(n2037), .B1(n1197), .B2(n1293), .ZN(n7341)
         );
  OAI22_X1 U2953 ( .A1(n2011), .A2(n2038), .B1(n1199), .B2(n1293), .ZN(n7342)
         );
  OAI22_X1 U2955 ( .A1(n2011), .A2(n2039), .B1(n1201), .B2(n1293), .ZN(n7343)
         );
  OAI22_X1 U2957 ( .A1(n2011), .A2(n2040), .B1(n1203), .B2(n1293), .ZN(n7344)
         );
  OAI22_X1 U2959 ( .A1(n2011), .A2(n2041), .B1(n1205), .B2(n1293), .ZN(n7345)
         );
  OAI22_X1 U2963 ( .A1(n2042), .A2(n2043), .B1(n1147), .B2(n2044), .ZN(n7346)
         );
  OAI22_X1 U2964 ( .A1(n2042), .A2(n2045), .B1(n1150), .B2(n2044), .ZN(n7347)
         );
  OAI22_X1 U2965 ( .A1(n2042), .A2(n2046), .B1(n1152), .B2(n2044), .ZN(n7348)
         );
  OAI22_X1 U2966 ( .A1(n2042), .A2(n2047), .B1(n1154), .B2(n2044), .ZN(n7349)
         );
  OAI22_X1 U2967 ( .A1(n2042), .A2(n2048), .B1(n1156), .B2(n2044), .ZN(n7350)
         );
  OAI22_X1 U2968 ( .A1(n2042), .A2(n2049), .B1(n1158), .B2(n2044), .ZN(n7351)
         );
  OAI22_X1 U2969 ( .A1(n2042), .A2(n2050), .B1(n1160), .B2(n2044), .ZN(n7352)
         );
  OAI22_X1 U2970 ( .A1(n2042), .A2(n2051), .B1(n1162), .B2(n2044), .ZN(n7353)
         );
  OAI22_X1 U2971 ( .A1(n2042), .A2(n2052), .B1(n1164), .B2(n2044), .ZN(n7354)
         );
  OAI22_X1 U2972 ( .A1(n2042), .A2(n2053), .B1(n1166), .B2(n2044), .ZN(n7355)
         );
  OAI22_X1 U2973 ( .A1(n2042), .A2(n2054), .B1(n1168), .B2(n2044), .ZN(n7356)
         );
  OAI22_X1 U2974 ( .A1(n2042), .A2(n2055), .B1(n1170), .B2(n2044), .ZN(n7357)
         );
  OAI22_X1 U2975 ( .A1(n2042), .A2(n2056), .B1(n1172), .B2(n2044), .ZN(n7358)
         );
  OAI22_X1 U2977 ( .A1(n2042), .A2(n2058), .B1(n1496), .B2(n2044), .ZN(n7360)
         );
  OAI22_X1 U2978 ( .A1(n2042), .A2(n2059), .B1(n1496), .B2(n2044), .ZN(n7361)
         );
  OAI22_X1 U2981 ( .A1(n2042), .A2(n2062), .B1(n1179), .B2(n2044), .ZN(n7364)
         );
  OAI22_X1 U2982 ( .A1(n2042), .A2(n2063), .B1(n1181), .B2(n2044), .ZN(n7365)
         );
  OAI22_X1 U2983 ( .A1(n2042), .A2(n2064), .B1(n1183), .B2(n2044), .ZN(n7366)
         );
  OAI22_X1 U2984 ( .A1(n2042), .A2(n2065), .B1(n1185), .B2(n2044), .ZN(n7367)
         );
  OAI22_X1 U2985 ( .A1(n2042), .A2(n2066), .B1(n1187), .B2(n2044), .ZN(n7368)
         );
  OAI22_X1 U2986 ( .A1(n2042), .A2(n2067), .B1(n1189), .B2(n2044), .ZN(n7369)
         );
  OAI22_X1 U2987 ( .A1(n2042), .A2(n2068), .B1(n1191), .B2(n2044), .ZN(n7370)
         );
  OAI22_X1 U2988 ( .A1(n2042), .A2(n2069), .B1(n1193), .B2(n2044), .ZN(n7371)
         );
  OAI22_X1 U2989 ( .A1(n2042), .A2(n2070), .B1(n1195), .B2(n2044), .ZN(n7372)
         );
  OAI22_X1 U2990 ( .A1(n2042), .A2(n2071), .B1(n1197), .B2(n2044), .ZN(n7373)
         );
  OAI22_X1 U2991 ( .A1(n2042), .A2(n2072), .B1(n1199), .B2(n2044), .ZN(n7374)
         );
  OAI22_X1 U2992 ( .A1(n2042), .A2(n2073), .B1(n1201), .B2(n2044), .ZN(n7375)
         );
  OAI22_X1 U2993 ( .A1(n2042), .A2(n2074), .B1(n1203), .B2(n2044), .ZN(n7376)
         );
  OAI22_X1 U2994 ( .A1(n2042), .A2(n2075), .B1(n1205), .B2(n2044), .ZN(n7377)
         );
  OAI22_X1 U2997 ( .A1(n2076), .A2(n2077), .B1(n1147), .B2(n2078), .ZN(n7378)
         );
  OAI22_X1 U2998 ( .A1(n2076), .A2(n2079), .B1(n1150), .B2(n2078), .ZN(n7379)
         );
  OAI22_X1 U2999 ( .A1(n2076), .A2(n2080), .B1(n1152), .B2(n2078), .ZN(n7380)
         );
  OAI22_X1 U3000 ( .A1(n2076), .A2(n2081), .B1(n1154), .B2(n2078), .ZN(n7381)
         );
  OAI22_X1 U3001 ( .A1(n2076), .A2(n2082), .B1(n1156), .B2(n2078), .ZN(n7382)
         );
  OAI22_X1 U3002 ( .A1(n2076), .A2(n2083), .B1(n1158), .B2(n2078), .ZN(n7383)
         );
  OAI22_X1 U3003 ( .A1(n2076), .A2(n2084), .B1(n1160), .B2(n2078), .ZN(n7384)
         );
  OAI22_X1 U3004 ( .A1(n2076), .A2(n2085), .B1(n1162), .B2(n2078), .ZN(n7385)
         );
  OAI22_X1 U3005 ( .A1(n2076), .A2(n2086), .B1(n1164), .B2(n2078), .ZN(n7386)
         );
  OAI22_X1 U3006 ( .A1(n2076), .A2(n2087), .B1(n1166), .B2(n2078), .ZN(n7387)
         );
  OAI22_X1 U3007 ( .A1(n2076), .A2(n2088), .B1(n1168), .B2(n2078), .ZN(n7388)
         );
  OAI22_X1 U3008 ( .A1(n2076), .A2(n2089), .B1(n1170), .B2(n2078), .ZN(n7389)
         );
  OAI22_X1 U3009 ( .A1(n2076), .A2(n2090), .B1(n1172), .B2(n2078), .ZN(n7390)
         );
  OAI22_X1 U3011 ( .A1(n2076), .A2(n2092), .B1(n1496), .B2(n2078), .ZN(n7392)
         );
  OAI22_X1 U3015 ( .A1(n2076), .A2(n2096), .B1(n1179), .B2(n2078), .ZN(n7396)
         );
  OAI22_X1 U3016 ( .A1(n2076), .A2(n2097), .B1(n1181), .B2(n2078), .ZN(n7397)
         );
  OAI22_X1 U3017 ( .A1(n2076), .A2(n2098), .B1(n1183), .B2(n2078), .ZN(n7398)
         );
  OAI22_X1 U3018 ( .A1(n2076), .A2(n2099), .B1(n1185), .B2(n2078), .ZN(n7399)
         );
  OAI22_X1 U3019 ( .A1(n2076), .A2(n2100), .B1(n1187), .B2(n2078), .ZN(n7400)
         );
  OAI22_X1 U3020 ( .A1(n2076), .A2(n2101), .B1(n1189), .B2(n2078), .ZN(n7401)
         );
  OAI22_X1 U3021 ( .A1(n2076), .A2(n2102), .B1(n1191), .B2(n2078), .ZN(n7402)
         );
  OAI22_X1 U3022 ( .A1(n2076), .A2(n2103), .B1(n1193), .B2(n2078), .ZN(n7403)
         );
  OAI22_X1 U3023 ( .A1(n2076), .A2(n2104), .B1(n1195), .B2(n2078), .ZN(n7404)
         );
  OAI22_X1 U3024 ( .A1(n2076), .A2(n2105), .B1(n1197), .B2(n2078), .ZN(n7405)
         );
  OAI22_X1 U3025 ( .A1(n2076), .A2(n2106), .B1(n1199), .B2(n2078), .ZN(n7406)
         );
  OAI22_X1 U3026 ( .A1(n2076), .A2(n2107), .B1(n1201), .B2(n2078), .ZN(n7407)
         );
  OAI22_X1 U3027 ( .A1(n2076), .A2(n2108), .B1(n1203), .B2(n2078), .ZN(n7408)
         );
  OAI22_X1 U3028 ( .A1(n2076), .A2(n2109), .B1(n1205), .B2(n2078), .ZN(n7409)
         );
  AND2_X1 U3031 ( .A1(n1843), .A2(n454), .ZN(n2010) );
  NOR2_X1 U3032 ( .A1(n1845), .A2(PC_write[3]), .ZN(n454) );
  INV_X1 U3033 ( .A(PC_write[2]), .ZN(n1845) );
  OAI22_X1 U3034 ( .A1(n2110), .A2(n2111), .B1(n1147), .B2(n871), .ZN(n7410)
         );
  OAI22_X1 U3036 ( .A1(n2110), .A2(n2113), .B1(n1150), .B2(n973), .ZN(n7411)
         );
  OAI22_X1 U3038 ( .A1(n2110), .A2(n2114), .B1(n1152), .B2(n973), .ZN(n7412)
         );
  OAI22_X1 U3040 ( .A1(n2110), .A2(n2115), .B1(n1154), .B2(n973), .ZN(n7413)
         );
  OAI22_X1 U3042 ( .A1(n2110), .A2(n2116), .B1(n1156), .B2(n973), .ZN(n7414)
         );
  OAI22_X1 U3044 ( .A1(n2110), .A2(n2117), .B1(n1158), .B2(n973), .ZN(n7415)
         );
  OAI22_X1 U3046 ( .A1(n2110), .A2(n2118), .B1(n1160), .B2(n973), .ZN(n7416)
         );
  OAI22_X1 U3048 ( .A1(n2110), .A2(n2119), .B1(n1162), .B2(n973), .ZN(n7417)
         );
  OAI22_X1 U3050 ( .A1(n2110), .A2(n2120), .B1(n1164), .B2(n973), .ZN(n7418)
         );
  OAI22_X1 U3052 ( .A1(n2110), .A2(n2121), .B1(n1166), .B2(n973), .ZN(n7419)
         );
  OAI22_X1 U3054 ( .A1(n2110), .A2(n2122), .B1(n1168), .B2(n973), .ZN(n7420)
         );
  OAI22_X1 U3056 ( .A1(n2110), .A2(n2123), .B1(n1170), .B2(n973), .ZN(n7421)
         );
  OAI22_X1 U3058 ( .A1(n2110), .A2(n2124), .B1(n1172), .B2(n973), .ZN(n7422)
         );
  INV_X1 U3062 ( .A(n2125), .ZN(n7425) );
  AOI22_X1 U3063 ( .A1(n871), .A2(\pc_lut[3][0] ), .B1(n3521), .B2(n2110), 
        .ZN(n2125) );
  INV_X1 U3064 ( .A(n2126), .ZN(n7426) );
  AOI22_X1 U3065 ( .A1(n871), .A2(\pc_lut[3][1] ), .B1(n3521), .B2(n2110), 
        .ZN(n2126) );
  OAI22_X1 U3067 ( .A1(n2110), .A2(n2127), .B1(n1179), .B2(n973), .ZN(n7428)
         );
  OAI22_X1 U3069 ( .A1(n2110), .A2(n2128), .B1(n1181), .B2(n973), .ZN(n7429)
         );
  OAI22_X1 U3071 ( .A1(n2110), .A2(n2129), .B1(n1183), .B2(n973), .ZN(n7430)
         );
  OAI22_X1 U3073 ( .A1(n2110), .A2(n2130), .B1(n1185), .B2(n973), .ZN(n7431)
         );
  OAI22_X1 U3075 ( .A1(n2110), .A2(n2131), .B1(n1187), .B2(n973), .ZN(n7432)
         );
  OAI22_X1 U3077 ( .A1(n2110), .A2(n2132), .B1(n1189), .B2(n973), .ZN(n7433)
         );
  OAI22_X1 U3079 ( .A1(n2110), .A2(n2133), .B1(n1191), .B2(n973), .ZN(n7434)
         );
  OAI22_X1 U3081 ( .A1(n2110), .A2(n2134), .B1(n1193), .B2(n973), .ZN(n7435)
         );
  OAI22_X1 U3083 ( .A1(n2110), .A2(n2135), .B1(n1195), .B2(n973), .ZN(n7436)
         );
  OAI22_X1 U3085 ( .A1(n2110), .A2(n2136), .B1(n1197), .B2(n973), .ZN(n7437)
         );
  OAI22_X1 U3087 ( .A1(n2110), .A2(n2137), .B1(n1199), .B2(n973), .ZN(n7438)
         );
  OAI22_X1 U3089 ( .A1(n2110), .A2(n2138), .B1(n1201), .B2(n973), .ZN(n7439)
         );
  OAI22_X1 U3091 ( .A1(n2110), .A2(n2139), .B1(n1203), .B2(n973), .ZN(n7440)
         );
  OAI22_X1 U3093 ( .A1(n2110), .A2(n2140), .B1(n1205), .B2(n973), .ZN(n7441)
         );
  OAI22_X1 U3098 ( .A1(n2144), .A2(n2145), .B1(n1147), .B2(n3), .ZN(n7442) );
  OAI22_X1 U3100 ( .A1(n2144), .A2(n2147), .B1(n1150), .B2(n283), .ZN(n7443)
         );
  OAI22_X1 U3102 ( .A1(n2144), .A2(n2148), .B1(n1152), .B2(n283), .ZN(n7444)
         );
  OAI22_X1 U3104 ( .A1(n2144), .A2(n2149), .B1(n1154), .B2(n283), .ZN(n7445)
         );
  OAI22_X1 U3106 ( .A1(n2144), .A2(n2150), .B1(n1156), .B2(n283), .ZN(n7446)
         );
  OAI22_X1 U3108 ( .A1(n2144), .A2(n2151), .B1(n1158), .B2(n283), .ZN(n7447)
         );
  OAI22_X1 U3110 ( .A1(n2144), .A2(n2152), .B1(n1160), .B2(n283), .ZN(n7448)
         );
  OAI22_X1 U3112 ( .A1(n2144), .A2(n2153), .B1(n1162), .B2(n283), .ZN(n7449)
         );
  OAI22_X1 U3114 ( .A1(n2144), .A2(n2154), .B1(n1164), .B2(n283), .ZN(n7450)
         );
  OAI22_X1 U3116 ( .A1(n2144), .A2(n2155), .B1(n1166), .B2(n283), .ZN(n7451)
         );
  OAI22_X1 U3118 ( .A1(n2144), .A2(n2156), .B1(n1168), .B2(n283), .ZN(n7452)
         );
  OAI22_X1 U3120 ( .A1(n2144), .A2(n2157), .B1(n1170), .B2(n283), .ZN(n7453)
         );
  OAI22_X1 U3122 ( .A1(n2144), .A2(n2158), .B1(n1172), .B2(n283), .ZN(n7454)
         );
  INV_X1 U3127 ( .A(n2159), .ZN(n7458) );
  AOI22_X1 U3128 ( .A1(n3), .A2(\pc_lut[2][1] ), .B1(n3521), .B2(n2144), .ZN(
        n2159) );
  OAI22_X1 U3130 ( .A1(n2144), .A2(n2160), .B1(n1179), .B2(n283), .ZN(n7460)
         );
  OAI22_X1 U3132 ( .A1(n2144), .A2(n2161), .B1(n1181), .B2(n283), .ZN(n7461)
         );
  OAI22_X1 U3134 ( .A1(n2144), .A2(n2162), .B1(n1183), .B2(n283), .ZN(n7462)
         );
  OAI22_X1 U3136 ( .A1(n2144), .A2(n2163), .B1(n1185), .B2(n283), .ZN(n7463)
         );
  OAI22_X1 U3138 ( .A1(n2144), .A2(n2164), .B1(n1187), .B2(n283), .ZN(n7464)
         );
  OAI22_X1 U3140 ( .A1(n2144), .A2(n2165), .B1(n1189), .B2(n283), .ZN(n7465)
         );
  OAI22_X1 U3142 ( .A1(n2144), .A2(n2166), .B1(n1191), .B2(n283), .ZN(n7466)
         );
  OAI22_X1 U3144 ( .A1(n2144), .A2(n2167), .B1(n1193), .B2(n283), .ZN(n7467)
         );
  OAI22_X1 U3146 ( .A1(n2144), .A2(n2168), .B1(n1195), .B2(n283), .ZN(n7468)
         );
  OAI22_X1 U3148 ( .A1(n2144), .A2(n2169), .B1(n1197), .B2(n283), .ZN(n7469)
         );
  OAI22_X1 U3150 ( .A1(n2144), .A2(n2170), .B1(n1199), .B2(n283), .ZN(n7470)
         );
  OAI22_X1 U3152 ( .A1(n2144), .A2(n2171), .B1(n1201), .B2(n283), .ZN(n7471)
         );
  OAI22_X1 U3154 ( .A1(n2144), .A2(n2172), .B1(n1203), .B2(n283), .ZN(n7472)
         );
  OAI22_X1 U3156 ( .A1(n2144), .A2(n2173), .B1(n1205), .B2(n283), .ZN(n7473)
         );
  INV_X1 U3161 ( .A(PC_write[1]), .ZN(n2142) );
  OAI22_X1 U3162 ( .A1(n2174), .A2(n2175), .B1(n1147), .B2(n2176), .ZN(n7474)
         );
  OAI22_X1 U3163 ( .A1(n2174), .A2(n2177), .B1(n1150), .B2(n2176), .ZN(n7475)
         );
  OAI22_X1 U3164 ( .A1(n2174), .A2(n2178), .B1(n1152), .B2(n2176), .ZN(n7476)
         );
  OAI22_X1 U3165 ( .A1(n2174), .A2(n2179), .B1(n1154), .B2(n2176), .ZN(n7477)
         );
  OAI22_X1 U3166 ( .A1(n2174), .A2(n2180), .B1(n1156), .B2(n2176), .ZN(n7478)
         );
  OAI22_X1 U3167 ( .A1(n2174), .A2(n2181), .B1(n1158), .B2(n2176), .ZN(n7479)
         );
  OAI22_X1 U3168 ( .A1(n2174), .A2(n2182), .B1(n1160), .B2(n2176), .ZN(n7480)
         );
  OAI22_X1 U3169 ( .A1(n2174), .A2(n2183), .B1(n1162), .B2(n2176), .ZN(n7481)
         );
  OAI22_X1 U3170 ( .A1(n2174), .A2(n2184), .B1(n1164), .B2(n2176), .ZN(n7482)
         );
  OAI22_X1 U3171 ( .A1(n2174), .A2(n2185), .B1(n1166), .B2(n2176), .ZN(n7483)
         );
  OAI22_X1 U3172 ( .A1(n2174), .A2(n2186), .B1(n1168), .B2(n2176), .ZN(n7484)
         );
  OAI22_X1 U3173 ( .A1(n2174), .A2(n2187), .B1(n1170), .B2(n2176), .ZN(n7485)
         );
  OAI22_X1 U3174 ( .A1(n2174), .A2(n2188), .B1(n1172), .B2(n2176), .ZN(n7486)
         );
  OAI22_X1 U3177 ( .A1(n2174), .A2(n2191), .B1(n1496), .B2(n2176), .ZN(n7489)
         );
  OAI22_X1 U3180 ( .A1(n2174), .A2(n2194), .B1(n1179), .B2(n2176), .ZN(n7492)
         );
  OAI22_X1 U3181 ( .A1(n2174), .A2(n2195), .B1(n1181), .B2(n2176), .ZN(n7493)
         );
  OAI22_X1 U3182 ( .A1(n2174), .A2(n2196), .B1(n1183), .B2(n2176), .ZN(n7494)
         );
  OAI22_X1 U3183 ( .A1(n2174), .A2(n2197), .B1(n1185), .B2(n2176), .ZN(n7495)
         );
  OAI22_X1 U3184 ( .A1(n2174), .A2(n2198), .B1(n1187), .B2(n2176), .ZN(n7496)
         );
  OAI22_X1 U3185 ( .A1(n2174), .A2(n2199), .B1(n1189), .B2(n2176), .ZN(n7497)
         );
  OAI22_X1 U3186 ( .A1(n2174), .A2(n2200), .B1(n1191), .B2(n2176), .ZN(n7498)
         );
  OAI22_X1 U3187 ( .A1(n2174), .A2(n2201), .B1(n1193), .B2(n2176), .ZN(n7499)
         );
  OAI22_X1 U3188 ( .A1(n2174), .A2(n2202), .B1(n1195), .B2(n2176), .ZN(n7500)
         );
  OAI22_X1 U3189 ( .A1(n2174), .A2(n2203), .B1(n1197), .B2(n2176), .ZN(n7501)
         );
  OAI22_X1 U3190 ( .A1(n2174), .A2(n2204), .B1(n1199), .B2(n2176), .ZN(n7502)
         );
  OAI22_X1 U3191 ( .A1(n2174), .A2(n2205), .B1(n1201), .B2(n2176), .ZN(n7503)
         );
  OAI22_X1 U3192 ( .A1(n2174), .A2(n2206), .B1(n1203), .B2(n2176), .ZN(n7504)
         );
  OAI22_X1 U3193 ( .A1(n2174), .A2(n2207), .B1(n1205), .B2(n2176), .ZN(n7505)
         );
  INV_X1 U3197 ( .A(PC_write[0]), .ZN(n2143) );
  OAI22_X1 U3198 ( .A1(n2208), .A2(n2209), .B1(n1147), .B2(n2210), .ZN(n7506)
         );
  OAI22_X1 U3200 ( .A1(n2208), .A2(n2211), .B1(n1150), .B2(n2210), .ZN(n7507)
         );
  OAI22_X1 U3202 ( .A1(n2208), .A2(n2212), .B1(n1152), .B2(n2210), .ZN(n7508)
         );
  OAI22_X1 U3204 ( .A1(n2208), .A2(n2213), .B1(n1154), .B2(n2210), .ZN(n7509)
         );
  OAI22_X1 U3206 ( .A1(n2208), .A2(n2214), .B1(n1156), .B2(n2210), .ZN(n7510)
         );
  OAI22_X1 U3208 ( .A1(n2208), .A2(n2215), .B1(n1158), .B2(n2210), .ZN(n7511)
         );
  OAI22_X1 U3210 ( .A1(n2208), .A2(n2216), .B1(n1160), .B2(n2210), .ZN(n7512)
         );
  OAI22_X1 U3212 ( .A1(n2208), .A2(n2217), .B1(n1162), .B2(n2210), .ZN(n7513)
         );
  OAI22_X1 U3214 ( .A1(n2208), .A2(n2218), .B1(n1164), .B2(n2210), .ZN(n7514)
         );
  OAI22_X1 U3216 ( .A1(n2208), .A2(n2219), .B1(n1166), .B2(n2210), .ZN(n7515)
         );
  OAI22_X1 U3218 ( .A1(n2208), .A2(n2220), .B1(n1168), .B2(n2210), .ZN(n7516)
         );
  OAI22_X1 U3220 ( .A1(n2208), .A2(n2221), .B1(n1170), .B2(n2210), .ZN(n7517)
         );
  OAI22_X1 U3222 ( .A1(n2208), .A2(n2222), .B1(n1172), .B2(n2210), .ZN(n7518)
         );
  OAI22_X1 U3229 ( .A1(n2208), .A2(n2228), .B1(n1179), .B2(n2210), .ZN(n7524)
         );
  OAI22_X1 U3231 ( .A1(n2208), .A2(n2229), .B1(n1181), .B2(n2210), .ZN(n7525)
         );
  OAI22_X1 U3233 ( .A1(n2208), .A2(n2230), .B1(n1183), .B2(n2210), .ZN(n7526)
         );
  OAI22_X1 U3235 ( .A1(n2208), .A2(n2231), .B1(n1185), .B2(n2210), .ZN(n7527)
         );
  OAI22_X1 U3237 ( .A1(n2208), .A2(n2232), .B1(n1187), .B2(n2210), .ZN(n7528)
         );
  OAI22_X1 U3239 ( .A1(n2208), .A2(n2233), .B1(n1189), .B2(n2210), .ZN(n7529)
         );
  OAI22_X1 U3241 ( .A1(n2208), .A2(n2234), .B1(n1191), .B2(n2210), .ZN(n7530)
         );
  OAI22_X1 U3243 ( .A1(n2208), .A2(n2235), .B1(n1193), .B2(n2210), .ZN(n7531)
         );
  OAI22_X1 U3245 ( .A1(n2208), .A2(n2236), .B1(n1195), .B2(n2210), .ZN(n7532)
         );
  OAI22_X1 U3247 ( .A1(n2208), .A2(n2237), .B1(n1197), .B2(n2210), .ZN(n7533)
         );
  OAI22_X1 U3249 ( .A1(n2208), .A2(n2238), .B1(n1199), .B2(n2210), .ZN(n7534)
         );
  OAI22_X1 U3251 ( .A1(n2208), .A2(n2239), .B1(n1201), .B2(n2210), .ZN(n7535)
         );
  OAI22_X1 U3253 ( .A1(n2208), .A2(n2240), .B1(n1203), .B2(n2210), .ZN(n7536)
         );
  OAI22_X1 U3255 ( .A1(n2208), .A2(n2241), .B1(n1205), .B2(n2210), .ZN(n7537)
         );
  AND2_X1 U3260 ( .A1(n3794), .A2(n592), .ZN(n2141) );
  NOR2_X1 U3261 ( .A1(PC_write[2]), .A2(PC_write[3]), .ZN(n592) );
  NOR2_X1 U3262 ( .A1(n1708), .A2(PC_write[4]), .ZN(n1843) );
  OAI211_X1 U3263 ( .C1(n3528), .C2(n1144), .A(Enable), .B(WR), .ZN(n1708) );
  INV_X1 U3264 ( .A(prevT_NT), .ZN(n1144) );
  NAND2_X1 U3266 ( .A1(n2242), .A2(n2243), .ZN(N99) );
  NOR4_X1 U3267 ( .A1(n2244), .A2(n2245), .A3(n2246), .A4(n2247), .ZN(n2243)
         );
  OAI221_X1 U3268 ( .B1(n285), .B2(n2248), .C1(n251), .C2(n2249), .A(n2250), 
        .ZN(n2247) );
  AOI22_X1 U3269 ( .A1(n2251), .A2(\pc_target[26][28] ), .B1(n2252), .B2(
        \pc_target[27][28] ), .ZN(n2250) );
  OAI221_X1 U3272 ( .B1(n145), .B2(n2253), .C1(n80), .C2(n2254), .A(n2255), 
        .ZN(n2246) );
  AOI22_X1 U3273 ( .A1(n2256), .A2(\pc_target[30][28] ), .B1(n2257), .B2(
        \pc_target[31][28] ), .ZN(n2255) );
  OAI221_X1 U3276 ( .B1(n561), .B2(n2258), .C1(n527), .C2(n2259), .A(n2260), 
        .ZN(n2245) );
  AOI22_X1 U3277 ( .A1(n2261), .A2(\pc_target[18][28] ), .B1(n2262), .B2(
        \pc_target[19][28] ), .ZN(n2260) );
  OAI221_X1 U3280 ( .B1(n355), .B2(n2263), .C1(n320), .C2(n2264), .A(n2265), 
        .ZN(n2244) );
  AOI22_X1 U3281 ( .A1(n2266), .A2(\pc_target[20][28] ), .B1(n2267), .B2(
        \pc_target[21][28] ), .ZN(n2265) );
  NOR4_X1 U3284 ( .A1(n2268), .A2(n2269), .A3(n2270), .A4(n2271), .ZN(n2242)
         );
  OAI221_X1 U3285 ( .B1(n838), .B2(n2272), .C1(n804), .C2(n2273), .A(n2274), 
        .ZN(n2271) );
  AOI22_X1 U3286 ( .A1(n2275), .A2(\pc_target[10][28] ), .B1(n2276), .B2(
        \pc_target[11][28] ), .ZN(n2274) );
  OAI221_X1 U3289 ( .B1(n700), .B2(n2277), .C1(n666), .C2(n2278), .A(n2279), 
        .ZN(n2270) );
  AOI22_X1 U3290 ( .A1(n2280), .A2(\pc_target[14][28] ), .B1(n2281), .B2(
        \pc_target[15][28] ), .ZN(n2279) );
  OAI221_X1 U3293 ( .B1(n1112), .B2(n2282), .C1(n1078), .C2(n2283), .A(n2284), 
        .ZN(n2269) );
  AOI22_X1 U3294 ( .A1(n2285), .A2(\pc_target[2][28] ), .B1(n2286), .B2(
        \pc_target[3][28] ), .ZN(n2284) );
  OAI221_X1 U3297 ( .B1(n975), .B2(n2287), .C1(n941), .C2(n2288), .A(n2289), 
        .ZN(n2268) );
  AOI22_X1 U3298 ( .A1(n2290), .A2(\pc_target[6][28] ), .B1(n2291), .B2(
        \pc_target[7][28] ), .ZN(n2289) );
  NAND2_X1 U3301 ( .A1(n2292), .A2(n2293), .ZN(N98) );
  NOR4_X1 U3302 ( .A1(n2294), .A2(n2295), .A3(n2296), .A4(n2297), .ZN(n2293)
         );
  OAI221_X1 U3303 ( .B1(n314), .B2(n2248), .C1(n280), .C2(n2249), .A(n2298), 
        .ZN(n2297) );
  AOI22_X1 U3304 ( .A1(n2251), .A2(\pc_target[26][29] ), .B1(n2252), .B2(
        \pc_target[27][29] ), .ZN(n2298) );
  OAI221_X1 U3307 ( .B1(n174), .B2(n2253), .C1(n138), .C2(n2254), .A(n2299), 
        .ZN(n2296) );
  AOI22_X1 U3308 ( .A1(n2256), .A2(\pc_target[30][29] ), .B1(n2257), .B2(
        \pc_target[31][29] ), .ZN(n2299) );
  OAI221_X1 U3311 ( .B1(n590), .B2(n2258), .C1(n556), .C2(n2259), .A(n2300), 
        .ZN(n2295) );
  AOI22_X1 U3312 ( .A1(n2261), .A2(\pc_target[18][29] ), .B1(n2262), .B2(
        \pc_target[19][29] ), .ZN(n2300) );
  OAI221_X1 U3315 ( .B1(n384), .B2(n2263), .C1(n349), .C2(n2264), .A(n2301), 
        .ZN(n2294) );
  AOI22_X1 U3316 ( .A1(n2266), .A2(\pc_target[20][29] ), .B1(n2267), .B2(
        \pc_target[21][29] ), .ZN(n2301) );
  NOR4_X1 U3319 ( .A1(n2302), .A2(n2303), .A3(n2304), .A4(n2305), .ZN(n2292)
         );
  OAI221_X1 U3320 ( .B1(n867), .B2(n2272), .C1(n833), .C2(n2273), .A(n2306), 
        .ZN(n2305) );
  AOI22_X1 U3321 ( .A1(n2275), .A2(\pc_target[10][29] ), .B1(n2276), .B2(
        \pc_target[11][29] ), .ZN(n2306) );
  OAI221_X1 U3324 ( .B1(n729), .B2(n2277), .C1(n695), .C2(n2278), .A(n2307), 
        .ZN(n2304) );
  AOI22_X1 U3325 ( .A1(n2280), .A2(\pc_target[14][29] ), .B1(n2281), .B2(
        \pc_target[15][29] ), .ZN(n2307) );
  OAI221_X1 U3328 ( .B1(n1141), .B2(n2282), .C1(n1107), .C2(n2283), .A(n2308), 
        .ZN(n2303) );
  AOI22_X1 U3329 ( .A1(n2285), .A2(\pc_target[2][29] ), .B1(n2286), .B2(
        \pc_target[3][29] ), .ZN(n2308) );
  OAI221_X1 U3332 ( .B1(n1004), .B2(n2287), .C1(n970), .C2(n2288), .A(n2309), 
        .ZN(n2302) );
  AOI22_X1 U3333 ( .A1(n2290), .A2(\pc_target[6][29] ), .B1(n2291), .B2(
        \pc_target[7][29] ), .ZN(n2309) );
  NAND2_X1 U3336 ( .A1(n2310), .A2(n2311), .ZN(N97) );
  NOR4_X1 U3337 ( .A1(n2312), .A2(n2313), .A3(n2314), .A4(n2315), .ZN(n2311)
         );
  OAI221_X1 U3338 ( .B1(n284), .B2(n2248), .C1(n250), .C2(n2249), .A(n2316), 
        .ZN(n2315) );
  AOI22_X1 U3339 ( .A1(n2251), .A2(\pc_target[26][30] ), .B1(n2252), .B2(
        \pc_target[27][30] ), .ZN(n2316) );
  OAI221_X1 U3342 ( .B1(n144), .B2(n2253), .C1(n78), .C2(n2254), .A(n2317), 
        .ZN(n2314) );
  AOI22_X1 U3343 ( .A1(n2256), .A2(\pc_target[30][30] ), .B1(n2257), .B2(
        \pc_target[31][30] ), .ZN(n2317) );
  OAI221_X1 U3346 ( .B1(n560), .B2(n2258), .C1(n526), .C2(n2259), .A(n2318), 
        .ZN(n2313) );
  AOI22_X1 U3347 ( .A1(n2261), .A2(\pc_target[18][30] ), .B1(n2262), .B2(
        \pc_target[19][30] ), .ZN(n2318) );
  OAI221_X1 U3350 ( .B1(n354), .B2(n2263), .C1(n319), .C2(n2264), .A(n2319), 
        .ZN(n2312) );
  AOI22_X1 U3351 ( .A1(n2266), .A2(\pc_target[20][30] ), .B1(n2267), .B2(
        \pc_target[21][30] ), .ZN(n2319) );
  NOR4_X1 U3354 ( .A1(n2320), .A2(n2321), .A3(n2322), .A4(n2323), .ZN(n2310)
         );
  OAI221_X1 U3355 ( .B1(n837), .B2(n2272), .C1(n803), .C2(n2273), .A(n2324), 
        .ZN(n2323) );
  AOI22_X1 U3356 ( .A1(n2275), .A2(\pc_target[10][30] ), .B1(n2276), .B2(
        \pc_target[11][30] ), .ZN(n2324) );
  OAI221_X1 U3359 ( .B1(n699), .B2(n2277), .C1(n665), .C2(n2278), .A(n2325), 
        .ZN(n2322) );
  AOI22_X1 U3360 ( .A1(n2280), .A2(\pc_target[14][30] ), .B1(n2281), .B2(
        \pc_target[15][30] ), .ZN(n2325) );
  OAI221_X1 U3363 ( .B1(n1111), .B2(n2282), .C1(n1077), .C2(n2283), .A(n2326), 
        .ZN(n2321) );
  AOI22_X1 U3364 ( .A1(n2285), .A2(\pc_target[2][30] ), .B1(n2286), .B2(
        \pc_target[3][30] ), .ZN(n2326) );
  OAI221_X1 U3367 ( .B1(n974), .B2(n2287), .C1(n940), .C2(n2288), .A(n2327), 
        .ZN(n2320) );
  AOI22_X1 U3368 ( .A1(n2290), .A2(\pc_target[6][30] ), .B1(n2291), .B2(
        \pc_target[7][30] ), .ZN(n2327) );
  NAND2_X1 U3371 ( .A1(n2328), .A2(n2329), .ZN(N96) );
  NOR4_X1 U3372 ( .A1(n2330), .A2(n2331), .A3(n2332), .A4(n2333), .ZN(n2329)
         );
  OAI221_X1 U3373 ( .B1(n315), .B2(n2248), .C1(n281), .C2(n2249), .A(n2334), 
        .ZN(n2333) );
  AOI22_X1 U3374 ( .A1(n2251), .A2(\pc_target[26][31] ), .B1(n2252), .B2(
        \pc_target[27][31] ), .ZN(n2334) );
  OAI221_X1 U3377 ( .B1(n175), .B2(n2253), .C1(n140), .C2(n2254), .A(n2335), 
        .ZN(n2332) );
  AOI22_X1 U3378 ( .A1(n2256), .A2(\pc_target[30][31] ), .B1(n2257), .B2(
        \pc_target[31][31] ), .ZN(n2335) );
  OAI221_X1 U3381 ( .B1(n591), .B2(n2258), .C1(n557), .C2(n2259), .A(n2336), 
        .ZN(n2331) );
  AOI22_X1 U3382 ( .A1(n2261), .A2(\pc_target[18][31] ), .B1(n2262), .B2(
        \pc_target[19][31] ), .ZN(n2336) );
  OAI221_X1 U3385 ( .B1(n385), .B2(n2263), .C1(n350), .C2(n2264), .A(n2337), 
        .ZN(n2330) );
  AOI22_X1 U3386 ( .A1(n2266), .A2(\pc_target[20][31] ), .B1(n2267), .B2(
        \pc_target[21][31] ), .ZN(n2337) );
  NOR4_X1 U3389 ( .A1(n2338), .A2(n2339), .A3(n2340), .A4(n2341), .ZN(n2328)
         );
  OAI221_X1 U3390 ( .B1(n868), .B2(n2272), .C1(n834), .C2(n2273), .A(n2342), 
        .ZN(n2341) );
  AOI22_X1 U3391 ( .A1(n2275), .A2(\pc_target[10][31] ), .B1(n2276), .B2(
        \pc_target[11][31] ), .ZN(n2342) );
  OAI221_X1 U3394 ( .B1(n730), .B2(n2277), .C1(n696), .C2(n2278), .A(n2343), 
        .ZN(n2340) );
  AOI22_X1 U3395 ( .A1(n2280), .A2(\pc_target[14][31] ), .B1(n2281), .B2(
        \pc_target[15][31] ), .ZN(n2343) );
  OAI221_X1 U3398 ( .B1(n1142), .B2(n2282), .C1(n1108), .C2(n2283), .A(n2344), 
        .ZN(n2339) );
  AOI22_X1 U3399 ( .A1(n2285), .A2(\pc_target[2][31] ), .B1(n2286), .B2(
        \pc_target[3][31] ), .ZN(n2344) );
  OAI221_X1 U3402 ( .B1(n1005), .B2(n2287), .C1(n971), .C2(n2288), .A(n2345), 
        .ZN(n2338) );
  AOI22_X1 U3403 ( .A1(n2290), .A2(\pc_target[6][31] ), .B1(n2291), .B2(
        \pc_target[7][31] ), .ZN(n2345) );
  NAND2_X1 U3406 ( .A1(n2346), .A2(n2347), .ZN(N219) );
  NOR4_X1 U3407 ( .A1(n2348), .A2(n2349), .A3(n2350), .A4(n2351), .ZN(n2347)
         );
  NOR4_X1 U3424 ( .A1(n2356), .A2(n2357), .A3(n2358), .A4(n2359), .ZN(n2346)
         );
  NAND2_X1 U3441 ( .A1(n2364), .A2(n2365), .ZN(N218) );
  NOR4_X1 U3442 ( .A1(n2366), .A2(n2367), .A3(n2368), .A4(n2369), .ZN(n2365)
         );
  AOI22_X1 U3444 ( .A1(n2251), .A2(\pc_lut[26][1] ), .B1(n2252), .B2(
        \pc_lut[27][1] ), .ZN(n2370) );
  AOI22_X1 U3448 ( .A1(n2256), .A2(\pc_lut[30][1] ), .B1(n2257), .B2(
        \pc_lut[31][1] ), .ZN(n2371) );
  AOI22_X1 U3452 ( .A1(n2261), .A2(\pc_lut[18][1] ), .B1(n2262), .B2(
        \pc_lut[19][1] ), .ZN(n2372) );
  NOR4_X1 U3459 ( .A1(n2374), .A2(n2375), .A3(n2376), .A4(n2377), .ZN(n2364)
         );
  AOI22_X1 U3461 ( .A1(n2275), .A2(\pc_lut[10][1] ), .B1(n2276), .B2(
        \pc_lut[11][1] ), .ZN(n2378) );
  AOI22_X1 U3465 ( .A1(n2280), .A2(\pc_lut[14][1] ), .B1(n2281), .B2(
        \pc_lut[15][1] ), .ZN(n2379) );
  AOI22_X1 U3469 ( .A1(n2285), .A2(\pc_lut[2][1] ), .B1(n2286), .B2(
        \pc_lut[3][1] ), .ZN(n2380) );
  AOI22_X1 U3473 ( .A1(n2290), .A2(\pc_lut[6][1] ), .B1(n2291), .B2(
        \pc_lut[7][1] ), .ZN(n2381) );
  NAND2_X1 U3476 ( .A1(n2382), .A2(n2383), .ZN(N217) );
  OAI221_X1 U3482 ( .B1(n1291), .B2(n2253), .C1(n1257), .C2(n2254), .A(n2389), 
        .ZN(n2386) );
  AOI22_X1 U3483 ( .A1(n2256), .A2(\pc_lut[30][2] ), .B1(n2257), .B2(
        \pc_lut[31][2] ), .ZN(n2389) );
  OAI221_X1 U3490 ( .B1(n1495), .B2(n2263), .C1(n1460), .C2(n2264), .A(n2391), 
        .ZN(n2384) );
  AOI22_X1 U3491 ( .A1(n2266), .A2(\pc_lut[20][2] ), .B1(n2267), .B2(
        \pc_lut[21][2] ), .ZN(n2391) );
  OAI221_X1 U3499 ( .B1(n1825), .B2(n2277), .C1(n1791), .C2(n2278), .A(n2397), 
        .ZN(n2394) );
  AOI22_X1 U3500 ( .A1(n2280), .A2(\pc_lut[14][2] ), .B1(n2281), .B2(
        \pc_lut[15][2] ), .ZN(n2397) );
  OAI221_X1 U3507 ( .B1(n2092), .B2(n2287), .C1(n2058), .C2(n2288), .A(n2399), 
        .ZN(n2392) );
  AOI22_X1 U3508 ( .A1(n2290), .A2(\pc_lut[6][2] ), .B1(n2291), .B2(
        \pc_lut[7][2] ), .ZN(n2399) );
  NAND2_X1 U3511 ( .A1(n2400), .A2(n2401), .ZN(N216) );
  OAI221_X1 U3513 ( .B1(n1429), .B2(n2248), .C1(n1395), .C2(n2249), .A(n2406), 
        .ZN(n2405) );
  AOI22_X1 U3514 ( .A1(n2251), .A2(\pc_lut[26][3] ), .B1(n2252), .B2(
        \pc_lut[27][3] ), .ZN(n2406) );
  OAI221_X1 U3517 ( .B1(n1294), .B2(n2253), .C1(n1260), .C2(n2254), .A(n2407), 
        .ZN(n2404) );
  AOI22_X1 U3518 ( .A1(n2256), .A2(\pc_lut[30][3] ), .B1(n2257), .B2(
        \pc_lut[31][3] ), .ZN(n2407) );
  OAI221_X1 U3530 ( .B1(n1963), .B2(n2272), .C1(n1929), .C2(n2273), .A(n2414), 
        .ZN(n2413) );
  AOI22_X1 U3531 ( .A1(n2275), .A2(\pc_lut[10][3] ), .B1(n2276), .B2(
        \pc_lut[11][3] ), .ZN(n2414) );
  OAI221_X1 U3534 ( .B1(n1828), .B2(n2277), .C1(n1794), .C2(n2278), .A(n2415), 
        .ZN(n2412) );
  AOI22_X1 U3535 ( .A1(n2280), .A2(\pc_lut[14][3] ), .B1(n2281), .B2(
        \pc_lut[15][3] ), .ZN(n2415) );
  NOR4_X1 U3547 ( .A1(n2420), .A2(n2421), .A3(n2422), .A4(n2423), .ZN(n2419)
         );
  OAI221_X1 U3548 ( .B1(n1425), .B2(n2248), .C1(n1391), .C2(n2249), .A(n2424), 
        .ZN(n2423) );
  AOI22_X1 U3549 ( .A1(n2251), .A2(\pc_lut[26][4] ), .B1(n2252), .B2(
        \pc_lut[27][4] ), .ZN(n2424) );
  OAI221_X1 U3552 ( .B1(n1290), .B2(n2253), .C1(n1255), .C2(n2254), .A(n2425), 
        .ZN(n2422) );
  AOI22_X1 U3553 ( .A1(n2256), .A2(\pc_lut[30][4] ), .B1(n2257), .B2(
        \pc_lut[31][4] ), .ZN(n2425) );
  OAI221_X1 U3556 ( .B1(n1689), .B2(n2258), .C1(n1655), .C2(n2259), .A(n2426), 
        .ZN(n2421) );
  AOI22_X1 U3557 ( .A1(n2261), .A2(\pc_lut[18][4] ), .B1(n2262), .B2(
        \pc_lut[19][4] ), .ZN(n2426) );
  OAI221_X1 U3560 ( .B1(n1494), .B2(n2263), .C1(n1459), .C2(n2264), .A(n2427), 
        .ZN(n2420) );
  AOI22_X1 U3561 ( .A1(n2266), .A2(\pc_lut[20][4] ), .B1(n2267), .B2(
        \pc_lut[21][4] ), .ZN(n2427) );
  NAND2_X1 U3581 ( .A1(n2436), .A2(n2437), .ZN(N214) );
  NOR4_X1 U3582 ( .A1(n2438), .A2(n2439), .A3(n2440), .A4(n2441), .ZN(n2437)
         );
  OAI221_X1 U3583 ( .B1(n1430), .B2(n2248), .C1(n1396), .C2(n2249), .A(n2442), 
        .ZN(n2441) );
  AOI22_X1 U3584 ( .A1(n2251), .A2(\pc_lut[26][5] ), .B1(n2252), .B2(
        \pc_lut[27][5] ), .ZN(n2442) );
  OAI221_X1 U3587 ( .B1(n1295), .B2(n2253), .C1(n1261), .C2(n2254), .A(n2443), 
        .ZN(n2440) );
  AOI22_X1 U3588 ( .A1(n2256), .A2(\pc_lut[30][5] ), .B1(n2257), .B2(
        \pc_lut[31][5] ), .ZN(n2443) );
  OAI221_X1 U3591 ( .B1(n1694), .B2(n2258), .C1(n1660), .C2(n2259), .A(n2444), 
        .ZN(n2439) );
  AOI22_X1 U3592 ( .A1(n2261), .A2(\pc_lut[18][5] ), .B1(n2262), .B2(
        \pc_lut[19][5] ), .ZN(n2444) );
  OAI221_X1 U3595 ( .B1(n1499), .B2(n2263), .C1(n1464), .C2(n2264), .A(n2445), 
        .ZN(n2438) );
  AOI22_X1 U3596 ( .A1(n2266), .A2(\pc_lut[20][5] ), .B1(n2267), .B2(
        \pc_lut[21][5] ), .ZN(n2445) );
  NOR4_X1 U3599 ( .A1(n2446), .A2(n2447), .A3(n2448), .A4(n2449), .ZN(n2436)
         );
  OAI221_X1 U3600 ( .B1(n1964), .B2(n2272), .C1(n1930), .C2(n2273), .A(n2450), 
        .ZN(n2449) );
  AOI22_X1 U3601 ( .A1(n2275), .A2(\pc_lut[10][5] ), .B1(n2276), .B2(
        \pc_lut[11][5] ), .ZN(n2450) );
  OAI221_X1 U3604 ( .B1(n1829), .B2(n2277), .C1(n1795), .C2(n2278), .A(n2451), 
        .ZN(n2448) );
  AOI22_X1 U3605 ( .A1(n2280), .A2(\pc_lut[14][5] ), .B1(n2281), .B2(
        \pc_lut[15][5] ), .ZN(n2451) );
  OAI221_X1 U3608 ( .B1(n2228), .B2(n2282), .C1(n2194), .C2(n2283), .A(n2452), 
        .ZN(n2447) );
  AOI22_X1 U3609 ( .A1(n2285), .A2(\pc_lut[2][5] ), .B1(n2286), .B2(
        \pc_lut[3][5] ), .ZN(n2452) );
  OAI221_X1 U3612 ( .B1(n2096), .B2(n2287), .C1(n2062), .C2(n2288), .A(n2453), 
        .ZN(n2446) );
  AOI22_X1 U3613 ( .A1(n2290), .A2(\pc_lut[6][5] ), .B1(n2291), .B2(
        \pc_lut[7][5] ), .ZN(n2453) );
  NAND2_X1 U3616 ( .A1(n2454), .A2(n2455), .ZN(N213) );
  NOR4_X1 U3617 ( .A1(n2456), .A2(n2457), .A3(n2458), .A4(n2459), .ZN(n2455)
         );
  OAI221_X1 U3618 ( .B1(n1424), .B2(n2248), .C1(n1390), .C2(n2249), .A(n2460), 
        .ZN(n2459) );
  AOI22_X1 U3619 ( .A1(n2251), .A2(\pc_lut[26][6] ), .B1(n2252), .B2(
        \pc_lut[27][6] ), .ZN(n2460) );
  OAI221_X1 U3622 ( .B1(n1289), .B2(n2253), .C1(n1254), .C2(n2254), .A(n2461), 
        .ZN(n2458) );
  AOI22_X1 U3623 ( .A1(n2256), .A2(\pc_lut[30][6] ), .B1(n2257), .B2(
        \pc_lut[31][6] ), .ZN(n2461) );
  OAI221_X1 U3626 ( .B1(n1688), .B2(n2258), .C1(n1654), .C2(n2259), .A(n2462), 
        .ZN(n2457) );
  AOI22_X1 U3627 ( .A1(n2261), .A2(\pc_lut[18][6] ), .B1(n2262), .B2(
        \pc_lut[19][6] ), .ZN(n2462) );
  OAI221_X1 U3630 ( .B1(n1493), .B2(n2263), .C1(n1458), .C2(n2264), .A(n2463), 
        .ZN(n2456) );
  AOI22_X1 U3631 ( .A1(n2266), .A2(\pc_lut[20][6] ), .B1(n2267), .B2(
        \pc_lut[21][6] ), .ZN(n2463) );
  NOR4_X1 U3634 ( .A1(n2464), .A2(n2465), .A3(n2466), .A4(n2467), .ZN(n2454)
         );
  OAI221_X1 U3635 ( .B1(n1958), .B2(n2272), .C1(n1924), .C2(n2273), .A(n2468), 
        .ZN(n2467) );
  AOI22_X1 U3636 ( .A1(n2275), .A2(\pc_lut[10][6] ), .B1(n2276), .B2(
        \pc_lut[11][6] ), .ZN(n2468) );
  OAI221_X1 U3639 ( .B1(n1823), .B2(n2277), .C1(n1789), .C2(n2278), .A(n2469), 
        .ZN(n2466) );
  AOI22_X1 U3640 ( .A1(n2280), .A2(\pc_lut[14][6] ), .B1(n2281), .B2(
        \pc_lut[15][6] ), .ZN(n2469) );
  OAI221_X1 U3643 ( .B1(n2222), .B2(n2282), .C1(n2188), .C2(n2283), .A(n2470), 
        .ZN(n2465) );
  AOI22_X1 U3644 ( .A1(n2285), .A2(\pc_lut[2][6] ), .B1(n2286), .B2(
        \pc_lut[3][6] ), .ZN(n2470) );
  OAI221_X1 U3647 ( .B1(n2090), .B2(n2287), .C1(n2056), .C2(n2288), .A(n2471), 
        .ZN(n2464) );
  AOI22_X1 U3648 ( .A1(n2290), .A2(\pc_lut[6][6] ), .B1(n2291), .B2(
        \pc_lut[7][6] ), .ZN(n2471) );
  NAND2_X1 U3651 ( .A1(n2472), .A2(n2473), .ZN(N212) );
  NOR4_X1 U3652 ( .A1(n2474), .A2(n2475), .A3(n2476), .A4(n2477), .ZN(n2473)
         );
  OAI221_X1 U3653 ( .B1(n1431), .B2(n2248), .C1(n1397), .C2(n2249), .A(n2478), 
        .ZN(n2477) );
  AOI22_X1 U3654 ( .A1(n2251), .A2(\pc_lut[26][7] ), .B1(n2252), .B2(
        \pc_lut[27][7] ), .ZN(n2478) );
  OAI221_X1 U3657 ( .B1(n1296), .B2(n2253), .C1(n1262), .C2(n2254), .A(n2479), 
        .ZN(n2476) );
  AOI22_X1 U3658 ( .A1(n2256), .A2(\pc_lut[30][7] ), .B1(n2257), .B2(
        \pc_lut[31][7] ), .ZN(n2479) );
  OAI221_X1 U3661 ( .B1(n1695), .B2(n2258), .C1(n1661), .C2(n2259), .A(n2480), 
        .ZN(n2475) );
  AOI22_X1 U3662 ( .A1(n2261), .A2(\pc_lut[18][7] ), .B1(n2262), .B2(
        \pc_lut[19][7] ), .ZN(n2480) );
  OAI221_X1 U3665 ( .B1(n1500), .B2(n2263), .C1(n1465), .C2(n2264), .A(n2481), 
        .ZN(n2474) );
  AOI22_X1 U3666 ( .A1(n2266), .A2(\pc_lut[20][7] ), .B1(n2267), .B2(
        \pc_lut[21][7] ), .ZN(n2481) );
  NOR4_X1 U3669 ( .A1(n2482), .A2(n2483), .A3(n2484), .A4(n2485), .ZN(n2472)
         );
  OAI221_X1 U3670 ( .B1(n1965), .B2(n2272), .C1(n1931), .C2(n2273), .A(n2486), 
        .ZN(n2485) );
  AOI22_X1 U3671 ( .A1(n2275), .A2(\pc_lut[10][7] ), .B1(n2276), .B2(
        \pc_lut[11][7] ), .ZN(n2486) );
  OAI221_X1 U3674 ( .B1(n1830), .B2(n2277), .C1(n1796), .C2(n2278), .A(n2487), 
        .ZN(n2484) );
  AOI22_X1 U3675 ( .A1(n2280), .A2(\pc_lut[14][7] ), .B1(n2281), .B2(
        \pc_lut[15][7] ), .ZN(n2487) );
  OAI221_X1 U3678 ( .B1(n2229), .B2(n2282), .C1(n2195), .C2(n2283), .A(n2488), 
        .ZN(n2483) );
  AOI22_X1 U3679 ( .A1(n2285), .A2(\pc_lut[2][7] ), .B1(n2286), .B2(
        \pc_lut[3][7] ), .ZN(n2488) );
  OAI221_X1 U3682 ( .B1(n2097), .B2(n2287), .C1(n2063), .C2(n2288), .A(n2489), 
        .ZN(n2482) );
  AOI22_X1 U3683 ( .A1(n2290), .A2(\pc_lut[6][7] ), .B1(n2291), .B2(
        \pc_lut[7][7] ), .ZN(n2489) );
  NAND2_X1 U3686 ( .A1(n2490), .A2(n2491), .ZN(N211) );
  NOR4_X1 U3687 ( .A1(n2492), .A2(n2493), .A3(n2494), .A4(n2495), .ZN(n2491)
         );
  OAI221_X1 U3688 ( .B1(n1423), .B2(n2248), .C1(n1389), .C2(n2249), .A(n2496), 
        .ZN(n2495) );
  AOI22_X1 U3689 ( .A1(n2251), .A2(\pc_lut[26][8] ), .B1(n2252), .B2(
        \pc_lut[27][8] ), .ZN(n2496) );
  OAI221_X1 U3692 ( .B1(n1288), .B2(n2253), .C1(n1253), .C2(n2254), .A(n2497), 
        .ZN(n2494) );
  AOI22_X1 U3693 ( .A1(n2256), .A2(\pc_lut[30][8] ), .B1(n2257), .B2(
        \pc_lut[31][8] ), .ZN(n2497) );
  OAI221_X1 U3696 ( .B1(n1687), .B2(n2258), .C1(n1653), .C2(n2259), .A(n2498), 
        .ZN(n2493) );
  AOI22_X1 U3697 ( .A1(n2261), .A2(\pc_lut[18][8] ), .B1(n2262), .B2(
        \pc_lut[19][8] ), .ZN(n2498) );
  OAI221_X1 U3700 ( .B1(n1492), .B2(n2263), .C1(n1457), .C2(n2264), .A(n2499), 
        .ZN(n2492) );
  AOI22_X1 U3701 ( .A1(n2266), .A2(\pc_lut[20][8] ), .B1(n2267), .B2(
        \pc_lut[21][8] ), .ZN(n2499) );
  NOR4_X1 U3704 ( .A1(n2500), .A2(n2501), .A3(n2502), .A4(n2503), .ZN(n2490)
         );
  OAI221_X1 U3705 ( .B1(n1957), .B2(n2272), .C1(n1923), .C2(n2273), .A(n2504), 
        .ZN(n2503) );
  AOI22_X1 U3706 ( .A1(n2275), .A2(\pc_lut[10][8] ), .B1(n2276), .B2(
        \pc_lut[11][8] ), .ZN(n2504) );
  OAI221_X1 U3709 ( .B1(n1822), .B2(n2277), .C1(n1788), .C2(n2278), .A(n2505), 
        .ZN(n2502) );
  AOI22_X1 U3710 ( .A1(n2280), .A2(\pc_lut[14][8] ), .B1(n2281), .B2(
        \pc_lut[15][8] ), .ZN(n2505) );
  OAI221_X1 U3713 ( .B1(n2221), .B2(n2282), .C1(n2187), .C2(n2283), .A(n2506), 
        .ZN(n2501) );
  AOI22_X1 U3714 ( .A1(n2285), .A2(\pc_lut[2][8] ), .B1(n2286), .B2(
        \pc_lut[3][8] ), .ZN(n2506) );
  OAI221_X1 U3717 ( .B1(n2089), .B2(n2287), .C1(n2055), .C2(n2288), .A(n2507), 
        .ZN(n2500) );
  AOI22_X1 U3718 ( .A1(n2290), .A2(\pc_lut[6][8] ), .B1(n2291), .B2(
        \pc_lut[7][8] ), .ZN(n2507) );
  NAND2_X1 U3721 ( .A1(n2508), .A2(n2509), .ZN(N210) );
  NOR4_X1 U3722 ( .A1(n2510), .A2(n2511), .A3(n2512), .A4(n2513), .ZN(n2509)
         );
  OAI221_X1 U3723 ( .B1(n1432), .B2(n2248), .C1(n1398), .C2(n2249), .A(n2514), 
        .ZN(n2513) );
  AOI22_X1 U3724 ( .A1(n2251), .A2(\pc_lut[26][9] ), .B1(n2252), .B2(
        \pc_lut[27][9] ), .ZN(n2514) );
  OAI221_X1 U3727 ( .B1(n1297), .B2(n2253), .C1(n1263), .C2(n2254), .A(n2515), 
        .ZN(n2512) );
  AOI22_X1 U3728 ( .A1(n2256), .A2(\pc_lut[30][9] ), .B1(n2257), .B2(
        \pc_lut[31][9] ), .ZN(n2515) );
  OAI221_X1 U3731 ( .B1(n1696), .B2(n2258), .C1(n1662), .C2(n2259), .A(n2516), 
        .ZN(n2511) );
  AOI22_X1 U3732 ( .A1(n2261), .A2(\pc_lut[18][9] ), .B1(n2262), .B2(
        \pc_lut[19][9] ), .ZN(n2516) );
  OAI221_X1 U3735 ( .B1(n1501), .B2(n2263), .C1(n1466), .C2(n2264), .A(n2517), 
        .ZN(n2510) );
  AOI22_X1 U3736 ( .A1(n2266), .A2(\pc_lut[20][9] ), .B1(n2267), .B2(
        \pc_lut[21][9] ), .ZN(n2517) );
  NOR4_X1 U3739 ( .A1(n2518), .A2(n2519), .A3(n2520), .A4(n2521), .ZN(n2508)
         );
  OAI221_X1 U3740 ( .B1(n1966), .B2(n2272), .C1(n1932), .C2(n2273), .A(n2522), 
        .ZN(n2521) );
  AOI22_X1 U3741 ( .A1(n2275), .A2(\pc_lut[10][9] ), .B1(n2276), .B2(
        \pc_lut[11][9] ), .ZN(n2522) );
  OAI221_X1 U3744 ( .B1(n1831), .B2(n2277), .C1(n1797), .C2(n2278), .A(n2523), 
        .ZN(n2520) );
  AOI22_X1 U3745 ( .A1(n2280), .A2(\pc_lut[14][9] ), .B1(n2281), .B2(
        \pc_lut[15][9] ), .ZN(n2523) );
  OAI221_X1 U3748 ( .B1(n2230), .B2(n2282), .C1(n2196), .C2(n2283), .A(n2524), 
        .ZN(n2519) );
  AOI22_X1 U3749 ( .A1(n2285), .A2(\pc_lut[2][9] ), .B1(n2286), .B2(
        \pc_lut[3][9] ), .ZN(n2524) );
  OAI221_X1 U3752 ( .B1(n2098), .B2(n2287), .C1(n2064), .C2(n2288), .A(n2525), 
        .ZN(n2518) );
  AOI22_X1 U3753 ( .A1(n2290), .A2(\pc_lut[6][9] ), .B1(n2291), .B2(
        \pc_lut[7][9] ), .ZN(n2525) );
  NAND2_X1 U3756 ( .A1(n2526), .A2(n2527), .ZN(N209) );
  NOR4_X1 U3757 ( .A1(n2528), .A2(n2529), .A3(n2530), .A4(n2531), .ZN(n2527)
         );
  OAI221_X1 U3758 ( .B1(n1422), .B2(n2248), .C1(n1388), .C2(n2249), .A(n2532), 
        .ZN(n2531) );
  AOI22_X1 U3759 ( .A1(n2251), .A2(\pc_lut[26][10] ), .B1(n2252), .B2(
        \pc_lut[27][10] ), .ZN(n2532) );
  OAI221_X1 U3762 ( .B1(n1287), .B2(n2253), .C1(n1252), .C2(n2254), .A(n2533), 
        .ZN(n2530) );
  AOI22_X1 U3763 ( .A1(n2256), .A2(\pc_lut[30][10] ), .B1(n2257), .B2(
        \pc_lut[31][10] ), .ZN(n2533) );
  OAI221_X1 U3766 ( .B1(n1686), .B2(n2258), .C1(n1652), .C2(n2259), .A(n2534), 
        .ZN(n2529) );
  AOI22_X1 U3767 ( .A1(n2261), .A2(\pc_lut[18][10] ), .B1(n2262), .B2(
        \pc_lut[19][10] ), .ZN(n2534) );
  OAI221_X1 U3770 ( .B1(n1491), .B2(n2263), .C1(n1456), .C2(n2264), .A(n2535), 
        .ZN(n2528) );
  AOI22_X1 U3771 ( .A1(n2266), .A2(\pc_lut[20][10] ), .B1(n2267), .B2(
        \pc_lut[21][10] ), .ZN(n2535) );
  NOR4_X1 U3774 ( .A1(n2536), .A2(n2537), .A3(n2538), .A4(n2539), .ZN(n2526)
         );
  OAI221_X1 U3775 ( .B1(n1956), .B2(n2272), .C1(n1922), .C2(n2273), .A(n2540), 
        .ZN(n2539) );
  AOI22_X1 U3776 ( .A1(n2275), .A2(\pc_lut[10][10] ), .B1(n2276), .B2(
        \pc_lut[11][10] ), .ZN(n2540) );
  OAI221_X1 U3779 ( .B1(n1821), .B2(n2277), .C1(n1787), .C2(n2278), .A(n2541), 
        .ZN(n2538) );
  AOI22_X1 U3780 ( .A1(n2280), .A2(\pc_lut[14][10] ), .B1(n2281), .B2(
        \pc_lut[15][10] ), .ZN(n2541) );
  OAI221_X1 U3783 ( .B1(n2220), .B2(n2282), .C1(n2186), .C2(n2283), .A(n2542), 
        .ZN(n2537) );
  AOI22_X1 U3784 ( .A1(n2285), .A2(\pc_lut[2][10] ), .B1(n2286), .B2(
        \pc_lut[3][10] ), .ZN(n2542) );
  OAI221_X1 U3787 ( .B1(n2088), .B2(n2287), .C1(n2054), .C2(n2288), .A(n2543), 
        .ZN(n2536) );
  AOI22_X1 U3788 ( .A1(n2290), .A2(\pc_lut[6][10] ), .B1(n2291), .B2(
        \pc_lut[7][10] ), .ZN(n2543) );
  NAND2_X1 U3791 ( .A1(n2544), .A2(n2545), .ZN(N208) );
  NOR4_X1 U3792 ( .A1(n2546), .A2(n2547), .A3(n2548), .A4(n2549), .ZN(n2545)
         );
  OAI221_X1 U3793 ( .B1(n1433), .B2(n2248), .C1(n1399), .C2(n2249), .A(n2550), 
        .ZN(n2549) );
  AOI22_X1 U3794 ( .A1(n2251), .A2(\pc_lut[26][11] ), .B1(n2252), .B2(
        \pc_lut[27][11] ), .ZN(n2550) );
  OAI221_X1 U3797 ( .B1(n1298), .B2(n2253), .C1(n1264), .C2(n2254), .A(n2551), 
        .ZN(n2548) );
  AOI22_X1 U3798 ( .A1(n2256), .A2(\pc_lut[30][11] ), .B1(n2257), .B2(
        \pc_lut[31][11] ), .ZN(n2551) );
  OAI221_X1 U3801 ( .B1(n1697), .B2(n2258), .C1(n1663), .C2(n2259), .A(n2552), 
        .ZN(n2547) );
  AOI22_X1 U3802 ( .A1(n2261), .A2(\pc_lut[18][11] ), .B1(n2262), .B2(
        \pc_lut[19][11] ), .ZN(n2552) );
  OAI221_X1 U3805 ( .B1(n1502), .B2(n2263), .C1(n1467), .C2(n2264), .A(n2553), 
        .ZN(n2546) );
  AOI22_X1 U3806 ( .A1(n2266), .A2(\pc_lut[20][11] ), .B1(n2267), .B2(
        \pc_lut[21][11] ), .ZN(n2553) );
  NOR4_X1 U3809 ( .A1(n2554), .A2(n2555), .A3(n2556), .A4(n2557), .ZN(n2544)
         );
  OAI221_X1 U3810 ( .B1(n1967), .B2(n2272), .C1(n1933), .C2(n2273), .A(n2558), 
        .ZN(n2557) );
  AOI22_X1 U3811 ( .A1(n2275), .A2(\pc_lut[10][11] ), .B1(n2276), .B2(
        \pc_lut[11][11] ), .ZN(n2558) );
  OAI221_X1 U3814 ( .B1(n1832), .B2(n2277), .C1(n1798), .C2(n2278), .A(n2559), 
        .ZN(n2556) );
  AOI22_X1 U3815 ( .A1(n2280), .A2(\pc_lut[14][11] ), .B1(n2281), .B2(
        \pc_lut[15][11] ), .ZN(n2559) );
  OAI221_X1 U3818 ( .B1(n2231), .B2(n2282), .C1(n2197), .C2(n2283), .A(n2560), 
        .ZN(n2555) );
  AOI22_X1 U3819 ( .A1(n2285), .A2(\pc_lut[2][11] ), .B1(n2286), .B2(
        \pc_lut[3][11] ), .ZN(n2560) );
  OAI221_X1 U3822 ( .B1(n2099), .B2(n2287), .C1(n2065), .C2(n2288), .A(n2561), 
        .ZN(n2554) );
  AOI22_X1 U3823 ( .A1(n2290), .A2(\pc_lut[6][11] ), .B1(n2291), .B2(
        \pc_lut[7][11] ), .ZN(n2561) );
  NAND2_X1 U3826 ( .A1(n2562), .A2(n2563), .ZN(N207) );
  NOR4_X1 U3827 ( .A1(n2564), .A2(n2565), .A3(n2566), .A4(n2567), .ZN(n2563)
         );
  OAI221_X1 U3828 ( .B1(n1421), .B2(n2248), .C1(n1387), .C2(n2249), .A(n2568), 
        .ZN(n2567) );
  AOI22_X1 U3829 ( .A1(n2251), .A2(\pc_lut[26][12] ), .B1(n2252), .B2(
        \pc_lut[27][12] ), .ZN(n2568) );
  OAI221_X1 U3832 ( .B1(n1286), .B2(n2253), .C1(n1251), .C2(n2254), .A(n2569), 
        .ZN(n2566) );
  AOI22_X1 U3833 ( .A1(n2256), .A2(\pc_lut[30][12] ), .B1(n2257), .B2(
        \pc_lut[31][12] ), .ZN(n2569) );
  OAI221_X1 U3836 ( .B1(n1685), .B2(n2258), .C1(n1651), .C2(n2259), .A(n2570), 
        .ZN(n2565) );
  AOI22_X1 U3837 ( .A1(n2261), .A2(\pc_lut[18][12] ), .B1(n2262), .B2(
        \pc_lut[19][12] ), .ZN(n2570) );
  OAI221_X1 U3840 ( .B1(n1490), .B2(n2263), .C1(n1455), .C2(n2264), .A(n2571), 
        .ZN(n2564) );
  AOI22_X1 U3841 ( .A1(n2266), .A2(\pc_lut[20][12] ), .B1(n2267), .B2(
        \pc_lut[21][12] ), .ZN(n2571) );
  NOR4_X1 U3844 ( .A1(n2572), .A2(n2573), .A3(n2574), .A4(n2575), .ZN(n2562)
         );
  OAI221_X1 U3845 ( .B1(n1955), .B2(n2272), .C1(n1921), .C2(n2273), .A(n2576), 
        .ZN(n2575) );
  AOI22_X1 U3846 ( .A1(n2275), .A2(\pc_lut[10][12] ), .B1(n2276), .B2(
        \pc_lut[11][12] ), .ZN(n2576) );
  OAI221_X1 U3849 ( .B1(n1820), .B2(n2277), .C1(n1786), .C2(n2278), .A(n2577), 
        .ZN(n2574) );
  AOI22_X1 U3850 ( .A1(n2280), .A2(\pc_lut[14][12] ), .B1(n2281), .B2(
        \pc_lut[15][12] ), .ZN(n2577) );
  OAI221_X1 U3853 ( .B1(n2219), .B2(n2282), .C1(n2185), .C2(n2283), .A(n2578), 
        .ZN(n2573) );
  AOI22_X1 U3854 ( .A1(n2285), .A2(\pc_lut[2][12] ), .B1(n2286), .B2(
        \pc_lut[3][12] ), .ZN(n2578) );
  OAI221_X1 U3857 ( .B1(n2087), .B2(n2287), .C1(n2053), .C2(n2288), .A(n2579), 
        .ZN(n2572) );
  AOI22_X1 U3858 ( .A1(n2290), .A2(\pc_lut[6][12] ), .B1(n2291), .B2(
        \pc_lut[7][12] ), .ZN(n2579) );
  NAND2_X1 U3861 ( .A1(n2580), .A2(n2581), .ZN(N206) );
  NOR4_X1 U3862 ( .A1(n2582), .A2(n2583), .A3(n2584), .A4(n2585), .ZN(n2581)
         );
  OAI221_X1 U3863 ( .B1(n1434), .B2(n2248), .C1(n1400), .C2(n2249), .A(n2586), 
        .ZN(n2585) );
  AOI22_X1 U3864 ( .A1(n2251), .A2(\pc_lut[26][13] ), .B1(n2252), .B2(
        \pc_lut[27][13] ), .ZN(n2586) );
  OAI221_X1 U3867 ( .B1(n1299), .B2(n2253), .C1(n1265), .C2(n2254), .A(n2587), 
        .ZN(n2584) );
  AOI22_X1 U3868 ( .A1(n2256), .A2(\pc_lut[30][13] ), .B1(n2257), .B2(
        \pc_lut[31][13] ), .ZN(n2587) );
  OAI221_X1 U3871 ( .B1(n1698), .B2(n2258), .C1(n1664), .C2(n2259), .A(n2588), 
        .ZN(n2583) );
  AOI22_X1 U3872 ( .A1(n2261), .A2(\pc_lut[18][13] ), .B1(n2262), .B2(
        \pc_lut[19][13] ), .ZN(n2588) );
  OAI221_X1 U3875 ( .B1(n1503), .B2(n2263), .C1(n1468), .C2(n2264), .A(n2589), 
        .ZN(n2582) );
  AOI22_X1 U3876 ( .A1(n2266), .A2(\pc_lut[20][13] ), .B1(n2267), .B2(
        \pc_lut[21][13] ), .ZN(n2589) );
  NOR4_X1 U3879 ( .A1(n2590), .A2(n2591), .A3(n2592), .A4(n2593), .ZN(n2580)
         );
  OAI221_X1 U3880 ( .B1(n1968), .B2(n2272), .C1(n1934), .C2(n2273), .A(n2594), 
        .ZN(n2593) );
  AOI22_X1 U3881 ( .A1(n2275), .A2(\pc_lut[10][13] ), .B1(n2276), .B2(
        \pc_lut[11][13] ), .ZN(n2594) );
  OAI221_X1 U3884 ( .B1(n1833), .B2(n2277), .C1(n1799), .C2(n2278), .A(n2595), 
        .ZN(n2592) );
  AOI22_X1 U3885 ( .A1(n2280), .A2(\pc_lut[14][13] ), .B1(n2281), .B2(
        \pc_lut[15][13] ), .ZN(n2595) );
  OAI221_X1 U3888 ( .B1(n2232), .B2(n2282), .C1(n2198), .C2(n2283), .A(n2596), 
        .ZN(n2591) );
  AOI22_X1 U3889 ( .A1(n2285), .A2(\pc_lut[2][13] ), .B1(n2286), .B2(
        \pc_lut[3][13] ), .ZN(n2596) );
  OAI221_X1 U3892 ( .B1(n2100), .B2(n2287), .C1(n2066), .C2(n2288), .A(n2597), 
        .ZN(n2590) );
  AOI22_X1 U3893 ( .A1(n2290), .A2(\pc_lut[6][13] ), .B1(n2291), .B2(
        \pc_lut[7][13] ), .ZN(n2597) );
  NAND2_X1 U3896 ( .A1(n2598), .A2(n2599), .ZN(N205) );
  NOR4_X1 U3897 ( .A1(n2600), .A2(n2601), .A3(n2602), .A4(n2603), .ZN(n2599)
         );
  OAI221_X1 U3898 ( .B1(n1420), .B2(n2248), .C1(n1386), .C2(n2249), .A(n2604), 
        .ZN(n2603) );
  AOI22_X1 U3899 ( .A1(n2251), .A2(\pc_lut[26][14] ), .B1(n2252), .B2(
        \pc_lut[27][14] ), .ZN(n2604) );
  OAI221_X1 U3902 ( .B1(n1285), .B2(n2253), .C1(n1250), .C2(n2254), .A(n2605), 
        .ZN(n2602) );
  AOI22_X1 U3903 ( .A1(n2256), .A2(\pc_lut[30][14] ), .B1(n2257), .B2(
        \pc_lut[31][14] ), .ZN(n2605) );
  OAI221_X1 U3906 ( .B1(n1684), .B2(n2258), .C1(n1650), .C2(n2259), .A(n2606), 
        .ZN(n2601) );
  AOI22_X1 U3907 ( .A1(n2261), .A2(\pc_lut[18][14] ), .B1(n2262), .B2(
        \pc_lut[19][14] ), .ZN(n2606) );
  OAI221_X1 U3910 ( .B1(n1489), .B2(n2263), .C1(n1454), .C2(n2264), .A(n2607), 
        .ZN(n2600) );
  AOI22_X1 U3911 ( .A1(n2266), .A2(\pc_lut[20][14] ), .B1(n2267), .B2(
        \pc_lut[21][14] ), .ZN(n2607) );
  NOR4_X1 U3914 ( .A1(n2608), .A2(n2609), .A3(n2610), .A4(n2611), .ZN(n2598)
         );
  OAI221_X1 U3915 ( .B1(n1954), .B2(n2272), .C1(n1920), .C2(n2273), .A(n2612), 
        .ZN(n2611) );
  AOI22_X1 U3916 ( .A1(n2275), .A2(\pc_lut[10][14] ), .B1(n2276), .B2(
        \pc_lut[11][14] ), .ZN(n2612) );
  OAI221_X1 U3919 ( .B1(n1819), .B2(n2277), .C1(n1785), .C2(n2278), .A(n2613), 
        .ZN(n2610) );
  AOI22_X1 U3920 ( .A1(n2280), .A2(\pc_lut[14][14] ), .B1(n2281), .B2(
        \pc_lut[15][14] ), .ZN(n2613) );
  OAI221_X1 U3923 ( .B1(n2218), .B2(n2282), .C1(n2184), .C2(n2283), .A(n2614), 
        .ZN(n2609) );
  AOI22_X1 U3924 ( .A1(n2285), .A2(\pc_lut[2][14] ), .B1(n2286), .B2(
        \pc_lut[3][14] ), .ZN(n2614) );
  OAI221_X1 U3927 ( .B1(n2086), .B2(n2287), .C1(n2052), .C2(n2288), .A(n2615), 
        .ZN(n2608) );
  AOI22_X1 U3928 ( .A1(n2290), .A2(\pc_lut[6][14] ), .B1(n2291), .B2(
        \pc_lut[7][14] ), .ZN(n2615) );
  NAND2_X1 U3931 ( .A1(n2616), .A2(n2617), .ZN(N204) );
  NOR4_X1 U3932 ( .A1(n2618), .A2(n2619), .A3(n2620), .A4(n2621), .ZN(n2617)
         );
  OAI221_X1 U3933 ( .B1(n1435), .B2(n2248), .C1(n1401), .C2(n2249), .A(n2622), 
        .ZN(n2621) );
  AOI22_X1 U3934 ( .A1(n2251), .A2(\pc_lut[26][15] ), .B1(n2252), .B2(
        \pc_lut[27][15] ), .ZN(n2622) );
  OAI221_X1 U3937 ( .B1(n1300), .B2(n2253), .C1(n1266), .C2(n2254), .A(n2623), 
        .ZN(n2620) );
  AOI22_X1 U3938 ( .A1(n2256), .A2(\pc_lut[30][15] ), .B1(n2257), .B2(
        \pc_lut[31][15] ), .ZN(n2623) );
  OAI221_X1 U3941 ( .B1(n1699), .B2(n2258), .C1(n1665), .C2(n2259), .A(n2624), 
        .ZN(n2619) );
  AOI22_X1 U3942 ( .A1(n2261), .A2(\pc_lut[18][15] ), .B1(n2262), .B2(
        \pc_lut[19][15] ), .ZN(n2624) );
  OAI221_X1 U3945 ( .B1(n1504), .B2(n2263), .C1(n1469), .C2(n2264), .A(n2625), 
        .ZN(n2618) );
  AOI22_X1 U3946 ( .A1(n2266), .A2(\pc_lut[20][15] ), .B1(n2267), .B2(
        \pc_lut[21][15] ), .ZN(n2625) );
  NOR4_X1 U3949 ( .A1(n2626), .A2(n2627), .A3(n2628), .A4(n2629), .ZN(n2616)
         );
  OAI221_X1 U3950 ( .B1(n1969), .B2(n2272), .C1(n1935), .C2(n2273), .A(n2630), 
        .ZN(n2629) );
  AOI22_X1 U3951 ( .A1(n2275), .A2(\pc_lut[10][15] ), .B1(n2276), .B2(
        \pc_lut[11][15] ), .ZN(n2630) );
  OAI221_X1 U3954 ( .B1(n1834), .B2(n2277), .C1(n1800), .C2(n2278), .A(n2631), 
        .ZN(n2628) );
  AOI22_X1 U3955 ( .A1(n2280), .A2(\pc_lut[14][15] ), .B1(n2281), .B2(
        \pc_lut[15][15] ), .ZN(n2631) );
  OAI221_X1 U3958 ( .B1(n2233), .B2(n2282), .C1(n2199), .C2(n2283), .A(n2632), 
        .ZN(n2627) );
  AOI22_X1 U3959 ( .A1(n2285), .A2(\pc_lut[2][15] ), .B1(n2286), .B2(
        \pc_lut[3][15] ), .ZN(n2632) );
  OAI221_X1 U3962 ( .B1(n2101), .B2(n2287), .C1(n2067), .C2(n2288), .A(n2633), 
        .ZN(n2626) );
  AOI22_X1 U3963 ( .A1(n2290), .A2(\pc_lut[6][15] ), .B1(n2291), .B2(
        \pc_lut[7][15] ), .ZN(n2633) );
  NAND2_X1 U3966 ( .A1(n2634), .A2(n2635), .ZN(N203) );
  NOR4_X1 U3967 ( .A1(n2636), .A2(n2637), .A3(n2638), .A4(n2639), .ZN(n2635)
         );
  OAI221_X1 U3968 ( .B1(n1419), .B2(n2248), .C1(n1385), .C2(n2249), .A(n2640), 
        .ZN(n2639) );
  AOI22_X1 U3969 ( .A1(n2251), .A2(\pc_lut[26][16] ), .B1(n2252), .B2(
        \pc_lut[27][16] ), .ZN(n2640) );
  OAI221_X1 U3972 ( .B1(n1284), .B2(n2253), .C1(n1249), .C2(n2254), .A(n2641), 
        .ZN(n2638) );
  AOI22_X1 U3973 ( .A1(n2256), .A2(\pc_lut[30][16] ), .B1(n2257), .B2(
        \pc_lut[31][16] ), .ZN(n2641) );
  OAI221_X1 U3976 ( .B1(n1683), .B2(n2258), .C1(n1649), .C2(n2259), .A(n2642), 
        .ZN(n2637) );
  AOI22_X1 U3977 ( .A1(n2261), .A2(\pc_lut[18][16] ), .B1(n2262), .B2(
        \pc_lut[19][16] ), .ZN(n2642) );
  OAI221_X1 U3980 ( .B1(n1488), .B2(n2263), .C1(n1453), .C2(n2264), .A(n2643), 
        .ZN(n2636) );
  AOI22_X1 U3981 ( .A1(n2266), .A2(\pc_lut[20][16] ), .B1(n2267), .B2(
        \pc_lut[21][16] ), .ZN(n2643) );
  NOR4_X1 U3984 ( .A1(n2644), .A2(n2645), .A3(n2646), .A4(n2647), .ZN(n2634)
         );
  OAI221_X1 U3985 ( .B1(n1953), .B2(n2272), .C1(n1919), .C2(n2273), .A(n2648), 
        .ZN(n2647) );
  AOI22_X1 U3986 ( .A1(n2275), .A2(\pc_lut[10][16] ), .B1(n2276), .B2(
        \pc_lut[11][16] ), .ZN(n2648) );
  OAI221_X1 U3989 ( .B1(n1818), .B2(n2277), .C1(n1784), .C2(n2278), .A(n2649), 
        .ZN(n2646) );
  AOI22_X1 U3990 ( .A1(n2280), .A2(\pc_lut[14][16] ), .B1(n2281), .B2(
        \pc_lut[15][16] ), .ZN(n2649) );
  OAI221_X1 U3993 ( .B1(n2217), .B2(n2282), .C1(n2183), .C2(n2283), .A(n2650), 
        .ZN(n2645) );
  AOI22_X1 U3994 ( .A1(n2285), .A2(\pc_lut[2][16] ), .B1(n2286), .B2(
        \pc_lut[3][16] ), .ZN(n2650) );
  OAI221_X1 U3997 ( .B1(n2085), .B2(n2287), .C1(n2051), .C2(n2288), .A(n2651), 
        .ZN(n2644) );
  AOI22_X1 U3998 ( .A1(n2290), .A2(\pc_lut[6][16] ), .B1(n2291), .B2(
        \pc_lut[7][16] ), .ZN(n2651) );
  NAND2_X1 U4001 ( .A1(n2652), .A2(n2653), .ZN(N202) );
  NOR4_X1 U4002 ( .A1(n2654), .A2(n2655), .A3(n2656), .A4(n2657), .ZN(n2653)
         );
  OAI221_X1 U4003 ( .B1(n1436), .B2(n2248), .C1(n1402), .C2(n2249), .A(n2658), 
        .ZN(n2657) );
  AOI22_X1 U4004 ( .A1(n2251), .A2(\pc_lut[26][17] ), .B1(n2252), .B2(
        \pc_lut[27][17] ), .ZN(n2658) );
  OAI221_X1 U4007 ( .B1(n1301), .B2(n2253), .C1(n1267), .C2(n2254), .A(n2659), 
        .ZN(n2656) );
  AOI22_X1 U4008 ( .A1(n2256), .A2(\pc_lut[30][17] ), .B1(n2257), .B2(
        \pc_lut[31][17] ), .ZN(n2659) );
  OAI221_X1 U4011 ( .B1(n1700), .B2(n2258), .C1(n1666), .C2(n2259), .A(n2660), 
        .ZN(n2655) );
  AOI22_X1 U4012 ( .A1(n2261), .A2(\pc_lut[18][17] ), .B1(n2262), .B2(
        \pc_lut[19][17] ), .ZN(n2660) );
  OAI221_X1 U4015 ( .B1(n1505), .B2(n2263), .C1(n1470), .C2(n2264), .A(n2661), 
        .ZN(n2654) );
  AOI22_X1 U4016 ( .A1(n2266), .A2(\pc_lut[20][17] ), .B1(n2267), .B2(
        \pc_lut[21][17] ), .ZN(n2661) );
  NOR4_X1 U4019 ( .A1(n2662), .A2(n2663), .A3(n2664), .A4(n2665), .ZN(n2652)
         );
  OAI221_X1 U4020 ( .B1(n1970), .B2(n2272), .C1(n1936), .C2(n2273), .A(n2666), 
        .ZN(n2665) );
  AOI22_X1 U4021 ( .A1(n2275), .A2(\pc_lut[10][17] ), .B1(n2276), .B2(
        \pc_lut[11][17] ), .ZN(n2666) );
  OAI221_X1 U4024 ( .B1(n1835), .B2(n2277), .C1(n1801), .C2(n2278), .A(n2667), 
        .ZN(n2664) );
  AOI22_X1 U4025 ( .A1(n2280), .A2(\pc_lut[14][17] ), .B1(n2281), .B2(
        \pc_lut[15][17] ), .ZN(n2667) );
  OAI221_X1 U4028 ( .B1(n2234), .B2(n2282), .C1(n2200), .C2(n2283), .A(n2668), 
        .ZN(n2663) );
  AOI22_X1 U4029 ( .A1(n2285), .A2(\pc_lut[2][17] ), .B1(n2286), .B2(
        \pc_lut[3][17] ), .ZN(n2668) );
  OAI221_X1 U4032 ( .B1(n2102), .B2(n2287), .C1(n2068), .C2(n2288), .A(n2669), 
        .ZN(n2662) );
  AOI22_X1 U4033 ( .A1(n2290), .A2(\pc_lut[6][17] ), .B1(n2291), .B2(
        \pc_lut[7][17] ), .ZN(n2669) );
  NAND2_X1 U4036 ( .A1(n2670), .A2(n2671), .ZN(N201) );
  NOR4_X1 U4037 ( .A1(n2672), .A2(n2673), .A3(n2674), .A4(n2675), .ZN(n2671)
         );
  OAI221_X1 U4038 ( .B1(n1418), .B2(n2248), .C1(n1384), .C2(n2249), .A(n2676), 
        .ZN(n2675) );
  AOI22_X1 U4039 ( .A1(n2251), .A2(\pc_lut[26][18] ), .B1(n2252), .B2(
        \pc_lut[27][18] ), .ZN(n2676) );
  OAI221_X1 U4042 ( .B1(n1283), .B2(n2253), .C1(n1248), .C2(n2254), .A(n2677), 
        .ZN(n2674) );
  AOI22_X1 U4043 ( .A1(n2256), .A2(\pc_lut[30][18] ), .B1(n2257), .B2(
        \pc_lut[31][18] ), .ZN(n2677) );
  OAI221_X1 U4046 ( .B1(n1682), .B2(n2258), .C1(n1648), .C2(n2259), .A(n2678), 
        .ZN(n2673) );
  AOI22_X1 U4047 ( .A1(n2261), .A2(\pc_lut[18][18] ), .B1(n2262), .B2(
        \pc_lut[19][18] ), .ZN(n2678) );
  OAI221_X1 U4050 ( .B1(n1487), .B2(n2263), .C1(n1452), .C2(n2264), .A(n2679), 
        .ZN(n2672) );
  AOI22_X1 U4051 ( .A1(n2266), .A2(\pc_lut[20][18] ), .B1(n2267), .B2(
        \pc_lut[21][18] ), .ZN(n2679) );
  NOR4_X1 U4054 ( .A1(n2680), .A2(n2681), .A3(n2682), .A4(n2683), .ZN(n2670)
         );
  OAI221_X1 U4055 ( .B1(n1952), .B2(n2272), .C1(n1918), .C2(n2273), .A(n2684), 
        .ZN(n2683) );
  AOI22_X1 U4056 ( .A1(n2275), .A2(\pc_lut[10][18] ), .B1(n2276), .B2(
        \pc_lut[11][18] ), .ZN(n2684) );
  OAI221_X1 U4059 ( .B1(n1817), .B2(n2277), .C1(n1783), .C2(n2278), .A(n2685), 
        .ZN(n2682) );
  AOI22_X1 U4060 ( .A1(n2280), .A2(\pc_lut[14][18] ), .B1(n2281), .B2(
        \pc_lut[15][18] ), .ZN(n2685) );
  OAI221_X1 U4063 ( .B1(n2216), .B2(n2282), .C1(n2182), .C2(n2283), .A(n2686), 
        .ZN(n2681) );
  AOI22_X1 U4064 ( .A1(n2285), .A2(\pc_lut[2][18] ), .B1(n2286), .B2(
        \pc_lut[3][18] ), .ZN(n2686) );
  OAI221_X1 U4067 ( .B1(n2084), .B2(n2287), .C1(n2050), .C2(n2288), .A(n2687), 
        .ZN(n2680) );
  AOI22_X1 U4068 ( .A1(n2290), .A2(\pc_lut[6][18] ), .B1(n2291), .B2(
        \pc_lut[7][18] ), .ZN(n2687) );
  NAND2_X1 U4071 ( .A1(n2688), .A2(n2689), .ZN(N200) );
  NOR4_X1 U4072 ( .A1(n2690), .A2(n2691), .A3(n2692), .A4(n2693), .ZN(n2689)
         );
  OAI221_X1 U4073 ( .B1(n1437), .B2(n2248), .C1(n1403), .C2(n2249), .A(n2694), 
        .ZN(n2693) );
  AOI22_X1 U4074 ( .A1(n2251), .A2(\pc_lut[26][19] ), .B1(n2252), .B2(
        \pc_lut[27][19] ), .ZN(n2694) );
  OAI221_X1 U4077 ( .B1(n1302), .B2(n2253), .C1(n1268), .C2(n2254), .A(n2695), 
        .ZN(n2692) );
  AOI22_X1 U4078 ( .A1(n2256), .A2(\pc_lut[30][19] ), .B1(n2257), .B2(
        \pc_lut[31][19] ), .ZN(n2695) );
  OAI221_X1 U4081 ( .B1(n1701), .B2(n2258), .C1(n1667), .C2(n2259), .A(n2696), 
        .ZN(n2691) );
  AOI22_X1 U4082 ( .A1(n2261), .A2(\pc_lut[18][19] ), .B1(n2262), .B2(
        \pc_lut[19][19] ), .ZN(n2696) );
  OAI221_X1 U4085 ( .B1(n1506), .B2(n2263), .C1(n1471), .C2(n2264), .A(n2697), 
        .ZN(n2690) );
  AOI22_X1 U4086 ( .A1(n2266), .A2(\pc_lut[20][19] ), .B1(n2267), .B2(
        \pc_lut[21][19] ), .ZN(n2697) );
  NOR4_X1 U4089 ( .A1(n2698), .A2(n2699), .A3(n2700), .A4(n2701), .ZN(n2688)
         );
  OAI221_X1 U4090 ( .B1(n1971), .B2(n2272), .C1(n1937), .C2(n2273), .A(n2702), 
        .ZN(n2701) );
  AOI22_X1 U4091 ( .A1(n2275), .A2(\pc_lut[10][19] ), .B1(n2276), .B2(
        \pc_lut[11][19] ), .ZN(n2702) );
  OAI221_X1 U4094 ( .B1(n1836), .B2(n2277), .C1(n1802), .C2(n2278), .A(n2703), 
        .ZN(n2700) );
  AOI22_X1 U4095 ( .A1(n2280), .A2(\pc_lut[14][19] ), .B1(n2281), .B2(
        \pc_lut[15][19] ), .ZN(n2703) );
  OAI221_X1 U4098 ( .B1(n2235), .B2(n2282), .C1(n2201), .C2(n2283), .A(n2704), 
        .ZN(n2699) );
  AOI22_X1 U4099 ( .A1(n2285), .A2(\pc_lut[2][19] ), .B1(n2286), .B2(
        \pc_lut[3][19] ), .ZN(n2704) );
  OAI221_X1 U4102 ( .B1(n2103), .B2(n2287), .C1(n2069), .C2(n2288), .A(n2705), 
        .ZN(n2698) );
  AOI22_X1 U4103 ( .A1(n2290), .A2(\pc_lut[6][19] ), .B1(n2291), .B2(
        \pc_lut[7][19] ), .ZN(n2705) );
  NAND2_X1 U4106 ( .A1(n2706), .A2(n2707), .ZN(N199) );
  NOR4_X1 U4107 ( .A1(n2708), .A2(n2709), .A3(n2710), .A4(n2711), .ZN(n2707)
         );
  OAI221_X1 U4108 ( .B1(n1417), .B2(n2248), .C1(n1383), .C2(n2249), .A(n2712), 
        .ZN(n2711) );
  AOI22_X1 U4109 ( .A1(n2251), .A2(\pc_lut[26][20] ), .B1(n2252), .B2(
        \pc_lut[27][20] ), .ZN(n2712) );
  OAI221_X1 U4112 ( .B1(n1282), .B2(n2253), .C1(n1247), .C2(n2254), .A(n2713), 
        .ZN(n2710) );
  AOI22_X1 U4113 ( .A1(n2256), .A2(\pc_lut[30][20] ), .B1(n2257), .B2(
        \pc_lut[31][20] ), .ZN(n2713) );
  OAI221_X1 U4116 ( .B1(n1681), .B2(n2258), .C1(n1647), .C2(n2259), .A(n2714), 
        .ZN(n2709) );
  AOI22_X1 U4117 ( .A1(n2261), .A2(\pc_lut[18][20] ), .B1(n2262), .B2(
        \pc_lut[19][20] ), .ZN(n2714) );
  OAI221_X1 U4120 ( .B1(n1486), .B2(n2263), .C1(n1451), .C2(n2264), .A(n2715), 
        .ZN(n2708) );
  AOI22_X1 U4121 ( .A1(n2266), .A2(\pc_lut[20][20] ), .B1(n2267), .B2(
        \pc_lut[21][20] ), .ZN(n2715) );
  NOR4_X1 U4124 ( .A1(n2716), .A2(n2717), .A3(n2718), .A4(n2719), .ZN(n2706)
         );
  OAI221_X1 U4125 ( .B1(n1951), .B2(n2272), .C1(n1917), .C2(n2273), .A(n2720), 
        .ZN(n2719) );
  AOI22_X1 U4126 ( .A1(n2275), .A2(\pc_lut[10][20] ), .B1(n2276), .B2(
        \pc_lut[11][20] ), .ZN(n2720) );
  OAI221_X1 U4129 ( .B1(n1816), .B2(n2277), .C1(n1782), .C2(n2278), .A(n2721), 
        .ZN(n2718) );
  AOI22_X1 U4130 ( .A1(n2280), .A2(\pc_lut[14][20] ), .B1(n2281), .B2(
        \pc_lut[15][20] ), .ZN(n2721) );
  OAI221_X1 U4133 ( .B1(n2215), .B2(n2282), .C1(n2181), .C2(n2283), .A(n2722), 
        .ZN(n2717) );
  AOI22_X1 U4134 ( .A1(n2285), .A2(\pc_lut[2][20] ), .B1(n2286), .B2(
        \pc_lut[3][20] ), .ZN(n2722) );
  OAI221_X1 U4137 ( .B1(n2083), .B2(n2287), .C1(n2049), .C2(n2288), .A(n2723), 
        .ZN(n2716) );
  AOI22_X1 U4138 ( .A1(n2290), .A2(\pc_lut[6][20] ), .B1(n2291), .B2(
        \pc_lut[7][20] ), .ZN(n2723) );
  NAND2_X1 U4141 ( .A1(n2724), .A2(n2725), .ZN(N198) );
  NOR4_X1 U4142 ( .A1(n2726), .A2(n2727), .A3(n2728), .A4(n2729), .ZN(n2725)
         );
  OAI221_X1 U4143 ( .B1(n1438), .B2(n2248), .C1(n1404), .C2(n2249), .A(n2730), 
        .ZN(n2729) );
  AOI22_X1 U4144 ( .A1(n2251), .A2(\pc_lut[26][21] ), .B1(n2252), .B2(
        \pc_lut[27][21] ), .ZN(n2730) );
  OAI221_X1 U4147 ( .B1(n1303), .B2(n2253), .C1(n1269), .C2(n2254), .A(n2731), 
        .ZN(n2728) );
  AOI22_X1 U4148 ( .A1(n2256), .A2(\pc_lut[30][21] ), .B1(n2257), .B2(
        \pc_lut[31][21] ), .ZN(n2731) );
  OAI221_X1 U4151 ( .B1(n1702), .B2(n2258), .C1(n1668), .C2(n2259), .A(n2732), 
        .ZN(n2727) );
  AOI22_X1 U4152 ( .A1(n2261), .A2(\pc_lut[18][21] ), .B1(n2262), .B2(
        \pc_lut[19][21] ), .ZN(n2732) );
  OAI221_X1 U4155 ( .B1(n1507), .B2(n2263), .C1(n1472), .C2(n2264), .A(n2733), 
        .ZN(n2726) );
  AOI22_X1 U4156 ( .A1(n2266), .A2(\pc_lut[20][21] ), .B1(n2267), .B2(
        \pc_lut[21][21] ), .ZN(n2733) );
  NOR4_X1 U4159 ( .A1(n2734), .A2(n2735), .A3(n2736), .A4(n2737), .ZN(n2724)
         );
  OAI221_X1 U4160 ( .B1(n1972), .B2(n2272), .C1(n1938), .C2(n2273), .A(n2738), 
        .ZN(n2737) );
  AOI22_X1 U4161 ( .A1(n2275), .A2(\pc_lut[10][21] ), .B1(n2276), .B2(
        \pc_lut[11][21] ), .ZN(n2738) );
  OAI221_X1 U4164 ( .B1(n1837), .B2(n2277), .C1(n1803), .C2(n2278), .A(n2739), 
        .ZN(n2736) );
  AOI22_X1 U4165 ( .A1(n2280), .A2(\pc_lut[14][21] ), .B1(n2281), .B2(
        \pc_lut[15][21] ), .ZN(n2739) );
  OAI221_X1 U4168 ( .B1(n2236), .B2(n2282), .C1(n2202), .C2(n2283), .A(n2740), 
        .ZN(n2735) );
  AOI22_X1 U4169 ( .A1(n2285), .A2(\pc_lut[2][21] ), .B1(n2286), .B2(
        \pc_lut[3][21] ), .ZN(n2740) );
  OAI221_X1 U4172 ( .B1(n2104), .B2(n2287), .C1(n2070), .C2(n2288), .A(n2741), 
        .ZN(n2734) );
  AOI22_X1 U4173 ( .A1(n2290), .A2(\pc_lut[6][21] ), .B1(n2291), .B2(
        \pc_lut[7][21] ), .ZN(n2741) );
  NAND2_X1 U4176 ( .A1(n2742), .A2(n2743), .ZN(N197) );
  NOR4_X1 U4177 ( .A1(n2744), .A2(n2745), .A3(n2746), .A4(n2747), .ZN(n2743)
         );
  OAI221_X1 U4178 ( .B1(n1416), .B2(n2248), .C1(n1382), .C2(n2249), .A(n2748), 
        .ZN(n2747) );
  AOI22_X1 U4179 ( .A1(n2251), .A2(\pc_lut[26][22] ), .B1(n2252), .B2(
        \pc_lut[27][22] ), .ZN(n2748) );
  OAI221_X1 U4182 ( .B1(n1281), .B2(n2253), .C1(n1246), .C2(n2254), .A(n2749), 
        .ZN(n2746) );
  AOI22_X1 U4183 ( .A1(n2256), .A2(\pc_lut[30][22] ), .B1(n2257), .B2(
        \pc_lut[31][22] ), .ZN(n2749) );
  OAI221_X1 U4186 ( .B1(n1680), .B2(n2258), .C1(n1646), .C2(n2259), .A(n2750), 
        .ZN(n2745) );
  AOI22_X1 U4187 ( .A1(n2261), .A2(\pc_lut[18][22] ), .B1(n2262), .B2(
        \pc_lut[19][22] ), .ZN(n2750) );
  OAI221_X1 U4190 ( .B1(n1485), .B2(n2263), .C1(n1450), .C2(n2264), .A(n2751), 
        .ZN(n2744) );
  AOI22_X1 U4191 ( .A1(n2266), .A2(\pc_lut[20][22] ), .B1(n2267), .B2(
        \pc_lut[21][22] ), .ZN(n2751) );
  NOR4_X1 U4194 ( .A1(n2752), .A2(n2753), .A3(n2754), .A4(n2755), .ZN(n2742)
         );
  OAI221_X1 U4195 ( .B1(n1950), .B2(n2272), .C1(n1916), .C2(n2273), .A(n2756), 
        .ZN(n2755) );
  AOI22_X1 U4196 ( .A1(n2275), .A2(\pc_lut[10][22] ), .B1(n2276), .B2(
        \pc_lut[11][22] ), .ZN(n2756) );
  OAI221_X1 U4199 ( .B1(n1815), .B2(n2277), .C1(n1781), .C2(n2278), .A(n2757), 
        .ZN(n2754) );
  AOI22_X1 U4200 ( .A1(n2280), .A2(\pc_lut[14][22] ), .B1(n2281), .B2(
        \pc_lut[15][22] ), .ZN(n2757) );
  OAI221_X1 U4203 ( .B1(n2214), .B2(n2282), .C1(n2180), .C2(n2283), .A(n2758), 
        .ZN(n2753) );
  AOI22_X1 U4204 ( .A1(n2285), .A2(\pc_lut[2][22] ), .B1(n2286), .B2(
        \pc_lut[3][22] ), .ZN(n2758) );
  OAI221_X1 U4207 ( .B1(n2082), .B2(n2287), .C1(n2048), .C2(n2288), .A(n2759), 
        .ZN(n2752) );
  AOI22_X1 U4208 ( .A1(n2290), .A2(\pc_lut[6][22] ), .B1(n2291), .B2(
        \pc_lut[7][22] ), .ZN(n2759) );
  NAND2_X1 U4211 ( .A1(n2760), .A2(n2761), .ZN(N196) );
  NOR4_X1 U4212 ( .A1(n2762), .A2(n2763), .A3(n2764), .A4(n2765), .ZN(n2761)
         );
  OAI221_X1 U4213 ( .B1(n1439), .B2(n2248), .C1(n1405), .C2(n2249), .A(n2766), 
        .ZN(n2765) );
  AOI22_X1 U4214 ( .A1(n2251), .A2(\pc_lut[26][23] ), .B1(n2252), .B2(
        \pc_lut[27][23] ), .ZN(n2766) );
  OAI221_X1 U4217 ( .B1(n1304), .B2(n2253), .C1(n1270), .C2(n2254), .A(n2767), 
        .ZN(n2764) );
  AOI22_X1 U4218 ( .A1(n2256), .A2(\pc_lut[30][23] ), .B1(n2257), .B2(
        \pc_lut[31][23] ), .ZN(n2767) );
  OAI221_X1 U4221 ( .B1(n1703), .B2(n2258), .C1(n1669), .C2(n2259), .A(n2768), 
        .ZN(n2763) );
  AOI22_X1 U4222 ( .A1(n2261), .A2(\pc_lut[18][23] ), .B1(n2262), .B2(
        \pc_lut[19][23] ), .ZN(n2768) );
  OAI221_X1 U4225 ( .B1(n1508), .B2(n2263), .C1(n1473), .C2(n2264), .A(n2769), 
        .ZN(n2762) );
  AOI22_X1 U4226 ( .A1(n2266), .A2(\pc_lut[20][23] ), .B1(n2267), .B2(
        \pc_lut[21][23] ), .ZN(n2769) );
  NOR4_X1 U4229 ( .A1(n2770), .A2(n2771), .A3(n2772), .A4(n2773), .ZN(n2760)
         );
  OAI221_X1 U4230 ( .B1(n1973), .B2(n2272), .C1(n1939), .C2(n2273), .A(n2774), 
        .ZN(n2773) );
  AOI22_X1 U4231 ( .A1(n2275), .A2(\pc_lut[10][23] ), .B1(n2276), .B2(
        \pc_lut[11][23] ), .ZN(n2774) );
  OAI221_X1 U4234 ( .B1(n1838), .B2(n2277), .C1(n1804), .C2(n2278), .A(n2775), 
        .ZN(n2772) );
  AOI22_X1 U4235 ( .A1(n2280), .A2(\pc_lut[14][23] ), .B1(n2281), .B2(
        \pc_lut[15][23] ), .ZN(n2775) );
  OAI221_X1 U4238 ( .B1(n2237), .B2(n2282), .C1(n2203), .C2(n2283), .A(n2776), 
        .ZN(n2771) );
  AOI22_X1 U4239 ( .A1(n2285), .A2(\pc_lut[2][23] ), .B1(n2286), .B2(
        \pc_lut[3][23] ), .ZN(n2776) );
  OAI221_X1 U4242 ( .B1(n2105), .B2(n2287), .C1(n2071), .C2(n2288), .A(n2777), 
        .ZN(n2770) );
  AOI22_X1 U4243 ( .A1(n2290), .A2(\pc_lut[6][23] ), .B1(n2291), .B2(
        \pc_lut[7][23] ), .ZN(n2777) );
  NAND2_X1 U4246 ( .A1(n2778), .A2(n2779), .ZN(N195) );
  NOR4_X1 U4247 ( .A1(n2780), .A2(n2781), .A3(n2782), .A4(n2783), .ZN(n2779)
         );
  OAI221_X1 U4248 ( .B1(n1415), .B2(n2248), .C1(n1381), .C2(n2249), .A(n2784), 
        .ZN(n2783) );
  AOI22_X1 U4249 ( .A1(n2251), .A2(\pc_lut[26][24] ), .B1(n2252), .B2(
        \pc_lut[27][24] ), .ZN(n2784) );
  OAI221_X1 U4252 ( .B1(n1280), .B2(n2253), .C1(n1245), .C2(n2254), .A(n2785), 
        .ZN(n2782) );
  AOI22_X1 U4253 ( .A1(n2256), .A2(\pc_lut[30][24] ), .B1(n2257), .B2(
        \pc_lut[31][24] ), .ZN(n2785) );
  OAI221_X1 U4256 ( .B1(n1679), .B2(n2258), .C1(n1645), .C2(n2259), .A(n2786), 
        .ZN(n2781) );
  AOI22_X1 U4257 ( .A1(n2261), .A2(\pc_lut[18][24] ), .B1(n2262), .B2(
        \pc_lut[19][24] ), .ZN(n2786) );
  OAI221_X1 U4260 ( .B1(n1484), .B2(n2263), .C1(n1449), .C2(n2264), .A(n2787), 
        .ZN(n2780) );
  AOI22_X1 U4261 ( .A1(n2266), .A2(\pc_lut[20][24] ), .B1(n2267), .B2(
        \pc_lut[21][24] ), .ZN(n2787) );
  NOR4_X1 U4264 ( .A1(n2788), .A2(n2789), .A3(n2790), .A4(n2791), .ZN(n2778)
         );
  OAI221_X1 U4265 ( .B1(n1949), .B2(n2272), .C1(n1915), .C2(n2273), .A(n2792), 
        .ZN(n2791) );
  AOI22_X1 U4266 ( .A1(n2275), .A2(\pc_lut[10][24] ), .B1(n2276), .B2(
        \pc_lut[11][24] ), .ZN(n2792) );
  OAI221_X1 U4269 ( .B1(n1814), .B2(n2277), .C1(n1780), .C2(n2278), .A(n2793), 
        .ZN(n2790) );
  AOI22_X1 U4270 ( .A1(n2280), .A2(\pc_lut[14][24] ), .B1(n2281), .B2(
        \pc_lut[15][24] ), .ZN(n2793) );
  OAI221_X1 U4273 ( .B1(n2213), .B2(n2282), .C1(n2179), .C2(n2283), .A(n2794), 
        .ZN(n2789) );
  AOI22_X1 U4274 ( .A1(n2285), .A2(\pc_lut[2][24] ), .B1(n2286), .B2(
        \pc_lut[3][24] ), .ZN(n2794) );
  OAI221_X1 U4277 ( .B1(n2081), .B2(n2287), .C1(n2047), .C2(n2288), .A(n2795), 
        .ZN(n2788) );
  AOI22_X1 U4278 ( .A1(n2290), .A2(\pc_lut[6][24] ), .B1(n2291), .B2(
        \pc_lut[7][24] ), .ZN(n2795) );
  NAND2_X1 U4281 ( .A1(n2796), .A2(n2797), .ZN(N194) );
  NOR4_X1 U4282 ( .A1(n2798), .A2(n2799), .A3(n2800), .A4(n2801), .ZN(n2797)
         );
  OAI221_X1 U4283 ( .B1(n1440), .B2(n2248), .C1(n1406), .C2(n2249), .A(n2802), 
        .ZN(n2801) );
  AOI22_X1 U4284 ( .A1(n2251), .A2(\pc_lut[26][25] ), .B1(n2252), .B2(
        \pc_lut[27][25] ), .ZN(n2802) );
  OAI221_X1 U4287 ( .B1(n1305), .B2(n2253), .C1(n1271), .C2(n2254), .A(n2803), 
        .ZN(n2800) );
  AOI22_X1 U4288 ( .A1(n2256), .A2(\pc_lut[30][25] ), .B1(n2257), .B2(
        \pc_lut[31][25] ), .ZN(n2803) );
  OAI221_X1 U4291 ( .B1(n1704), .B2(n2258), .C1(n1670), .C2(n2259), .A(n2804), 
        .ZN(n2799) );
  AOI22_X1 U4292 ( .A1(n2261), .A2(\pc_lut[18][25] ), .B1(n2262), .B2(
        \pc_lut[19][25] ), .ZN(n2804) );
  OAI221_X1 U4295 ( .B1(n1509), .B2(n2263), .C1(n1474), .C2(n2264), .A(n2805), 
        .ZN(n2798) );
  AOI22_X1 U4296 ( .A1(n2266), .A2(\pc_lut[20][25] ), .B1(n2267), .B2(
        \pc_lut[21][25] ), .ZN(n2805) );
  NOR4_X1 U4299 ( .A1(n2806), .A2(n2807), .A3(n2808), .A4(n2809), .ZN(n2796)
         );
  OAI221_X1 U4300 ( .B1(n1974), .B2(n2272), .C1(n1940), .C2(n2273), .A(n2810), 
        .ZN(n2809) );
  AOI22_X1 U4301 ( .A1(n2275), .A2(\pc_lut[10][25] ), .B1(n2276), .B2(
        \pc_lut[11][25] ), .ZN(n2810) );
  OAI221_X1 U4304 ( .B1(n1839), .B2(n2277), .C1(n1805), .C2(n2278), .A(n2811), 
        .ZN(n2808) );
  AOI22_X1 U4305 ( .A1(n2280), .A2(\pc_lut[14][25] ), .B1(n2281), .B2(
        \pc_lut[15][25] ), .ZN(n2811) );
  OAI221_X1 U4308 ( .B1(n2238), .B2(n2282), .C1(n2204), .C2(n2283), .A(n2812), 
        .ZN(n2807) );
  AOI22_X1 U4309 ( .A1(n2285), .A2(\pc_lut[2][25] ), .B1(n2286), .B2(
        \pc_lut[3][25] ), .ZN(n2812) );
  OAI221_X1 U4312 ( .B1(n2106), .B2(n2287), .C1(n2072), .C2(n2288), .A(n2813), 
        .ZN(n2806) );
  AOI22_X1 U4313 ( .A1(n2290), .A2(\pc_lut[6][25] ), .B1(n2291), .B2(
        \pc_lut[7][25] ), .ZN(n2813) );
  NAND2_X1 U4316 ( .A1(n2814), .A2(n2815), .ZN(N193) );
  NOR4_X1 U4317 ( .A1(n2816), .A2(n2817), .A3(n2818), .A4(n2819), .ZN(n2815)
         );
  OAI221_X1 U4318 ( .B1(n1414), .B2(n2248), .C1(n1380), .C2(n2249), .A(n2820), 
        .ZN(n2819) );
  AOI22_X1 U4319 ( .A1(n2251), .A2(\pc_lut[26][26] ), .B1(n2252), .B2(
        \pc_lut[27][26] ), .ZN(n2820) );
  OAI221_X1 U4322 ( .B1(n1279), .B2(n2253), .C1(n1244), .C2(n2254), .A(n2821), 
        .ZN(n2818) );
  AOI22_X1 U4323 ( .A1(n2256), .A2(\pc_lut[30][26] ), .B1(n2257), .B2(
        \pc_lut[31][26] ), .ZN(n2821) );
  OAI221_X1 U4326 ( .B1(n1678), .B2(n2258), .C1(n1644), .C2(n2259), .A(n2822), 
        .ZN(n2817) );
  AOI22_X1 U4327 ( .A1(n2261), .A2(\pc_lut[18][26] ), .B1(n2262), .B2(
        \pc_lut[19][26] ), .ZN(n2822) );
  OAI221_X1 U4330 ( .B1(n1483), .B2(n2263), .C1(n1448), .C2(n2264), .A(n2823), 
        .ZN(n2816) );
  AOI22_X1 U4331 ( .A1(n2266), .A2(\pc_lut[20][26] ), .B1(n2267), .B2(
        \pc_lut[21][26] ), .ZN(n2823) );
  NOR4_X1 U4334 ( .A1(n2824), .A2(n2825), .A3(n2826), .A4(n2827), .ZN(n2814)
         );
  OAI221_X1 U4335 ( .B1(n1948), .B2(n2272), .C1(n1914), .C2(n2273), .A(n2828), 
        .ZN(n2827) );
  AOI22_X1 U4336 ( .A1(n2275), .A2(\pc_lut[10][26] ), .B1(n2276), .B2(
        \pc_lut[11][26] ), .ZN(n2828) );
  OAI221_X1 U4339 ( .B1(n1813), .B2(n2277), .C1(n1779), .C2(n2278), .A(n2829), 
        .ZN(n2826) );
  AOI22_X1 U4340 ( .A1(n2280), .A2(\pc_lut[14][26] ), .B1(n2281), .B2(
        \pc_lut[15][26] ), .ZN(n2829) );
  OAI221_X1 U4343 ( .B1(n2212), .B2(n2282), .C1(n2178), .C2(n2283), .A(n2830), 
        .ZN(n2825) );
  AOI22_X1 U4344 ( .A1(n2285), .A2(\pc_lut[2][26] ), .B1(n2286), .B2(
        \pc_lut[3][26] ), .ZN(n2830) );
  OAI221_X1 U4347 ( .B1(n2080), .B2(n2287), .C1(n2046), .C2(n2288), .A(n2831), 
        .ZN(n2824) );
  AOI22_X1 U4348 ( .A1(n2290), .A2(\pc_lut[6][26] ), .B1(n2291), .B2(
        \pc_lut[7][26] ), .ZN(n2831) );
  NAND2_X1 U4351 ( .A1(n2832), .A2(n2833), .ZN(N192) );
  NOR4_X1 U4352 ( .A1(n2834), .A2(n2835), .A3(n2836), .A4(n2837), .ZN(n2833)
         );
  OAI221_X1 U4353 ( .B1(n1441), .B2(n2248), .C1(n1407), .C2(n2249), .A(n2838), 
        .ZN(n2837) );
  AOI22_X1 U4354 ( .A1(n2251), .A2(\pc_lut[26][27] ), .B1(n2252), .B2(
        \pc_lut[27][27] ), .ZN(n2838) );
  OAI221_X1 U4357 ( .B1(n1306), .B2(n2253), .C1(n1272), .C2(n2254), .A(n2839), 
        .ZN(n2836) );
  AOI22_X1 U4358 ( .A1(n2256), .A2(\pc_lut[30][27] ), .B1(n2257), .B2(
        \pc_lut[31][27] ), .ZN(n2839) );
  OAI221_X1 U4361 ( .B1(n1705), .B2(n2258), .C1(n1671), .C2(n2259), .A(n2840), 
        .ZN(n2835) );
  AOI22_X1 U4362 ( .A1(n2261), .A2(\pc_lut[18][27] ), .B1(n2262), .B2(
        \pc_lut[19][27] ), .ZN(n2840) );
  OAI221_X1 U4365 ( .B1(n1510), .B2(n2263), .C1(n1475), .C2(n2264), .A(n2841), 
        .ZN(n2834) );
  AOI22_X1 U4366 ( .A1(n2266), .A2(\pc_lut[20][27] ), .B1(n2267), .B2(
        \pc_lut[21][27] ), .ZN(n2841) );
  NOR4_X1 U4369 ( .A1(n2842), .A2(n2843), .A3(n2844), .A4(n2845), .ZN(n2832)
         );
  OAI221_X1 U4370 ( .B1(n1975), .B2(n2272), .C1(n1941), .C2(n2273), .A(n2846), 
        .ZN(n2845) );
  AOI22_X1 U4371 ( .A1(n2275), .A2(\pc_lut[10][27] ), .B1(n2276), .B2(
        \pc_lut[11][27] ), .ZN(n2846) );
  OAI221_X1 U4374 ( .B1(n1840), .B2(n2277), .C1(n1806), .C2(n2278), .A(n2847), 
        .ZN(n2844) );
  AOI22_X1 U4375 ( .A1(n2280), .A2(\pc_lut[14][27] ), .B1(n2281), .B2(
        \pc_lut[15][27] ), .ZN(n2847) );
  OAI221_X1 U4378 ( .B1(n2239), .B2(n2282), .C1(n2205), .C2(n2283), .A(n2848), 
        .ZN(n2843) );
  AOI22_X1 U4379 ( .A1(n2285), .A2(\pc_lut[2][27] ), .B1(n2286), .B2(
        \pc_lut[3][27] ), .ZN(n2848) );
  OAI221_X1 U4382 ( .B1(n2107), .B2(n2287), .C1(n2073), .C2(n2288), .A(n2849), 
        .ZN(n2842) );
  AOI22_X1 U4383 ( .A1(n2290), .A2(\pc_lut[6][27] ), .B1(n2291), .B2(
        \pc_lut[7][27] ), .ZN(n2849) );
  NAND2_X1 U4386 ( .A1(n2850), .A2(n2851), .ZN(N191) );
  NOR4_X1 U4387 ( .A1(n2852), .A2(n2853), .A3(n2854), .A4(n2855), .ZN(n2851)
         );
  OAI221_X1 U4388 ( .B1(n1413), .B2(n2248), .C1(n1379), .C2(n2249), .A(n2856), 
        .ZN(n2855) );
  AOI22_X1 U4389 ( .A1(n2251), .A2(\pc_lut[26][28] ), .B1(n2252), .B2(
        \pc_lut[27][28] ), .ZN(n2856) );
  OAI221_X1 U4392 ( .B1(n1278), .B2(n2253), .C1(n1243), .C2(n2254), .A(n2857), 
        .ZN(n2854) );
  AOI22_X1 U4393 ( .A1(n2256), .A2(\pc_lut[30][28] ), .B1(n2257), .B2(
        \pc_lut[31][28] ), .ZN(n2857) );
  OAI221_X1 U4396 ( .B1(n1677), .B2(n2258), .C1(n1643), .C2(n2259), .A(n2858), 
        .ZN(n2853) );
  AOI22_X1 U4397 ( .A1(n2261), .A2(\pc_lut[18][28] ), .B1(n2262), .B2(
        \pc_lut[19][28] ), .ZN(n2858) );
  OAI221_X1 U4400 ( .B1(n1482), .B2(n2263), .C1(n1447), .C2(n2264), .A(n2859), 
        .ZN(n2852) );
  AOI22_X1 U4401 ( .A1(n2266), .A2(\pc_lut[20][28] ), .B1(n2267), .B2(
        \pc_lut[21][28] ), .ZN(n2859) );
  NOR4_X1 U4404 ( .A1(n2860), .A2(n2861), .A3(n2862), .A4(n2863), .ZN(n2850)
         );
  OAI221_X1 U4405 ( .B1(n1947), .B2(n2272), .C1(n1913), .C2(n2273), .A(n2864), 
        .ZN(n2863) );
  AOI22_X1 U4406 ( .A1(n2275), .A2(\pc_lut[10][28] ), .B1(n2276), .B2(
        \pc_lut[11][28] ), .ZN(n2864) );
  OAI221_X1 U4409 ( .B1(n1812), .B2(n2277), .C1(n1778), .C2(n2278), .A(n2865), 
        .ZN(n2862) );
  AOI22_X1 U4410 ( .A1(n2280), .A2(\pc_lut[14][28] ), .B1(n2281), .B2(
        \pc_lut[15][28] ), .ZN(n2865) );
  OAI221_X1 U4413 ( .B1(n2211), .B2(n2282), .C1(n2177), .C2(n2283), .A(n2866), 
        .ZN(n2861) );
  AOI22_X1 U4414 ( .A1(n2285), .A2(\pc_lut[2][28] ), .B1(n2286), .B2(
        \pc_lut[3][28] ), .ZN(n2866) );
  OAI221_X1 U4417 ( .B1(n2079), .B2(n2287), .C1(n2045), .C2(n2288), .A(n2867), 
        .ZN(n2860) );
  AOI22_X1 U4418 ( .A1(n2290), .A2(\pc_lut[6][28] ), .B1(n2291), .B2(
        \pc_lut[7][28] ), .ZN(n2867) );
  NAND2_X1 U4421 ( .A1(n2868), .A2(n2869), .ZN(N190) );
  NOR4_X1 U4422 ( .A1(n2870), .A2(n2871), .A3(n2872), .A4(n2873), .ZN(n2869)
         );
  OAI221_X1 U4423 ( .B1(n1442), .B2(n2248), .C1(n1408), .C2(n2249), .A(n2874), 
        .ZN(n2873) );
  AOI22_X1 U4424 ( .A1(n2251), .A2(\pc_lut[26][29] ), .B1(n2252), .B2(
        \pc_lut[27][29] ), .ZN(n2874) );
  OAI221_X1 U4427 ( .B1(n1307), .B2(n2253), .C1(n1273), .C2(n2254), .A(n2875), 
        .ZN(n2872) );
  AOI22_X1 U4428 ( .A1(n2256), .A2(\pc_lut[30][29] ), .B1(n2257), .B2(
        \pc_lut[31][29] ), .ZN(n2875) );
  OAI221_X1 U4431 ( .B1(n1706), .B2(n2258), .C1(n1672), .C2(n2259), .A(n2876), 
        .ZN(n2871) );
  AOI22_X1 U4432 ( .A1(n2261), .A2(\pc_lut[18][29] ), .B1(n2262), .B2(
        \pc_lut[19][29] ), .ZN(n2876) );
  OAI221_X1 U4435 ( .B1(n1511), .B2(n2263), .C1(n1476), .C2(n2264), .A(n2877), 
        .ZN(n2870) );
  AOI22_X1 U4436 ( .A1(n2266), .A2(\pc_lut[20][29] ), .B1(n2267), .B2(
        \pc_lut[21][29] ), .ZN(n2877) );
  NOR4_X1 U4439 ( .A1(n2878), .A2(n2879), .A3(n2880), .A4(n2881), .ZN(n2868)
         );
  OAI221_X1 U4440 ( .B1(n1976), .B2(n2272), .C1(n1942), .C2(n2273), .A(n2882), 
        .ZN(n2881) );
  AOI22_X1 U4441 ( .A1(n2275), .A2(\pc_lut[10][29] ), .B1(n2276), .B2(
        \pc_lut[11][29] ), .ZN(n2882) );
  OAI221_X1 U4444 ( .B1(n1841), .B2(n2277), .C1(n1807), .C2(n2278), .A(n2883), 
        .ZN(n2880) );
  AOI22_X1 U4445 ( .A1(n2280), .A2(\pc_lut[14][29] ), .B1(n2281), .B2(
        \pc_lut[15][29] ), .ZN(n2883) );
  OAI221_X1 U4448 ( .B1(n2240), .B2(n2282), .C1(n2206), .C2(n2283), .A(n2884), 
        .ZN(n2879) );
  AOI22_X1 U4449 ( .A1(n2285), .A2(\pc_lut[2][29] ), .B1(n2286), .B2(
        \pc_lut[3][29] ), .ZN(n2884) );
  OAI221_X1 U4452 ( .B1(n2108), .B2(n2287), .C1(n2074), .C2(n2288), .A(n2885), 
        .ZN(n2878) );
  AOI22_X1 U4453 ( .A1(n2290), .A2(\pc_lut[6][29] ), .B1(n2291), .B2(
        \pc_lut[7][29] ), .ZN(n2885) );
  NAND2_X1 U4456 ( .A1(n2886), .A2(n2887), .ZN(N189) );
  NOR4_X1 U4457 ( .A1(n2888), .A2(n2889), .A3(n2890), .A4(n2891), .ZN(n2887)
         );
  OAI221_X1 U4458 ( .B1(n1411), .B2(n2248), .C1(n1377), .C2(n2249), .A(n2892), 
        .ZN(n2891) );
  AOI22_X1 U4459 ( .A1(n2251), .A2(\pc_lut[26][30] ), .B1(n2252), .B2(
        \pc_lut[27][30] ), .ZN(n2892) );
  OAI221_X1 U4462 ( .B1(n1276), .B2(n2253), .C1(n1241), .C2(n2254), .A(n2893), 
        .ZN(n2890) );
  AOI22_X1 U4463 ( .A1(n2256), .A2(\pc_lut[30][30] ), .B1(n2257), .B2(
        \pc_lut[31][30] ), .ZN(n2893) );
  OAI221_X1 U4466 ( .B1(n1675), .B2(n2258), .C1(n1641), .C2(n2259), .A(n2894), 
        .ZN(n2889) );
  AOI22_X1 U4467 ( .A1(n2261), .A2(\pc_lut[18][30] ), .B1(n2262), .B2(
        \pc_lut[19][30] ), .ZN(n2894) );
  OAI221_X1 U4470 ( .B1(n1480), .B2(n2263), .C1(n1445), .C2(n2264), .A(n2895), 
        .ZN(n2888) );
  AOI22_X1 U4471 ( .A1(n2266), .A2(\pc_lut[20][30] ), .B1(n2267), .B2(
        \pc_lut[21][30] ), .ZN(n2895) );
  NOR4_X1 U4474 ( .A1(n2896), .A2(n2897), .A3(n2898), .A4(n2899), .ZN(n2886)
         );
  OAI221_X1 U4475 ( .B1(n1945), .B2(n2272), .C1(n1911), .C2(n2273), .A(n2900), 
        .ZN(n2899) );
  AOI22_X1 U4476 ( .A1(n2275), .A2(\pc_lut[10][30] ), .B1(n2276), .B2(
        \pc_lut[11][30] ), .ZN(n2900) );
  OAI221_X1 U4479 ( .B1(n1810), .B2(n2277), .C1(n1776), .C2(n2278), .A(n2901), 
        .ZN(n2898) );
  AOI22_X1 U4480 ( .A1(n2280), .A2(\pc_lut[14][30] ), .B1(n2281), .B2(
        \pc_lut[15][30] ), .ZN(n2901) );
  OAI221_X1 U4483 ( .B1(n2209), .B2(n2282), .C1(n2175), .C2(n2283), .A(n2902), 
        .ZN(n2897) );
  AOI22_X1 U4484 ( .A1(n2285), .A2(\pc_lut[2][30] ), .B1(n2286), .B2(
        \pc_lut[3][30] ), .ZN(n2902) );
  OAI221_X1 U4487 ( .B1(n2077), .B2(n2287), .C1(n2043), .C2(n2288), .A(n2903), 
        .ZN(n2896) );
  AOI22_X1 U4488 ( .A1(n2290), .A2(\pc_lut[6][30] ), .B1(n2291), .B2(
        \pc_lut[7][30] ), .ZN(n2903) );
  NAND2_X1 U4491 ( .A1(n2904), .A2(n2905), .ZN(N188) );
  NOR4_X1 U4492 ( .A1(n2906), .A2(n2907), .A3(n2908), .A4(n2909), .ZN(n2905)
         );
  OAI221_X1 U4493 ( .B1(n1443), .B2(n2248), .C1(n1409), .C2(n2249), .A(n2910), 
        .ZN(n2909) );
  AOI22_X1 U4494 ( .A1(n2251), .A2(\pc_lut[26][31] ), .B1(n2252), .B2(
        \pc_lut[27][31] ), .ZN(n2910) );
  OAI221_X1 U4497 ( .B1(n1308), .B2(n2253), .C1(n1274), .C2(n2254), .A(n2911), 
        .ZN(n2908) );
  AOI22_X1 U4498 ( .A1(n2256), .A2(\pc_lut[30][31] ), .B1(n2257), .B2(
        \pc_lut[31][31] ), .ZN(n2911) );
  OAI221_X1 U4501 ( .B1(n1707), .B2(n2258), .C1(n1673), .C2(n2259), .A(n2912), 
        .ZN(n2907) );
  AOI22_X1 U4502 ( .A1(n2261), .A2(\pc_lut[18][31] ), .B1(n2262), .B2(
        \pc_lut[19][31] ), .ZN(n2912) );
  OAI221_X1 U4505 ( .B1(n1512), .B2(n2263), .C1(n1477), .C2(n2264), .A(n2913), 
        .ZN(n2906) );
  AOI22_X1 U4506 ( .A1(n2266), .A2(\pc_lut[20][31] ), .B1(n2267), .B2(
        \pc_lut[21][31] ), .ZN(n2913) );
  NOR4_X1 U4509 ( .A1(n2914), .A2(n2915), .A3(n2916), .A4(n2917), .ZN(n2904)
         );
  OAI221_X1 U4510 ( .B1(n1977), .B2(n2272), .C1(n1943), .C2(n2273), .A(n2918), 
        .ZN(n2917) );
  AOI22_X1 U4511 ( .A1(n2275), .A2(\pc_lut[10][31] ), .B1(n2276), .B2(
        \pc_lut[11][31] ), .ZN(n2918) );
  OAI221_X1 U4514 ( .B1(n1842), .B2(n2277), .C1(n1808), .C2(n2278), .A(n2919), 
        .ZN(n2916) );
  AOI22_X1 U4515 ( .A1(n2280), .A2(\pc_lut[14][31] ), .B1(n2281), .B2(
        \pc_lut[15][31] ), .ZN(n2919) );
  OAI221_X1 U4518 ( .B1(n2241), .B2(n2282), .C1(n2207), .C2(n2283), .A(n2920), 
        .ZN(n2915) );
  AOI22_X1 U4519 ( .A1(n2285), .A2(\pc_lut[2][31] ), .B1(n2286), .B2(
        \pc_lut[3][31] ), .ZN(n2920) );
  OAI221_X1 U4522 ( .B1(n2109), .B2(n2287), .C1(n2075), .C2(n2288), .A(n2921), 
        .ZN(n2914) );
  AOI22_X1 U4523 ( .A1(n2290), .A2(\pc_lut[6][31] ), .B1(n2291), .B2(
        \pc_lut[7][31] ), .ZN(n2921) );
  NAND2_X1 U4526 ( .A1(n2922), .A2(n2923), .ZN(N127) );
  NOR4_X1 U4527 ( .A1(n2924), .A2(n2925), .A3(n2926), .A4(n2927), .ZN(n2923)
         );
  OAI221_X1 U4528 ( .B1(n299), .B2(n2248), .C1(n265), .C2(n2249), .A(n2928), 
        .ZN(n2927) );
  AOI22_X1 U4529 ( .A1(n2251), .A2(\pc_target[26][0] ), .B1(n2252), .B2(
        \pc_target[27][0] ), .ZN(n2928) );
  OAI221_X1 U4532 ( .B1(n159), .B2(n2253), .C1(n108), .C2(n2254), .A(n2929), 
        .ZN(n2926) );
  AOI22_X1 U4533 ( .A1(n2256), .A2(\pc_target[30][0] ), .B1(n2257), .B2(
        \pc_target[31][0] ), .ZN(n2929) );
  OAI221_X1 U4536 ( .B1(n575), .B2(n2258), .C1(n541), .C2(n2259), .A(n2930), 
        .ZN(n2925) );
  AOI22_X1 U4537 ( .A1(n2261), .A2(\pc_target[18][0] ), .B1(n2262), .B2(
        \pc_target[19][0] ), .ZN(n2930) );
  OAI221_X1 U4540 ( .B1(n369), .B2(n2263), .C1(n334), .C2(n2264), .A(n2931), 
        .ZN(n2924) );
  AOI22_X1 U4541 ( .A1(n2266), .A2(\pc_target[20][0] ), .B1(n2267), .B2(
        \pc_target[21][0] ), .ZN(n2931) );
  NOR4_X1 U4544 ( .A1(n2932), .A2(n2933), .A3(n2934), .A4(n2935), .ZN(n2922)
         );
  OAI221_X1 U4545 ( .B1(n852), .B2(n2272), .C1(n818), .C2(n2273), .A(n2936), 
        .ZN(n2935) );
  AOI22_X1 U4546 ( .A1(n2275), .A2(\pc_target[10][0] ), .B1(n2276), .B2(
        \pc_target[11][0] ), .ZN(n2936) );
  OAI221_X1 U4549 ( .B1(n714), .B2(n2277), .C1(n680), .C2(n2278), .A(n2937), 
        .ZN(n2934) );
  AOI22_X1 U4550 ( .A1(n2280), .A2(\pc_target[14][0] ), .B1(n2281), .B2(
        \pc_target[15][0] ), .ZN(n2937) );
  OAI221_X1 U4553 ( .B1(n1126), .B2(n2282), .C1(n1092), .C2(n2283), .A(n2938), 
        .ZN(n2933) );
  AOI22_X1 U4554 ( .A1(n2285), .A2(\pc_target[2][0] ), .B1(n2286), .B2(
        \pc_target[3][0] ), .ZN(n2938) );
  OAI221_X1 U4557 ( .B1(n989), .B2(n2287), .C1(n955), .C2(n2288), .A(n2939), 
        .ZN(n2932) );
  AOI22_X1 U4558 ( .A1(n2290), .A2(\pc_target[6][0] ), .B1(n2291), .B2(
        \pc_target[7][0] ), .ZN(n2939) );
  NAND2_X1 U4561 ( .A1(n2940), .A2(n2941), .ZN(N126) );
  NOR4_X1 U4562 ( .A1(n2942), .A2(n2943), .A3(n2944), .A4(n2945), .ZN(n2941)
         );
  OAI221_X1 U4563 ( .B1(n300), .B2(n2248), .C1(n266), .C2(n2249), .A(n2946), 
        .ZN(n2945) );
  AOI22_X1 U4564 ( .A1(n2251), .A2(\pc_target[26][1] ), .B1(n2252), .B2(
        \pc_target[27][1] ), .ZN(n2946) );
  OAI221_X1 U4567 ( .B1(n160), .B2(n2253), .C1(n110), .C2(n2254), .A(n2947), 
        .ZN(n2944) );
  AOI22_X1 U4568 ( .A1(n2256), .A2(\pc_target[30][1] ), .B1(n2257), .B2(
        \pc_target[31][1] ), .ZN(n2947) );
  OAI221_X1 U4571 ( .B1(n576), .B2(n2258), .C1(n542), .C2(n2259), .A(n2948), 
        .ZN(n2943) );
  AOI22_X1 U4572 ( .A1(n2261), .A2(\pc_target[18][1] ), .B1(n2262), .B2(
        \pc_target[19][1] ), .ZN(n2948) );
  OAI221_X1 U4575 ( .B1(n370), .B2(n2263), .C1(n335), .C2(n2264), .A(n2949), 
        .ZN(n2942) );
  AOI22_X1 U4576 ( .A1(n2266), .A2(\pc_target[20][1] ), .B1(n2267), .B2(
        \pc_target[21][1] ), .ZN(n2949) );
  NOR4_X1 U4579 ( .A1(n2950), .A2(n2951), .A3(n2952), .A4(n2953), .ZN(n2940)
         );
  OAI221_X1 U4580 ( .B1(n853), .B2(n2272), .C1(n819), .C2(n2273), .A(n2954), 
        .ZN(n2953) );
  AOI22_X1 U4581 ( .A1(n2275), .A2(\pc_target[10][1] ), .B1(n2276), .B2(
        \pc_target[11][1] ), .ZN(n2954) );
  OAI221_X1 U4584 ( .B1(n715), .B2(n2277), .C1(n681), .C2(n2278), .A(n2955), 
        .ZN(n2952) );
  AOI22_X1 U4585 ( .A1(n2280), .A2(\pc_target[14][1] ), .B1(n2281), .B2(
        \pc_target[15][1] ), .ZN(n2955) );
  OAI221_X1 U4588 ( .B1(n1127), .B2(n2282), .C1(n1093), .C2(n2283), .A(n2956), 
        .ZN(n2951) );
  AOI22_X1 U4589 ( .A1(n2285), .A2(\pc_target[2][1] ), .B1(n2286), .B2(
        \pc_target[3][1] ), .ZN(n2956) );
  OAI221_X1 U4592 ( .B1(n990), .B2(n2287), .C1(n956), .C2(n2288), .A(n2957), 
        .ZN(n2950) );
  AOI22_X1 U4593 ( .A1(n2290), .A2(\pc_target[6][1] ), .B1(n2291), .B2(
        \pc_target[7][1] ), .ZN(n2957) );
  NAND2_X1 U4596 ( .A1(n2958), .A2(n2959), .ZN(N125) );
  NOR4_X1 U4597 ( .A1(n2960), .A2(n2961), .A3(n2962), .A4(n2963), .ZN(n2959)
         );
  OAI221_X1 U4598 ( .B1(n298), .B2(n2248), .C1(n264), .C2(n2249), .A(n2964), 
        .ZN(n2963) );
  AOI22_X1 U4599 ( .A1(n2251), .A2(\pc_target[26][2] ), .B1(n2252), .B2(
        \pc_target[27][2] ), .ZN(n2964) );
  OAI221_X1 U4602 ( .B1(n158), .B2(n2253), .C1(n106), .C2(n2254), .A(n2965), 
        .ZN(n2962) );
  AOI22_X1 U4603 ( .A1(n2256), .A2(\pc_target[30][2] ), .B1(n2257), .B2(
        \pc_target[31][2] ), .ZN(n2965) );
  OAI221_X1 U4606 ( .B1(n574), .B2(n2258), .C1(n540), .C2(n2259), .A(n2966), 
        .ZN(n2961) );
  AOI22_X1 U4607 ( .A1(n2261), .A2(\pc_target[18][2] ), .B1(n2262), .B2(
        \pc_target[19][2] ), .ZN(n2966) );
  OAI221_X1 U4610 ( .B1(n368), .B2(n2263), .C1(n333), .C2(n2264), .A(n2967), 
        .ZN(n2960) );
  AOI22_X1 U4611 ( .A1(n2266), .A2(\pc_target[20][2] ), .B1(n2267), .B2(
        \pc_target[21][2] ), .ZN(n2967) );
  NOR4_X1 U4614 ( .A1(n2968), .A2(n2969), .A3(n2970), .A4(n2971), .ZN(n2958)
         );
  OAI221_X1 U4615 ( .B1(n851), .B2(n2272), .C1(n817), .C2(n2273), .A(n2972), 
        .ZN(n2971) );
  AOI22_X1 U4616 ( .A1(n2275), .A2(\pc_target[10][2] ), .B1(n2276), .B2(
        \pc_target[11][2] ), .ZN(n2972) );
  OAI221_X1 U4619 ( .B1(n713), .B2(n2277), .C1(n679), .C2(n2278), .A(n2973), 
        .ZN(n2970) );
  AOI22_X1 U4620 ( .A1(n2280), .A2(\pc_target[14][2] ), .B1(n2281), .B2(
        \pc_target[15][2] ), .ZN(n2973) );
  OAI221_X1 U4623 ( .B1(n1125), .B2(n2282), .C1(n1091), .C2(n2283), .A(n2974), 
        .ZN(n2969) );
  AOI22_X1 U4624 ( .A1(n2285), .A2(\pc_target[2][2] ), .B1(n2286), .B2(
        \pc_target[3][2] ), .ZN(n2974) );
  OAI221_X1 U4627 ( .B1(n988), .B2(n2287), .C1(n954), .C2(n2288), .A(n2975), 
        .ZN(n2968) );
  AOI22_X1 U4628 ( .A1(n2290), .A2(\pc_target[6][2] ), .B1(n2291), .B2(
        \pc_target[7][2] ), .ZN(n2975) );
  NAND2_X1 U4631 ( .A1(n2976), .A2(n2977), .ZN(N124) );
  NOR4_X1 U4632 ( .A1(n2978), .A2(n2979), .A3(n2980), .A4(n2981), .ZN(n2977)
         );
  OAI221_X1 U4633 ( .B1(n301), .B2(n2248), .C1(n267), .C2(n2249), .A(n2982), 
        .ZN(n2981) );
  AOI22_X1 U4634 ( .A1(n2251), .A2(\pc_target[26][3] ), .B1(n2252), .B2(
        \pc_target[27][3] ), .ZN(n2982) );
  OAI221_X1 U4637 ( .B1(n161), .B2(n2253), .C1(n112), .C2(n2254), .A(n2983), 
        .ZN(n2980) );
  AOI22_X1 U4638 ( .A1(n2256), .A2(\pc_target[30][3] ), .B1(n2257), .B2(
        \pc_target[31][3] ), .ZN(n2983) );
  OAI221_X1 U4641 ( .B1(n577), .B2(n2258), .C1(n543), .C2(n2259), .A(n2984), 
        .ZN(n2979) );
  AOI22_X1 U4642 ( .A1(n2261), .A2(\pc_target[18][3] ), .B1(n2262), .B2(
        \pc_target[19][3] ), .ZN(n2984) );
  OAI221_X1 U4645 ( .B1(n371), .B2(n2263), .C1(n336), .C2(n2264), .A(n2985), 
        .ZN(n2978) );
  AOI22_X1 U4646 ( .A1(n2266), .A2(\pc_target[20][3] ), .B1(n2267), .B2(
        \pc_target[21][3] ), .ZN(n2985) );
  NOR4_X1 U4649 ( .A1(n2986), .A2(n2987), .A3(n2988), .A4(n2989), .ZN(n2976)
         );
  OAI221_X1 U4650 ( .B1(n854), .B2(n2272), .C1(n820), .C2(n2273), .A(n2990), 
        .ZN(n2989) );
  AOI22_X1 U4651 ( .A1(n2275), .A2(\pc_target[10][3] ), .B1(n2276), .B2(
        \pc_target[11][3] ), .ZN(n2990) );
  OAI221_X1 U4654 ( .B1(n716), .B2(n2277), .C1(n682), .C2(n2278), .A(n2991), 
        .ZN(n2988) );
  AOI22_X1 U4655 ( .A1(n2280), .A2(\pc_target[14][3] ), .B1(n2281), .B2(
        \pc_target[15][3] ), .ZN(n2991) );
  OAI221_X1 U4658 ( .B1(n1128), .B2(n2282), .C1(n1094), .C2(n2283), .A(n2992), 
        .ZN(n2987) );
  AOI22_X1 U4659 ( .A1(n2285), .A2(\pc_target[2][3] ), .B1(n2286), .B2(
        \pc_target[3][3] ), .ZN(n2992) );
  OAI221_X1 U4662 ( .B1(n991), .B2(n2287), .C1(n957), .C2(n2288), .A(n2993), 
        .ZN(n2986) );
  AOI22_X1 U4663 ( .A1(n2290), .A2(\pc_target[6][3] ), .B1(n2291), .B2(
        \pc_target[7][3] ), .ZN(n2993) );
  NAND2_X1 U4666 ( .A1(n2994), .A2(n2995), .ZN(N123) );
  NOR4_X1 U4667 ( .A1(n2996), .A2(n2997), .A3(n2998), .A4(n2999), .ZN(n2995)
         );
  OAI221_X1 U4668 ( .B1(n297), .B2(n2248), .C1(n263), .C2(n2249), .A(n3000), 
        .ZN(n2999) );
  AOI22_X1 U4669 ( .A1(n2251), .A2(\pc_target[26][4] ), .B1(n2252), .B2(
        \pc_target[27][4] ), .ZN(n3000) );
  OAI221_X1 U4672 ( .B1(n157), .B2(n2253), .C1(n104), .C2(n2254), .A(n3001), 
        .ZN(n2998) );
  AOI22_X1 U4673 ( .A1(n2256), .A2(\pc_target[30][4] ), .B1(n2257), .B2(
        \pc_target[31][4] ), .ZN(n3001) );
  OAI221_X1 U4676 ( .B1(n573), .B2(n2258), .C1(n539), .C2(n2259), .A(n3002), 
        .ZN(n2997) );
  AOI22_X1 U4677 ( .A1(n2261), .A2(\pc_target[18][4] ), .B1(n2262), .B2(
        \pc_target[19][4] ), .ZN(n3002) );
  OAI221_X1 U4680 ( .B1(n367), .B2(n2263), .C1(n332), .C2(n2264), .A(n3003), 
        .ZN(n2996) );
  AOI22_X1 U4681 ( .A1(n2266), .A2(\pc_target[20][4] ), .B1(n2267), .B2(
        \pc_target[21][4] ), .ZN(n3003) );
  NOR4_X1 U4684 ( .A1(n3004), .A2(n3005), .A3(n3006), .A4(n3007), .ZN(n2994)
         );
  OAI221_X1 U4685 ( .B1(n850), .B2(n2272), .C1(n816), .C2(n2273), .A(n3008), 
        .ZN(n3007) );
  AOI22_X1 U4686 ( .A1(n2275), .A2(\pc_target[10][4] ), .B1(n2276), .B2(
        \pc_target[11][4] ), .ZN(n3008) );
  OAI221_X1 U4689 ( .B1(n712), .B2(n2277), .C1(n678), .C2(n2278), .A(n3009), 
        .ZN(n3006) );
  AOI22_X1 U4690 ( .A1(n2280), .A2(\pc_target[14][4] ), .B1(n2281), .B2(
        \pc_target[15][4] ), .ZN(n3009) );
  OAI221_X1 U4693 ( .B1(n1124), .B2(n2282), .C1(n1090), .C2(n2283), .A(n3010), 
        .ZN(n3005) );
  AOI22_X1 U4694 ( .A1(n2285), .A2(\pc_target[2][4] ), .B1(n2286), .B2(
        \pc_target[3][4] ), .ZN(n3010) );
  OAI221_X1 U4697 ( .B1(n987), .B2(n2287), .C1(n953), .C2(n2288), .A(n3011), 
        .ZN(n3004) );
  AOI22_X1 U4698 ( .A1(n2290), .A2(\pc_target[6][4] ), .B1(n2291), .B2(
        \pc_target[7][4] ), .ZN(n3011) );
  NAND2_X1 U4701 ( .A1(n3012), .A2(n3013), .ZN(N122) );
  NOR4_X1 U4702 ( .A1(n3014), .A2(n3015), .A3(n3016), .A4(n3017), .ZN(n3013)
         );
  OAI221_X1 U4703 ( .B1(n302), .B2(n2248), .C1(n268), .C2(n2249), .A(n3018), 
        .ZN(n3017) );
  AOI22_X1 U4704 ( .A1(n2251), .A2(\pc_target[26][5] ), .B1(n2252), .B2(
        \pc_target[27][5] ), .ZN(n3018) );
  OAI221_X1 U4707 ( .B1(n162), .B2(n2253), .C1(n114), .C2(n2254), .A(n3019), 
        .ZN(n3016) );
  AOI22_X1 U4708 ( .A1(n2256), .A2(\pc_target[30][5] ), .B1(n2257), .B2(
        \pc_target[31][5] ), .ZN(n3019) );
  OAI221_X1 U4711 ( .B1(n578), .B2(n2258), .C1(n544), .C2(n2259), .A(n3020), 
        .ZN(n3015) );
  AOI22_X1 U4712 ( .A1(n2261), .A2(\pc_target[18][5] ), .B1(n2262), .B2(
        \pc_target[19][5] ), .ZN(n3020) );
  OAI221_X1 U4715 ( .B1(n372), .B2(n2263), .C1(n337), .C2(n2264), .A(n3021), 
        .ZN(n3014) );
  AOI22_X1 U4716 ( .A1(n2266), .A2(\pc_target[20][5] ), .B1(n2267), .B2(
        \pc_target[21][5] ), .ZN(n3021) );
  NOR4_X1 U4719 ( .A1(n3022), .A2(n3023), .A3(n3024), .A4(n3025), .ZN(n3012)
         );
  OAI221_X1 U4720 ( .B1(n855), .B2(n2272), .C1(n821), .C2(n2273), .A(n3026), 
        .ZN(n3025) );
  AOI22_X1 U4721 ( .A1(n2275), .A2(\pc_target[10][5] ), .B1(n2276), .B2(
        \pc_target[11][5] ), .ZN(n3026) );
  OAI221_X1 U4724 ( .B1(n717), .B2(n2277), .C1(n683), .C2(n2278), .A(n3027), 
        .ZN(n3024) );
  AOI22_X1 U4725 ( .A1(n2280), .A2(\pc_target[14][5] ), .B1(n2281), .B2(
        \pc_target[15][5] ), .ZN(n3027) );
  OAI221_X1 U4728 ( .B1(n1129), .B2(n2282), .C1(n1095), .C2(n2283), .A(n3028), 
        .ZN(n3023) );
  AOI22_X1 U4729 ( .A1(n2285), .A2(\pc_target[2][5] ), .B1(n2286), .B2(
        \pc_target[3][5] ), .ZN(n3028) );
  OAI221_X1 U4732 ( .B1(n992), .B2(n2287), .C1(n958), .C2(n2288), .A(n3029), 
        .ZN(n3022) );
  AOI22_X1 U4733 ( .A1(n2290), .A2(\pc_target[6][5] ), .B1(n2291), .B2(
        \pc_target[7][5] ), .ZN(n3029) );
  NAND2_X1 U4736 ( .A1(n3030), .A2(n3031), .ZN(N121) );
  NOR4_X1 U4737 ( .A1(n3032), .A2(n3033), .A3(n3034), .A4(n3035), .ZN(n3031)
         );
  OAI221_X1 U4738 ( .B1(n296), .B2(n2248), .C1(n262), .C2(n2249), .A(n3036), 
        .ZN(n3035) );
  AOI22_X1 U4739 ( .A1(n2251), .A2(\pc_target[26][6] ), .B1(n2252), .B2(
        \pc_target[27][6] ), .ZN(n3036) );
  OAI221_X1 U4742 ( .B1(n156), .B2(n2253), .C1(n102), .C2(n2254), .A(n3037), 
        .ZN(n3034) );
  AOI22_X1 U4743 ( .A1(n2256), .A2(\pc_target[30][6] ), .B1(n2257), .B2(
        \pc_target[31][6] ), .ZN(n3037) );
  OAI221_X1 U4746 ( .B1(n572), .B2(n2258), .C1(n538), .C2(n2259), .A(n3038), 
        .ZN(n3033) );
  AOI22_X1 U4747 ( .A1(n2261), .A2(\pc_target[18][6] ), .B1(n2262), .B2(
        \pc_target[19][6] ), .ZN(n3038) );
  OAI221_X1 U4750 ( .B1(n366), .B2(n2263), .C1(n331), .C2(n2264), .A(n3039), 
        .ZN(n3032) );
  AOI22_X1 U4751 ( .A1(n2266), .A2(\pc_target[20][6] ), .B1(n2267), .B2(
        \pc_target[21][6] ), .ZN(n3039) );
  NOR4_X1 U4754 ( .A1(n3040), .A2(n3041), .A3(n3042), .A4(n3043), .ZN(n3030)
         );
  OAI221_X1 U4755 ( .B1(n849), .B2(n2272), .C1(n815), .C2(n2273), .A(n3044), 
        .ZN(n3043) );
  AOI22_X1 U4756 ( .A1(n2275), .A2(\pc_target[10][6] ), .B1(n2276), .B2(
        \pc_target[11][6] ), .ZN(n3044) );
  OAI221_X1 U4759 ( .B1(n711), .B2(n2277), .C1(n677), .C2(n2278), .A(n3045), 
        .ZN(n3042) );
  AOI22_X1 U4760 ( .A1(n2280), .A2(\pc_target[14][6] ), .B1(n2281), .B2(
        \pc_target[15][6] ), .ZN(n3045) );
  OAI221_X1 U4763 ( .B1(n1123), .B2(n2282), .C1(n1089), .C2(n2283), .A(n3046), 
        .ZN(n3041) );
  AOI22_X1 U4764 ( .A1(n2285), .A2(\pc_target[2][6] ), .B1(n2286), .B2(
        \pc_target[3][6] ), .ZN(n3046) );
  OAI221_X1 U4767 ( .B1(n986), .B2(n2287), .C1(n952), .C2(n2288), .A(n3047), 
        .ZN(n3040) );
  AOI22_X1 U4768 ( .A1(n2290), .A2(\pc_target[6][6] ), .B1(n2291), .B2(
        \pc_target[7][6] ), .ZN(n3047) );
  NAND2_X1 U4771 ( .A1(n3048), .A2(n3049), .ZN(N120) );
  NOR4_X1 U4772 ( .A1(n3050), .A2(n3051), .A3(n3052), .A4(n3053), .ZN(n3049)
         );
  OAI221_X1 U4773 ( .B1(n303), .B2(n2248), .C1(n269), .C2(n2249), .A(n3054), 
        .ZN(n3053) );
  AOI22_X1 U4774 ( .A1(n2251), .A2(\pc_target[26][7] ), .B1(n2252), .B2(
        \pc_target[27][7] ), .ZN(n3054) );
  OAI221_X1 U4777 ( .B1(n163), .B2(n2253), .C1(n116), .C2(n2254), .A(n3055), 
        .ZN(n3052) );
  AOI22_X1 U4778 ( .A1(n2256), .A2(\pc_target[30][7] ), .B1(n2257), .B2(
        \pc_target[31][7] ), .ZN(n3055) );
  OAI221_X1 U4781 ( .B1(n579), .B2(n2258), .C1(n545), .C2(n2259), .A(n3056), 
        .ZN(n3051) );
  AOI22_X1 U4782 ( .A1(n2261), .A2(\pc_target[18][7] ), .B1(n2262), .B2(
        \pc_target[19][7] ), .ZN(n3056) );
  OAI221_X1 U4785 ( .B1(n373), .B2(n2263), .C1(n338), .C2(n2264), .A(n3057), 
        .ZN(n3050) );
  AOI22_X1 U4786 ( .A1(n2266), .A2(\pc_target[20][7] ), .B1(n2267), .B2(
        \pc_target[21][7] ), .ZN(n3057) );
  NOR4_X1 U4789 ( .A1(n3058), .A2(n3059), .A3(n3060), .A4(n3061), .ZN(n3048)
         );
  OAI221_X1 U4790 ( .B1(n856), .B2(n2272), .C1(n822), .C2(n2273), .A(n3062), 
        .ZN(n3061) );
  AOI22_X1 U4791 ( .A1(n2275), .A2(\pc_target[10][7] ), .B1(n2276), .B2(
        \pc_target[11][7] ), .ZN(n3062) );
  OAI221_X1 U4794 ( .B1(n718), .B2(n2277), .C1(n684), .C2(n2278), .A(n3063), 
        .ZN(n3060) );
  AOI22_X1 U4795 ( .A1(n2280), .A2(\pc_target[14][7] ), .B1(n2281), .B2(
        \pc_target[15][7] ), .ZN(n3063) );
  OAI221_X1 U4798 ( .B1(n1130), .B2(n2282), .C1(n1096), .C2(n2283), .A(n3064), 
        .ZN(n3059) );
  AOI22_X1 U4799 ( .A1(n2285), .A2(\pc_target[2][7] ), .B1(n2286), .B2(
        \pc_target[3][7] ), .ZN(n3064) );
  OAI221_X1 U4802 ( .B1(n993), .B2(n2287), .C1(n959), .C2(n2288), .A(n3065), 
        .ZN(n3058) );
  AOI22_X1 U4803 ( .A1(n2290), .A2(\pc_target[6][7] ), .B1(n2291), .B2(
        \pc_target[7][7] ), .ZN(n3065) );
  NAND2_X1 U4806 ( .A1(n3066), .A2(n3067), .ZN(N119) );
  NOR4_X1 U4807 ( .A1(n3068), .A2(n3069), .A3(n3070), .A4(n3071), .ZN(n3067)
         );
  OAI221_X1 U4808 ( .B1(n295), .B2(n2248), .C1(n261), .C2(n2249), .A(n3072), 
        .ZN(n3071) );
  AOI22_X1 U4809 ( .A1(n2251), .A2(\pc_target[26][8] ), .B1(n2252), .B2(
        \pc_target[27][8] ), .ZN(n3072) );
  OAI221_X1 U4812 ( .B1(n155), .B2(n2253), .C1(n100), .C2(n2254), .A(n3073), 
        .ZN(n3070) );
  AOI22_X1 U4813 ( .A1(n2256), .A2(\pc_target[30][8] ), .B1(n2257), .B2(
        \pc_target[31][8] ), .ZN(n3073) );
  OAI221_X1 U4816 ( .B1(n571), .B2(n2258), .C1(n537), .C2(n2259), .A(n3074), 
        .ZN(n3069) );
  AOI22_X1 U4817 ( .A1(n2261), .A2(\pc_target[18][8] ), .B1(n2262), .B2(
        \pc_target[19][8] ), .ZN(n3074) );
  OAI221_X1 U4820 ( .B1(n365), .B2(n2263), .C1(n330), .C2(n2264), .A(n3075), 
        .ZN(n3068) );
  AOI22_X1 U4821 ( .A1(n2266), .A2(\pc_target[20][8] ), .B1(n2267), .B2(
        \pc_target[21][8] ), .ZN(n3075) );
  NOR4_X1 U4824 ( .A1(n3076), .A2(n3077), .A3(n3078), .A4(n3079), .ZN(n3066)
         );
  OAI221_X1 U4825 ( .B1(n848), .B2(n2272), .C1(n814), .C2(n2273), .A(n3080), 
        .ZN(n3079) );
  AOI22_X1 U4826 ( .A1(n2275), .A2(\pc_target[10][8] ), .B1(n2276), .B2(
        \pc_target[11][8] ), .ZN(n3080) );
  OAI221_X1 U4829 ( .B1(n710), .B2(n2277), .C1(n676), .C2(n2278), .A(n3081), 
        .ZN(n3078) );
  AOI22_X1 U4830 ( .A1(n2280), .A2(\pc_target[14][8] ), .B1(n2281), .B2(
        \pc_target[15][8] ), .ZN(n3081) );
  OAI221_X1 U4833 ( .B1(n1122), .B2(n2282), .C1(n1088), .C2(n2283), .A(n3082), 
        .ZN(n3077) );
  AOI22_X1 U4834 ( .A1(n2285), .A2(\pc_target[2][8] ), .B1(n2286), .B2(
        \pc_target[3][8] ), .ZN(n3082) );
  OAI221_X1 U4837 ( .B1(n985), .B2(n2287), .C1(n951), .C2(n2288), .A(n3083), 
        .ZN(n3076) );
  AOI22_X1 U4838 ( .A1(n2290), .A2(\pc_target[6][8] ), .B1(n2291), .B2(
        \pc_target[7][8] ), .ZN(n3083) );
  NAND2_X1 U4841 ( .A1(n3084), .A2(n3085), .ZN(N118) );
  NOR4_X1 U4842 ( .A1(n3086), .A2(n3087), .A3(n3088), .A4(n3089), .ZN(n3085)
         );
  OAI221_X1 U4843 ( .B1(n304), .B2(n2248), .C1(n270), .C2(n2249), .A(n3090), 
        .ZN(n3089) );
  AOI22_X1 U4844 ( .A1(n2251), .A2(\pc_target[26][9] ), .B1(n2252), .B2(
        \pc_target[27][9] ), .ZN(n3090) );
  OAI221_X1 U4847 ( .B1(n164), .B2(n2253), .C1(n118), .C2(n2254), .A(n3091), 
        .ZN(n3088) );
  AOI22_X1 U4848 ( .A1(n2256), .A2(\pc_target[30][9] ), .B1(n2257), .B2(
        \pc_target[31][9] ), .ZN(n3091) );
  OAI221_X1 U4851 ( .B1(n580), .B2(n2258), .C1(n546), .C2(n2259), .A(n3092), 
        .ZN(n3087) );
  AOI22_X1 U4852 ( .A1(n2261), .A2(\pc_target[18][9] ), .B1(n2262), .B2(
        \pc_target[19][9] ), .ZN(n3092) );
  OAI221_X1 U4855 ( .B1(n374), .B2(n2263), .C1(n339), .C2(n2264), .A(n3093), 
        .ZN(n3086) );
  AOI22_X1 U4856 ( .A1(n2266), .A2(\pc_target[20][9] ), .B1(n2267), .B2(
        \pc_target[21][9] ), .ZN(n3093) );
  NOR4_X1 U4859 ( .A1(n3094), .A2(n3095), .A3(n3096), .A4(n3097), .ZN(n3084)
         );
  OAI221_X1 U4860 ( .B1(n857), .B2(n2272), .C1(n823), .C2(n2273), .A(n3098), 
        .ZN(n3097) );
  AOI22_X1 U4861 ( .A1(n2275), .A2(\pc_target[10][9] ), .B1(n2276), .B2(
        \pc_target[11][9] ), .ZN(n3098) );
  OAI221_X1 U4864 ( .B1(n719), .B2(n2277), .C1(n685), .C2(n2278), .A(n3099), 
        .ZN(n3096) );
  AOI22_X1 U4865 ( .A1(n2280), .A2(\pc_target[14][9] ), .B1(n2281), .B2(
        \pc_target[15][9] ), .ZN(n3099) );
  OAI221_X1 U4868 ( .B1(n1131), .B2(n2282), .C1(n1097), .C2(n2283), .A(n3100), 
        .ZN(n3095) );
  AOI22_X1 U4869 ( .A1(n2285), .A2(\pc_target[2][9] ), .B1(n2286), .B2(
        \pc_target[3][9] ), .ZN(n3100) );
  OAI221_X1 U4872 ( .B1(n994), .B2(n2287), .C1(n960), .C2(n2288), .A(n3101), 
        .ZN(n3094) );
  AOI22_X1 U4873 ( .A1(n2290), .A2(\pc_target[6][9] ), .B1(n2291), .B2(
        \pc_target[7][9] ), .ZN(n3101) );
  NAND2_X1 U4876 ( .A1(n3102), .A2(n3103), .ZN(N117) );
  NOR4_X1 U4877 ( .A1(n3104), .A2(n3105), .A3(n3106), .A4(n3107), .ZN(n3103)
         );
  OAI221_X1 U4878 ( .B1(n294), .B2(n2248), .C1(n260), .C2(n2249), .A(n3108), 
        .ZN(n3107) );
  AOI22_X1 U4879 ( .A1(n2251), .A2(\pc_target[26][10] ), .B1(n2252), .B2(
        \pc_target[27][10] ), .ZN(n3108) );
  OAI221_X1 U4882 ( .B1(n154), .B2(n2253), .C1(n98), .C2(n2254), .A(n3109), 
        .ZN(n3106) );
  AOI22_X1 U4883 ( .A1(n2256), .A2(\pc_target[30][10] ), .B1(n2257), .B2(
        \pc_target[31][10] ), .ZN(n3109) );
  OAI221_X1 U4886 ( .B1(n570), .B2(n2258), .C1(n536), .C2(n2259), .A(n3110), 
        .ZN(n3105) );
  AOI22_X1 U4887 ( .A1(n2261), .A2(\pc_target[18][10] ), .B1(n2262), .B2(
        \pc_target[19][10] ), .ZN(n3110) );
  OAI221_X1 U4890 ( .B1(n364), .B2(n2263), .C1(n329), .C2(n2264), .A(n3111), 
        .ZN(n3104) );
  AOI22_X1 U4891 ( .A1(n2266), .A2(\pc_target[20][10] ), .B1(n2267), .B2(
        \pc_target[21][10] ), .ZN(n3111) );
  NOR4_X1 U4894 ( .A1(n3112), .A2(n3113), .A3(n3114), .A4(n3115), .ZN(n3102)
         );
  OAI221_X1 U4895 ( .B1(n847), .B2(n2272), .C1(n813), .C2(n2273), .A(n3116), 
        .ZN(n3115) );
  AOI22_X1 U4896 ( .A1(n2275), .A2(\pc_target[10][10] ), .B1(n2276), .B2(
        \pc_target[11][10] ), .ZN(n3116) );
  OAI221_X1 U4899 ( .B1(n709), .B2(n2277), .C1(n675), .C2(n2278), .A(n3117), 
        .ZN(n3114) );
  AOI22_X1 U4900 ( .A1(n2280), .A2(\pc_target[14][10] ), .B1(n2281), .B2(
        \pc_target[15][10] ), .ZN(n3117) );
  OAI221_X1 U4903 ( .B1(n1121), .B2(n2282), .C1(n1087), .C2(n2283), .A(n3118), 
        .ZN(n3113) );
  AOI22_X1 U4904 ( .A1(n2285), .A2(\pc_target[2][10] ), .B1(n2286), .B2(
        \pc_target[3][10] ), .ZN(n3118) );
  OAI221_X1 U4907 ( .B1(n984), .B2(n2287), .C1(n950), .C2(n2288), .A(n3119), 
        .ZN(n3112) );
  AOI22_X1 U4908 ( .A1(n2290), .A2(\pc_target[6][10] ), .B1(n2291), .B2(
        \pc_target[7][10] ), .ZN(n3119) );
  NAND2_X1 U4911 ( .A1(n3120), .A2(n3121), .ZN(N116) );
  NOR4_X1 U4912 ( .A1(n3122), .A2(n3123), .A3(n3124), .A4(n3125), .ZN(n3121)
         );
  OAI221_X1 U4913 ( .B1(n305), .B2(n2248), .C1(n271), .C2(n2249), .A(n3126), 
        .ZN(n3125) );
  AOI22_X1 U4914 ( .A1(n2251), .A2(\pc_target[26][11] ), .B1(n2252), .B2(
        \pc_target[27][11] ), .ZN(n3126) );
  OAI221_X1 U4917 ( .B1(n165), .B2(n2253), .C1(n120), .C2(n2254), .A(n3127), 
        .ZN(n3124) );
  AOI22_X1 U4918 ( .A1(n2256), .A2(\pc_target[30][11] ), .B1(n2257), .B2(
        \pc_target[31][11] ), .ZN(n3127) );
  OAI221_X1 U4921 ( .B1(n581), .B2(n2258), .C1(n547), .C2(n2259), .A(n3128), 
        .ZN(n3123) );
  AOI22_X1 U4922 ( .A1(n2261), .A2(\pc_target[18][11] ), .B1(n2262), .B2(
        \pc_target[19][11] ), .ZN(n3128) );
  OAI221_X1 U4925 ( .B1(n375), .B2(n2263), .C1(n340), .C2(n2264), .A(n3129), 
        .ZN(n3122) );
  AOI22_X1 U4926 ( .A1(n2266), .A2(\pc_target[20][11] ), .B1(n2267), .B2(
        \pc_target[21][11] ), .ZN(n3129) );
  NOR4_X1 U4929 ( .A1(n3130), .A2(n3131), .A3(n3132), .A4(n3133), .ZN(n3120)
         );
  OAI221_X1 U4930 ( .B1(n858), .B2(n2272), .C1(n824), .C2(n2273), .A(n3134), 
        .ZN(n3133) );
  AOI22_X1 U4931 ( .A1(n2275), .A2(\pc_target[10][11] ), .B1(n2276), .B2(
        \pc_target[11][11] ), .ZN(n3134) );
  OAI221_X1 U4934 ( .B1(n720), .B2(n2277), .C1(n686), .C2(n2278), .A(n3135), 
        .ZN(n3132) );
  AOI22_X1 U4935 ( .A1(n2280), .A2(\pc_target[14][11] ), .B1(n2281), .B2(
        \pc_target[15][11] ), .ZN(n3135) );
  OAI221_X1 U4938 ( .B1(n1132), .B2(n2282), .C1(n1098), .C2(n2283), .A(n3136), 
        .ZN(n3131) );
  AOI22_X1 U4939 ( .A1(n2285), .A2(\pc_target[2][11] ), .B1(n2286), .B2(
        \pc_target[3][11] ), .ZN(n3136) );
  OAI221_X1 U4942 ( .B1(n995), .B2(n2287), .C1(n961), .C2(n2288), .A(n3137), 
        .ZN(n3130) );
  AOI22_X1 U4943 ( .A1(n2290), .A2(\pc_target[6][11] ), .B1(n2291), .B2(
        \pc_target[7][11] ), .ZN(n3137) );
  NAND2_X1 U4946 ( .A1(n3138), .A2(n3139), .ZN(N115) );
  NOR4_X1 U4947 ( .A1(n3140), .A2(n3141), .A3(n3142), .A4(n3143), .ZN(n3139)
         );
  OAI221_X1 U4948 ( .B1(n293), .B2(n2248), .C1(n259), .C2(n2249), .A(n3144), 
        .ZN(n3143) );
  AOI22_X1 U4949 ( .A1(n2251), .A2(\pc_target[26][12] ), .B1(n2252), .B2(
        \pc_target[27][12] ), .ZN(n3144) );
  OAI221_X1 U4952 ( .B1(n153), .B2(n2253), .C1(n96), .C2(n2254), .A(n3145), 
        .ZN(n3142) );
  AOI22_X1 U4953 ( .A1(n2256), .A2(\pc_target[30][12] ), .B1(n2257), .B2(
        \pc_target[31][12] ), .ZN(n3145) );
  OAI221_X1 U4956 ( .B1(n569), .B2(n2258), .C1(n535), .C2(n2259), .A(n3146), 
        .ZN(n3141) );
  AOI22_X1 U4957 ( .A1(n2261), .A2(\pc_target[18][12] ), .B1(n2262), .B2(
        \pc_target[19][12] ), .ZN(n3146) );
  OAI221_X1 U4960 ( .B1(n363), .B2(n2263), .C1(n328), .C2(n2264), .A(n3147), 
        .ZN(n3140) );
  AOI22_X1 U4961 ( .A1(n2266), .A2(\pc_target[20][12] ), .B1(n2267), .B2(
        \pc_target[21][12] ), .ZN(n3147) );
  NOR4_X1 U4964 ( .A1(n3148), .A2(n3149), .A3(n3150), .A4(n3151), .ZN(n3138)
         );
  OAI221_X1 U4965 ( .B1(n846), .B2(n2272), .C1(n812), .C2(n2273), .A(n3152), 
        .ZN(n3151) );
  AOI22_X1 U4966 ( .A1(n2275), .A2(\pc_target[10][12] ), .B1(n2276), .B2(
        \pc_target[11][12] ), .ZN(n3152) );
  OAI221_X1 U4969 ( .B1(n708), .B2(n2277), .C1(n674), .C2(n2278), .A(n3153), 
        .ZN(n3150) );
  AOI22_X1 U4970 ( .A1(n2280), .A2(\pc_target[14][12] ), .B1(n2281), .B2(
        \pc_target[15][12] ), .ZN(n3153) );
  OAI221_X1 U4973 ( .B1(n1120), .B2(n2282), .C1(n1086), .C2(n2283), .A(n3154), 
        .ZN(n3149) );
  AOI22_X1 U4974 ( .A1(n2285), .A2(\pc_target[2][12] ), .B1(n2286), .B2(
        \pc_target[3][12] ), .ZN(n3154) );
  OAI221_X1 U4977 ( .B1(n983), .B2(n2287), .C1(n949), .C2(n2288), .A(n3155), 
        .ZN(n3148) );
  AOI22_X1 U4978 ( .A1(n2290), .A2(\pc_target[6][12] ), .B1(n2291), .B2(
        \pc_target[7][12] ), .ZN(n3155) );
  NAND2_X1 U4981 ( .A1(n3156), .A2(n3157), .ZN(N114) );
  NOR4_X1 U4982 ( .A1(n3158), .A2(n3159), .A3(n3160), .A4(n3161), .ZN(n3157)
         );
  OAI221_X1 U4983 ( .B1(n306), .B2(n2248), .C1(n272), .C2(n2249), .A(n3162), 
        .ZN(n3161) );
  AOI22_X1 U4984 ( .A1(n2251), .A2(\pc_target[26][13] ), .B1(n2252), .B2(
        \pc_target[27][13] ), .ZN(n3162) );
  OAI221_X1 U4987 ( .B1(n166), .B2(n2253), .C1(n122), .C2(n2254), .A(n3163), 
        .ZN(n3160) );
  AOI22_X1 U4988 ( .A1(n2256), .A2(\pc_target[30][13] ), .B1(n2257), .B2(
        \pc_target[31][13] ), .ZN(n3163) );
  OAI221_X1 U4991 ( .B1(n582), .B2(n2258), .C1(n548), .C2(n2259), .A(n3164), 
        .ZN(n3159) );
  AOI22_X1 U4992 ( .A1(n2261), .A2(\pc_target[18][13] ), .B1(n2262), .B2(
        \pc_target[19][13] ), .ZN(n3164) );
  OAI221_X1 U4995 ( .B1(n376), .B2(n2263), .C1(n341), .C2(n2264), .A(n3165), 
        .ZN(n3158) );
  AOI22_X1 U4996 ( .A1(n2266), .A2(\pc_target[20][13] ), .B1(n2267), .B2(
        \pc_target[21][13] ), .ZN(n3165) );
  NOR4_X1 U4999 ( .A1(n3166), .A2(n3167), .A3(n3168), .A4(n3169), .ZN(n3156)
         );
  OAI221_X1 U5000 ( .B1(n859), .B2(n2272), .C1(n825), .C2(n2273), .A(n3170), 
        .ZN(n3169) );
  AOI22_X1 U5001 ( .A1(n2275), .A2(\pc_target[10][13] ), .B1(n2276), .B2(
        \pc_target[11][13] ), .ZN(n3170) );
  OAI221_X1 U5004 ( .B1(n721), .B2(n2277), .C1(n687), .C2(n2278), .A(n3171), 
        .ZN(n3168) );
  AOI22_X1 U5005 ( .A1(n2280), .A2(\pc_target[14][13] ), .B1(n2281), .B2(
        \pc_target[15][13] ), .ZN(n3171) );
  OAI221_X1 U5008 ( .B1(n1133), .B2(n2282), .C1(n1099), .C2(n2283), .A(n3172), 
        .ZN(n3167) );
  AOI22_X1 U5009 ( .A1(n2285), .A2(\pc_target[2][13] ), .B1(n2286), .B2(
        \pc_target[3][13] ), .ZN(n3172) );
  OAI221_X1 U5012 ( .B1(n996), .B2(n2287), .C1(n962), .C2(n2288), .A(n3173), 
        .ZN(n3166) );
  AOI22_X1 U5013 ( .A1(n2290), .A2(\pc_target[6][13] ), .B1(n2291), .B2(
        \pc_target[7][13] ), .ZN(n3173) );
  NAND2_X1 U5016 ( .A1(n3174), .A2(n3175), .ZN(N113) );
  NOR4_X1 U5017 ( .A1(n3176), .A2(n3177), .A3(n3178), .A4(n3179), .ZN(n3175)
         );
  OAI221_X1 U5018 ( .B1(n292), .B2(n2248), .C1(n258), .C2(n2249), .A(n3180), 
        .ZN(n3179) );
  AOI22_X1 U5019 ( .A1(n2251), .A2(\pc_target[26][14] ), .B1(n2252), .B2(
        \pc_target[27][14] ), .ZN(n3180) );
  OAI221_X1 U5022 ( .B1(n152), .B2(n2253), .C1(n94), .C2(n2254), .A(n3181), 
        .ZN(n3178) );
  AOI22_X1 U5023 ( .A1(n2256), .A2(\pc_target[30][14] ), .B1(n2257), .B2(
        \pc_target[31][14] ), .ZN(n3181) );
  OAI221_X1 U5026 ( .B1(n568), .B2(n2258), .C1(n534), .C2(n2259), .A(n3182), 
        .ZN(n3177) );
  AOI22_X1 U5027 ( .A1(n2261), .A2(\pc_target[18][14] ), .B1(n2262), .B2(
        \pc_target[19][14] ), .ZN(n3182) );
  OAI221_X1 U5030 ( .B1(n362), .B2(n2263), .C1(n327), .C2(n2264), .A(n3183), 
        .ZN(n3176) );
  AOI22_X1 U5031 ( .A1(n2266), .A2(\pc_target[20][14] ), .B1(n2267), .B2(
        \pc_target[21][14] ), .ZN(n3183) );
  NOR4_X1 U5034 ( .A1(n3184), .A2(n3185), .A3(n3186), .A4(n3187), .ZN(n3174)
         );
  OAI221_X1 U5035 ( .B1(n845), .B2(n2272), .C1(n811), .C2(n2273), .A(n3188), 
        .ZN(n3187) );
  AOI22_X1 U5036 ( .A1(n2275), .A2(\pc_target[10][14] ), .B1(n2276), .B2(
        \pc_target[11][14] ), .ZN(n3188) );
  OAI221_X1 U5039 ( .B1(n707), .B2(n2277), .C1(n673), .C2(n2278), .A(n3189), 
        .ZN(n3186) );
  AOI22_X1 U5040 ( .A1(n2280), .A2(\pc_target[14][14] ), .B1(n2281), .B2(
        \pc_target[15][14] ), .ZN(n3189) );
  OAI221_X1 U5043 ( .B1(n1119), .B2(n2282), .C1(n1085), .C2(n2283), .A(n3190), 
        .ZN(n3185) );
  AOI22_X1 U5044 ( .A1(n2285), .A2(\pc_target[2][14] ), .B1(n2286), .B2(
        \pc_target[3][14] ), .ZN(n3190) );
  OAI221_X1 U5047 ( .B1(n982), .B2(n2287), .C1(n948), .C2(n2288), .A(n3191), 
        .ZN(n3184) );
  AOI22_X1 U5048 ( .A1(n2290), .A2(\pc_target[6][14] ), .B1(n2291), .B2(
        \pc_target[7][14] ), .ZN(n3191) );
  NAND2_X1 U5051 ( .A1(n3192), .A2(n3193), .ZN(N112) );
  NOR4_X1 U5052 ( .A1(n3194), .A2(n3195), .A3(n3196), .A4(n3197), .ZN(n3193)
         );
  OAI221_X1 U5053 ( .B1(n307), .B2(n2248), .C1(n273), .C2(n2249), .A(n3198), 
        .ZN(n3197) );
  AOI22_X1 U5054 ( .A1(n2251), .A2(\pc_target[26][15] ), .B1(n2252), .B2(
        \pc_target[27][15] ), .ZN(n3198) );
  OAI221_X1 U5057 ( .B1(n167), .B2(n2253), .C1(n124), .C2(n2254), .A(n3199), 
        .ZN(n3196) );
  AOI22_X1 U5058 ( .A1(n2256), .A2(\pc_target[30][15] ), .B1(n2257), .B2(
        \pc_target[31][15] ), .ZN(n3199) );
  OAI221_X1 U5061 ( .B1(n583), .B2(n2258), .C1(n549), .C2(n2259), .A(n3200), 
        .ZN(n3195) );
  AOI22_X1 U5062 ( .A1(n2261), .A2(\pc_target[18][15] ), .B1(n2262), .B2(
        \pc_target[19][15] ), .ZN(n3200) );
  OAI221_X1 U5065 ( .B1(n377), .B2(n2263), .C1(n342), .C2(n2264), .A(n3201), 
        .ZN(n3194) );
  AOI22_X1 U5066 ( .A1(n2266), .A2(\pc_target[20][15] ), .B1(n2267), .B2(
        \pc_target[21][15] ), .ZN(n3201) );
  NOR4_X1 U5069 ( .A1(n3202), .A2(n3203), .A3(n3204), .A4(n3205), .ZN(n3192)
         );
  OAI221_X1 U5070 ( .B1(n860), .B2(n2272), .C1(n826), .C2(n2273), .A(n3206), 
        .ZN(n3205) );
  AOI22_X1 U5071 ( .A1(n2275), .A2(\pc_target[10][15] ), .B1(n2276), .B2(
        \pc_target[11][15] ), .ZN(n3206) );
  OAI221_X1 U5074 ( .B1(n722), .B2(n2277), .C1(n688), .C2(n2278), .A(n3207), 
        .ZN(n3204) );
  AOI22_X1 U5075 ( .A1(n2280), .A2(\pc_target[14][15] ), .B1(n2281), .B2(
        \pc_target[15][15] ), .ZN(n3207) );
  OAI221_X1 U5078 ( .B1(n1134), .B2(n2282), .C1(n1100), .C2(n2283), .A(n3208), 
        .ZN(n3203) );
  AOI22_X1 U5079 ( .A1(n2285), .A2(\pc_target[2][15] ), .B1(n2286), .B2(
        \pc_target[3][15] ), .ZN(n3208) );
  OAI221_X1 U5082 ( .B1(n997), .B2(n2287), .C1(n963), .C2(n2288), .A(n3209), 
        .ZN(n3202) );
  AOI22_X1 U5083 ( .A1(n2290), .A2(\pc_target[6][15] ), .B1(n2291), .B2(
        \pc_target[7][15] ), .ZN(n3209) );
  NAND2_X1 U5086 ( .A1(n3210), .A2(n3211), .ZN(N111) );
  NOR4_X1 U5087 ( .A1(n3212), .A2(n3213), .A3(n3214), .A4(n3215), .ZN(n3211)
         );
  OAI221_X1 U5088 ( .B1(n291), .B2(n2248), .C1(n257), .C2(n2249), .A(n3216), 
        .ZN(n3215) );
  AOI22_X1 U5089 ( .A1(n2251), .A2(\pc_target[26][16] ), .B1(n2252), .B2(
        \pc_target[27][16] ), .ZN(n3216) );
  OAI221_X1 U5092 ( .B1(n151), .B2(n2253), .C1(n92), .C2(n2254), .A(n3217), 
        .ZN(n3214) );
  AOI22_X1 U5093 ( .A1(n2256), .A2(\pc_target[30][16] ), .B1(n2257), .B2(
        \pc_target[31][16] ), .ZN(n3217) );
  OAI221_X1 U5096 ( .B1(n567), .B2(n2258), .C1(n533), .C2(n2259), .A(n3218), 
        .ZN(n3213) );
  AOI22_X1 U5097 ( .A1(n2261), .A2(\pc_target[18][16] ), .B1(n2262), .B2(
        \pc_target[19][16] ), .ZN(n3218) );
  OAI221_X1 U5100 ( .B1(n361), .B2(n2263), .C1(n326), .C2(n2264), .A(n3219), 
        .ZN(n3212) );
  AOI22_X1 U5101 ( .A1(n2266), .A2(\pc_target[20][16] ), .B1(n2267), .B2(
        \pc_target[21][16] ), .ZN(n3219) );
  NOR4_X1 U5104 ( .A1(n3220), .A2(n3221), .A3(n3222), .A4(n3223), .ZN(n3210)
         );
  OAI221_X1 U5105 ( .B1(n844), .B2(n2272), .C1(n810), .C2(n2273), .A(n3224), 
        .ZN(n3223) );
  AOI22_X1 U5106 ( .A1(n2275), .A2(\pc_target[10][16] ), .B1(n2276), .B2(
        \pc_target[11][16] ), .ZN(n3224) );
  OAI221_X1 U5109 ( .B1(n706), .B2(n2277), .C1(n672), .C2(n2278), .A(n3225), 
        .ZN(n3222) );
  AOI22_X1 U5110 ( .A1(n2280), .A2(\pc_target[14][16] ), .B1(n2281), .B2(
        \pc_target[15][16] ), .ZN(n3225) );
  OAI221_X1 U5113 ( .B1(n1118), .B2(n2282), .C1(n1084), .C2(n2283), .A(n3226), 
        .ZN(n3221) );
  AOI22_X1 U5114 ( .A1(n2285), .A2(\pc_target[2][16] ), .B1(n2286), .B2(
        \pc_target[3][16] ), .ZN(n3226) );
  OAI221_X1 U5117 ( .B1(n981), .B2(n2287), .C1(n947), .C2(n2288), .A(n3227), 
        .ZN(n3220) );
  AOI22_X1 U5118 ( .A1(n2290), .A2(\pc_target[6][16] ), .B1(n2291), .B2(
        \pc_target[7][16] ), .ZN(n3227) );
  NAND2_X1 U5121 ( .A1(n3228), .A2(n3229), .ZN(N110) );
  NOR4_X1 U5122 ( .A1(n3230), .A2(n3231), .A3(n3232), .A4(n3233), .ZN(n3229)
         );
  OAI221_X1 U5123 ( .B1(n308), .B2(n2248), .C1(n274), .C2(n2249), .A(n3234), 
        .ZN(n3233) );
  AOI22_X1 U5124 ( .A1(n2251), .A2(\pc_target[26][17] ), .B1(n2252), .B2(
        \pc_target[27][17] ), .ZN(n3234) );
  OAI221_X1 U5127 ( .B1(n168), .B2(n2253), .C1(n126), .C2(n2254), .A(n3235), 
        .ZN(n3232) );
  AOI22_X1 U5128 ( .A1(n2256), .A2(\pc_target[30][17] ), .B1(n2257), .B2(
        \pc_target[31][17] ), .ZN(n3235) );
  OAI221_X1 U5131 ( .B1(n584), .B2(n2258), .C1(n550), .C2(n2259), .A(n3236), 
        .ZN(n3231) );
  AOI22_X1 U5132 ( .A1(n2261), .A2(\pc_target[18][17] ), .B1(n2262), .B2(
        \pc_target[19][17] ), .ZN(n3236) );
  OAI221_X1 U5135 ( .B1(n378), .B2(n2263), .C1(n343), .C2(n2264), .A(n3237), 
        .ZN(n3230) );
  AOI22_X1 U5136 ( .A1(n2266), .A2(\pc_target[20][17] ), .B1(n2267), .B2(
        \pc_target[21][17] ), .ZN(n3237) );
  NOR4_X1 U5139 ( .A1(n3238), .A2(n3239), .A3(n3240), .A4(n3241), .ZN(n3228)
         );
  OAI221_X1 U5140 ( .B1(n861), .B2(n2272), .C1(n827), .C2(n2273), .A(n3242), 
        .ZN(n3241) );
  AOI22_X1 U5141 ( .A1(n2275), .A2(\pc_target[10][17] ), .B1(n2276), .B2(
        \pc_target[11][17] ), .ZN(n3242) );
  OAI221_X1 U5144 ( .B1(n723), .B2(n2277), .C1(n689), .C2(n2278), .A(n3243), 
        .ZN(n3240) );
  AOI22_X1 U5145 ( .A1(n2280), .A2(\pc_target[14][17] ), .B1(n2281), .B2(
        \pc_target[15][17] ), .ZN(n3243) );
  OAI221_X1 U5148 ( .B1(n1135), .B2(n2282), .C1(n1101), .C2(n2283), .A(n3244), 
        .ZN(n3239) );
  AOI22_X1 U5149 ( .A1(n2285), .A2(\pc_target[2][17] ), .B1(n2286), .B2(
        \pc_target[3][17] ), .ZN(n3244) );
  OAI221_X1 U5152 ( .B1(n998), .B2(n2287), .C1(n964), .C2(n2288), .A(n3245), 
        .ZN(n3238) );
  AOI22_X1 U5153 ( .A1(n2290), .A2(\pc_target[6][17] ), .B1(n2291), .B2(
        \pc_target[7][17] ), .ZN(n3245) );
  NAND2_X1 U5156 ( .A1(n3246), .A2(n3247), .ZN(N109) );
  NOR4_X1 U5157 ( .A1(n3248), .A2(n3249), .A3(n3250), .A4(n3251), .ZN(n3247)
         );
  OAI221_X1 U5158 ( .B1(n290), .B2(n2248), .C1(n256), .C2(n2249), .A(n3252), 
        .ZN(n3251) );
  AOI22_X1 U5159 ( .A1(n2251), .A2(\pc_target[26][18] ), .B1(n2252), .B2(
        \pc_target[27][18] ), .ZN(n3252) );
  OAI221_X1 U5162 ( .B1(n150), .B2(n2253), .C1(n90), .C2(n2254), .A(n3253), 
        .ZN(n3250) );
  AOI22_X1 U5163 ( .A1(n2256), .A2(\pc_target[30][18] ), .B1(n2257), .B2(
        \pc_target[31][18] ), .ZN(n3253) );
  OAI221_X1 U5166 ( .B1(n566), .B2(n2258), .C1(n532), .C2(n2259), .A(n3254), 
        .ZN(n3249) );
  AOI22_X1 U5167 ( .A1(n2261), .A2(\pc_target[18][18] ), .B1(n2262), .B2(
        \pc_target[19][18] ), .ZN(n3254) );
  OAI221_X1 U5170 ( .B1(n360), .B2(n2263), .C1(n325), .C2(n2264), .A(n3255), 
        .ZN(n3248) );
  AOI22_X1 U5171 ( .A1(n2266), .A2(\pc_target[20][18] ), .B1(n2267), .B2(
        \pc_target[21][18] ), .ZN(n3255) );
  NOR4_X1 U5174 ( .A1(n3256), .A2(n3257), .A3(n3258), .A4(n3259), .ZN(n3246)
         );
  OAI221_X1 U5175 ( .B1(n843), .B2(n2272), .C1(n809), .C2(n2273), .A(n3260), 
        .ZN(n3259) );
  AOI22_X1 U5176 ( .A1(n2275), .A2(\pc_target[10][18] ), .B1(n2276), .B2(
        \pc_target[11][18] ), .ZN(n3260) );
  OAI221_X1 U5179 ( .B1(n705), .B2(n2277), .C1(n671), .C2(n2278), .A(n3261), 
        .ZN(n3258) );
  AOI22_X1 U5180 ( .A1(n2280), .A2(\pc_target[14][18] ), .B1(n2281), .B2(
        \pc_target[15][18] ), .ZN(n3261) );
  OAI221_X1 U5183 ( .B1(n1117), .B2(n2282), .C1(n1083), .C2(n2283), .A(n3262), 
        .ZN(n3257) );
  AOI22_X1 U5184 ( .A1(n2285), .A2(\pc_target[2][18] ), .B1(n2286), .B2(
        \pc_target[3][18] ), .ZN(n3262) );
  OAI221_X1 U5187 ( .B1(n980), .B2(n2287), .C1(n946), .C2(n2288), .A(n3263), 
        .ZN(n3256) );
  AOI22_X1 U5188 ( .A1(n2290), .A2(\pc_target[6][18] ), .B1(n2291), .B2(
        \pc_target[7][18] ), .ZN(n3263) );
  NAND2_X1 U5191 ( .A1(n3264), .A2(n3265), .ZN(N108) );
  NOR4_X1 U5192 ( .A1(n3266), .A2(n3267), .A3(n3268), .A4(n3269), .ZN(n3265)
         );
  OAI221_X1 U5193 ( .B1(n309), .B2(n2248), .C1(n275), .C2(n2249), .A(n3270), 
        .ZN(n3269) );
  AOI22_X1 U5194 ( .A1(n2251), .A2(\pc_target[26][19] ), .B1(n2252), .B2(
        \pc_target[27][19] ), .ZN(n3270) );
  OAI221_X1 U5197 ( .B1(n169), .B2(n2253), .C1(n128), .C2(n2254), .A(n3271), 
        .ZN(n3268) );
  AOI22_X1 U5198 ( .A1(n2256), .A2(\pc_target[30][19] ), .B1(n2257), .B2(
        \pc_target[31][19] ), .ZN(n3271) );
  OAI221_X1 U5201 ( .B1(n585), .B2(n2258), .C1(n551), .C2(n2259), .A(n3272), 
        .ZN(n3267) );
  AOI22_X1 U5202 ( .A1(n2261), .A2(\pc_target[18][19] ), .B1(n2262), .B2(
        \pc_target[19][19] ), .ZN(n3272) );
  OAI221_X1 U5205 ( .B1(n379), .B2(n2263), .C1(n344), .C2(n2264), .A(n3273), 
        .ZN(n3266) );
  AOI22_X1 U5206 ( .A1(n2266), .A2(\pc_target[20][19] ), .B1(n2267), .B2(
        \pc_target[21][19] ), .ZN(n3273) );
  NOR4_X1 U5209 ( .A1(n3274), .A2(n3275), .A3(n3276), .A4(n3277), .ZN(n3264)
         );
  OAI221_X1 U5210 ( .B1(n862), .B2(n2272), .C1(n828), .C2(n2273), .A(n3278), 
        .ZN(n3277) );
  AOI22_X1 U5211 ( .A1(n2275), .A2(\pc_target[10][19] ), .B1(n2276), .B2(
        \pc_target[11][19] ), .ZN(n3278) );
  OAI221_X1 U5214 ( .B1(n724), .B2(n2277), .C1(n690), .C2(n2278), .A(n3279), 
        .ZN(n3276) );
  AOI22_X1 U5215 ( .A1(n2280), .A2(\pc_target[14][19] ), .B1(n2281), .B2(
        \pc_target[15][19] ), .ZN(n3279) );
  OAI221_X1 U5218 ( .B1(n1136), .B2(n2282), .C1(n1102), .C2(n2283), .A(n3280), 
        .ZN(n3275) );
  AOI22_X1 U5219 ( .A1(n2285), .A2(\pc_target[2][19] ), .B1(n2286), .B2(
        \pc_target[3][19] ), .ZN(n3280) );
  OAI221_X1 U5222 ( .B1(n999), .B2(n2287), .C1(n965), .C2(n2288), .A(n3281), 
        .ZN(n3274) );
  AOI22_X1 U5223 ( .A1(n2290), .A2(\pc_target[6][19] ), .B1(n2291), .B2(
        \pc_target[7][19] ), .ZN(n3281) );
  NAND2_X1 U5226 ( .A1(n3282), .A2(n3283), .ZN(N107) );
  NOR4_X1 U5227 ( .A1(n3284), .A2(n3285), .A3(n3286), .A4(n3287), .ZN(n3283)
         );
  OAI221_X1 U5228 ( .B1(n289), .B2(n2248), .C1(n255), .C2(n2249), .A(n3288), 
        .ZN(n3287) );
  AOI22_X1 U5229 ( .A1(n2251), .A2(\pc_target[26][20] ), .B1(n2252), .B2(
        \pc_target[27][20] ), .ZN(n3288) );
  OAI221_X1 U5232 ( .B1(n149), .B2(n2253), .C1(n88), .C2(n2254), .A(n3289), 
        .ZN(n3286) );
  AOI22_X1 U5233 ( .A1(n2256), .A2(\pc_target[30][20] ), .B1(n2257), .B2(
        \pc_target[31][20] ), .ZN(n3289) );
  OAI221_X1 U5236 ( .B1(n565), .B2(n2258), .C1(n531), .C2(n2259), .A(n3290), 
        .ZN(n3285) );
  AOI22_X1 U5237 ( .A1(n2261), .A2(\pc_target[18][20] ), .B1(n2262), .B2(
        \pc_target[19][20] ), .ZN(n3290) );
  OAI221_X1 U5240 ( .B1(n359), .B2(n2263), .C1(n324), .C2(n2264), .A(n3291), 
        .ZN(n3284) );
  AOI22_X1 U5241 ( .A1(n2266), .A2(\pc_target[20][20] ), .B1(n2267), .B2(
        \pc_target[21][20] ), .ZN(n3291) );
  NOR4_X1 U5244 ( .A1(n3292), .A2(n3293), .A3(n3294), .A4(n3295), .ZN(n3282)
         );
  OAI221_X1 U5245 ( .B1(n842), .B2(n2272), .C1(n808), .C2(n2273), .A(n3296), 
        .ZN(n3295) );
  AOI22_X1 U5246 ( .A1(n2275), .A2(\pc_target[10][20] ), .B1(n2276), .B2(
        \pc_target[11][20] ), .ZN(n3296) );
  OAI221_X1 U5249 ( .B1(n704), .B2(n2277), .C1(n670), .C2(n2278), .A(n3297), 
        .ZN(n3294) );
  AOI22_X1 U5250 ( .A1(n2280), .A2(\pc_target[14][20] ), .B1(n2281), .B2(
        \pc_target[15][20] ), .ZN(n3297) );
  OAI221_X1 U5253 ( .B1(n1116), .B2(n2282), .C1(n1082), .C2(n2283), .A(n3298), 
        .ZN(n3293) );
  AOI22_X1 U5254 ( .A1(n2285), .A2(\pc_target[2][20] ), .B1(n2286), .B2(
        \pc_target[3][20] ), .ZN(n3298) );
  OAI221_X1 U5257 ( .B1(n979), .B2(n2287), .C1(n945), .C2(n2288), .A(n3299), 
        .ZN(n3292) );
  AOI22_X1 U5258 ( .A1(n2290), .A2(\pc_target[6][20] ), .B1(n2291), .B2(
        \pc_target[7][20] ), .ZN(n3299) );
  NAND2_X1 U5261 ( .A1(n3300), .A2(n3301), .ZN(N106) );
  NOR4_X1 U5262 ( .A1(n3302), .A2(n3303), .A3(n3304), .A4(n3305), .ZN(n3301)
         );
  OAI221_X1 U5263 ( .B1(n310), .B2(n2248), .C1(n276), .C2(n2249), .A(n3306), 
        .ZN(n3305) );
  AOI22_X1 U5264 ( .A1(n2251), .A2(\pc_target[26][21] ), .B1(n2252), .B2(
        \pc_target[27][21] ), .ZN(n3306) );
  OAI221_X1 U5267 ( .B1(n170), .B2(n2253), .C1(n130), .C2(n2254), .A(n3307), 
        .ZN(n3304) );
  AOI22_X1 U5268 ( .A1(n2256), .A2(\pc_target[30][21] ), .B1(n2257), .B2(
        \pc_target[31][21] ), .ZN(n3307) );
  OAI221_X1 U5271 ( .B1(n586), .B2(n2258), .C1(n552), .C2(n2259), .A(n3308), 
        .ZN(n3303) );
  AOI22_X1 U5272 ( .A1(n2261), .A2(\pc_target[18][21] ), .B1(n2262), .B2(
        \pc_target[19][21] ), .ZN(n3308) );
  OAI221_X1 U5275 ( .B1(n380), .B2(n2263), .C1(n345), .C2(n2264), .A(n3309), 
        .ZN(n3302) );
  AOI22_X1 U5276 ( .A1(n2266), .A2(\pc_target[20][21] ), .B1(n2267), .B2(
        \pc_target[21][21] ), .ZN(n3309) );
  NOR4_X1 U5279 ( .A1(n3310), .A2(n3311), .A3(n3312), .A4(n3313), .ZN(n3300)
         );
  OAI221_X1 U5280 ( .B1(n863), .B2(n2272), .C1(n829), .C2(n2273), .A(n3314), 
        .ZN(n3313) );
  AOI22_X1 U5281 ( .A1(n2275), .A2(\pc_target[10][21] ), .B1(n2276), .B2(
        \pc_target[11][21] ), .ZN(n3314) );
  OAI221_X1 U5284 ( .B1(n725), .B2(n2277), .C1(n691), .C2(n2278), .A(n3315), 
        .ZN(n3312) );
  AOI22_X1 U5285 ( .A1(n2280), .A2(\pc_target[14][21] ), .B1(n2281), .B2(
        \pc_target[15][21] ), .ZN(n3315) );
  OAI221_X1 U5288 ( .B1(n1137), .B2(n2282), .C1(n1103), .C2(n2283), .A(n3316), 
        .ZN(n3311) );
  AOI22_X1 U5289 ( .A1(n2285), .A2(\pc_target[2][21] ), .B1(n2286), .B2(
        \pc_target[3][21] ), .ZN(n3316) );
  OAI221_X1 U5292 ( .B1(n1000), .B2(n2287), .C1(n966), .C2(n2288), .A(n3317), 
        .ZN(n3310) );
  AOI22_X1 U5293 ( .A1(n2290), .A2(\pc_target[6][21] ), .B1(n2291), .B2(
        \pc_target[7][21] ), .ZN(n3317) );
  NAND2_X1 U5296 ( .A1(n3318), .A2(n3319), .ZN(N105) );
  NOR4_X1 U5297 ( .A1(n3320), .A2(n3321), .A3(n3322), .A4(n3323), .ZN(n3319)
         );
  OAI221_X1 U5298 ( .B1(n288), .B2(n2248), .C1(n254), .C2(n2249), .A(n3324), 
        .ZN(n3323) );
  AOI22_X1 U5299 ( .A1(n2251), .A2(\pc_target[26][22] ), .B1(n2252), .B2(
        \pc_target[27][22] ), .ZN(n3324) );
  OAI221_X1 U5302 ( .B1(n148), .B2(n2253), .C1(n86), .C2(n2254), .A(n3325), 
        .ZN(n3322) );
  AOI22_X1 U5303 ( .A1(n2256), .A2(\pc_target[30][22] ), .B1(n2257), .B2(
        \pc_target[31][22] ), .ZN(n3325) );
  OAI221_X1 U5306 ( .B1(n564), .B2(n2258), .C1(n530), .C2(n2259), .A(n3326), 
        .ZN(n3321) );
  AOI22_X1 U5307 ( .A1(n2261), .A2(\pc_target[18][22] ), .B1(n2262), .B2(
        \pc_target[19][22] ), .ZN(n3326) );
  OAI221_X1 U5310 ( .B1(n358), .B2(n2263), .C1(n323), .C2(n2264), .A(n3327), 
        .ZN(n3320) );
  AOI22_X1 U5311 ( .A1(n2266), .A2(\pc_target[20][22] ), .B1(n2267), .B2(
        \pc_target[21][22] ), .ZN(n3327) );
  NOR4_X1 U5314 ( .A1(n3328), .A2(n3329), .A3(n3330), .A4(n3331), .ZN(n3318)
         );
  OAI221_X1 U5315 ( .B1(n841), .B2(n2272), .C1(n807), .C2(n2273), .A(n3332), 
        .ZN(n3331) );
  AOI22_X1 U5316 ( .A1(n2275), .A2(\pc_target[10][22] ), .B1(n2276), .B2(
        \pc_target[11][22] ), .ZN(n3332) );
  OAI221_X1 U5319 ( .B1(n703), .B2(n2277), .C1(n669), .C2(n2278), .A(n3333), 
        .ZN(n3330) );
  AOI22_X1 U5320 ( .A1(n2280), .A2(\pc_target[14][22] ), .B1(n2281), .B2(
        \pc_target[15][22] ), .ZN(n3333) );
  OAI221_X1 U5323 ( .B1(n1115), .B2(n2282), .C1(n1081), .C2(n2283), .A(n3334), 
        .ZN(n3329) );
  AOI22_X1 U5324 ( .A1(n2285), .A2(\pc_target[2][22] ), .B1(n2286), .B2(
        \pc_target[3][22] ), .ZN(n3334) );
  OAI221_X1 U5327 ( .B1(n978), .B2(n2287), .C1(n944), .C2(n2288), .A(n3335), 
        .ZN(n3328) );
  AOI22_X1 U5328 ( .A1(n2290), .A2(\pc_target[6][22] ), .B1(n2291), .B2(
        \pc_target[7][22] ), .ZN(n3335) );
  NAND2_X1 U5331 ( .A1(n3336), .A2(n3337), .ZN(N104) );
  NOR4_X1 U5332 ( .A1(n3338), .A2(n3339), .A3(n3340), .A4(n3341), .ZN(n3337)
         );
  OAI221_X1 U5333 ( .B1(n311), .B2(n2248), .C1(n277), .C2(n2249), .A(n3342), 
        .ZN(n3341) );
  AOI22_X1 U5334 ( .A1(n2251), .A2(\pc_target[26][23] ), .B1(n2252), .B2(
        \pc_target[27][23] ), .ZN(n3342) );
  OAI221_X1 U5337 ( .B1(n171), .B2(n2253), .C1(n132), .C2(n2254), .A(n3343), 
        .ZN(n3340) );
  AOI22_X1 U5338 ( .A1(n2256), .A2(\pc_target[30][23] ), .B1(n2257), .B2(
        \pc_target[31][23] ), .ZN(n3343) );
  OAI221_X1 U5341 ( .B1(n587), .B2(n2258), .C1(n553), .C2(n2259), .A(n3344), 
        .ZN(n3339) );
  AOI22_X1 U5342 ( .A1(n2261), .A2(\pc_target[18][23] ), .B1(n2262), .B2(
        \pc_target[19][23] ), .ZN(n3344) );
  OAI221_X1 U5345 ( .B1(n381), .B2(n2263), .C1(n346), .C2(n2264), .A(n3345), 
        .ZN(n3338) );
  AOI22_X1 U5346 ( .A1(n2266), .A2(\pc_target[20][23] ), .B1(n2267), .B2(
        \pc_target[21][23] ), .ZN(n3345) );
  NOR4_X1 U5349 ( .A1(n3346), .A2(n3347), .A3(n3348), .A4(n3349), .ZN(n3336)
         );
  OAI221_X1 U5350 ( .B1(n864), .B2(n2272), .C1(n830), .C2(n2273), .A(n3350), 
        .ZN(n3349) );
  AOI22_X1 U5351 ( .A1(n2275), .A2(\pc_target[10][23] ), .B1(n2276), .B2(
        \pc_target[11][23] ), .ZN(n3350) );
  OAI221_X1 U5354 ( .B1(n726), .B2(n2277), .C1(n692), .C2(n2278), .A(n3351), 
        .ZN(n3348) );
  AOI22_X1 U5355 ( .A1(n2280), .A2(\pc_target[14][23] ), .B1(n2281), .B2(
        \pc_target[15][23] ), .ZN(n3351) );
  OAI221_X1 U5358 ( .B1(n1138), .B2(n2282), .C1(n1104), .C2(n2283), .A(n3352), 
        .ZN(n3347) );
  AOI22_X1 U5359 ( .A1(n2285), .A2(\pc_target[2][23] ), .B1(n2286), .B2(
        \pc_target[3][23] ), .ZN(n3352) );
  OAI221_X1 U5362 ( .B1(n1001), .B2(n2287), .C1(n967), .C2(n2288), .A(n3353), 
        .ZN(n3346) );
  AOI22_X1 U5363 ( .A1(n2290), .A2(\pc_target[6][23] ), .B1(n2291), .B2(
        \pc_target[7][23] ), .ZN(n3353) );
  NAND2_X1 U5366 ( .A1(n3354), .A2(n3355), .ZN(N103) );
  NOR4_X1 U5367 ( .A1(n3356), .A2(n3357), .A3(n3358), .A4(n3359), .ZN(n3355)
         );
  OAI221_X1 U5368 ( .B1(n287), .B2(n2248), .C1(n253), .C2(n2249), .A(n3360), 
        .ZN(n3359) );
  AOI22_X1 U5369 ( .A1(n2251), .A2(\pc_target[26][24] ), .B1(n2252), .B2(
        \pc_target[27][24] ), .ZN(n3360) );
  OAI221_X1 U5372 ( .B1(n147), .B2(n2253), .C1(n84), .C2(n2254), .A(n3361), 
        .ZN(n3358) );
  AOI22_X1 U5373 ( .A1(n2256), .A2(\pc_target[30][24] ), .B1(n2257), .B2(
        \pc_target[31][24] ), .ZN(n3361) );
  OAI221_X1 U5376 ( .B1(n563), .B2(n2258), .C1(n529), .C2(n2259), .A(n3362), 
        .ZN(n3357) );
  AOI22_X1 U5377 ( .A1(n2261), .A2(\pc_target[18][24] ), .B1(n2262), .B2(
        \pc_target[19][24] ), .ZN(n3362) );
  OAI221_X1 U5380 ( .B1(n357), .B2(n2263), .C1(n322), .C2(n2264), .A(n3363), 
        .ZN(n3356) );
  AOI22_X1 U5381 ( .A1(n2266), .A2(\pc_target[20][24] ), .B1(n2267), .B2(
        \pc_target[21][24] ), .ZN(n3363) );
  NOR4_X1 U5384 ( .A1(n3364), .A2(n3365), .A3(n3366), .A4(n3367), .ZN(n3354)
         );
  OAI221_X1 U5385 ( .B1(n840), .B2(n2272), .C1(n806), .C2(n2273), .A(n3368), 
        .ZN(n3367) );
  AOI22_X1 U5386 ( .A1(n2275), .A2(\pc_target[10][24] ), .B1(n2276), .B2(
        \pc_target[11][24] ), .ZN(n3368) );
  OAI221_X1 U5389 ( .B1(n702), .B2(n2277), .C1(n668), .C2(n2278), .A(n3369), 
        .ZN(n3366) );
  AOI22_X1 U5390 ( .A1(n2280), .A2(\pc_target[14][24] ), .B1(n2281), .B2(
        \pc_target[15][24] ), .ZN(n3369) );
  OAI221_X1 U5393 ( .B1(n1114), .B2(n2282), .C1(n1080), .C2(n2283), .A(n3370), 
        .ZN(n3365) );
  AOI22_X1 U5394 ( .A1(n2285), .A2(\pc_target[2][24] ), .B1(n2286), .B2(
        \pc_target[3][24] ), .ZN(n3370) );
  OAI221_X1 U5397 ( .B1(n977), .B2(n2287), .C1(n943), .C2(n2288), .A(n3371), 
        .ZN(n3364) );
  AOI22_X1 U5398 ( .A1(n2290), .A2(\pc_target[6][24] ), .B1(n2291), .B2(
        \pc_target[7][24] ), .ZN(n3371) );
  NAND2_X1 U5401 ( .A1(n3372), .A2(n3373), .ZN(N102) );
  NOR4_X1 U5402 ( .A1(n3374), .A2(n3375), .A3(n3376), .A4(n3377), .ZN(n3373)
         );
  OAI221_X1 U5403 ( .B1(n312), .B2(n2248), .C1(n278), .C2(n2249), .A(n3378), 
        .ZN(n3377) );
  AOI22_X1 U5404 ( .A1(n2251), .A2(\pc_target[26][25] ), .B1(n2252), .B2(
        \pc_target[27][25] ), .ZN(n3378) );
  OAI221_X1 U5407 ( .B1(n172), .B2(n2253), .C1(n134), .C2(n2254), .A(n3379), 
        .ZN(n3376) );
  AOI22_X1 U5408 ( .A1(n2256), .A2(\pc_target[30][25] ), .B1(n2257), .B2(
        \pc_target[31][25] ), .ZN(n3379) );
  OAI221_X1 U5411 ( .B1(n588), .B2(n2258), .C1(n554), .C2(n2259), .A(n3380), 
        .ZN(n3375) );
  AOI22_X1 U5412 ( .A1(n2261), .A2(\pc_target[18][25] ), .B1(n2262), .B2(
        \pc_target[19][25] ), .ZN(n3380) );
  OAI221_X1 U5415 ( .B1(n382), .B2(n2263), .C1(n347), .C2(n2264), .A(n3381), 
        .ZN(n3374) );
  AOI22_X1 U5416 ( .A1(n2266), .A2(\pc_target[20][25] ), .B1(n2267), .B2(
        \pc_target[21][25] ), .ZN(n3381) );
  NOR4_X1 U5419 ( .A1(n3382), .A2(n3383), .A3(n3384), .A4(n3385), .ZN(n3372)
         );
  OAI221_X1 U5420 ( .B1(n865), .B2(n2272), .C1(n831), .C2(n2273), .A(n3386), 
        .ZN(n3385) );
  AOI22_X1 U5421 ( .A1(n2275), .A2(\pc_target[10][25] ), .B1(n2276), .B2(
        \pc_target[11][25] ), .ZN(n3386) );
  OAI221_X1 U5424 ( .B1(n727), .B2(n2277), .C1(n693), .C2(n2278), .A(n3387), 
        .ZN(n3384) );
  AOI22_X1 U5425 ( .A1(n2280), .A2(\pc_target[14][25] ), .B1(n2281), .B2(
        \pc_target[15][25] ), .ZN(n3387) );
  OAI221_X1 U5428 ( .B1(n1139), .B2(n2282), .C1(n1105), .C2(n2283), .A(n3388), 
        .ZN(n3383) );
  AOI22_X1 U5429 ( .A1(n2285), .A2(\pc_target[2][25] ), .B1(n2286), .B2(
        \pc_target[3][25] ), .ZN(n3388) );
  OAI221_X1 U5432 ( .B1(n1002), .B2(n2287), .C1(n968), .C2(n2288), .A(n3389), 
        .ZN(n3382) );
  AOI22_X1 U5433 ( .A1(n2290), .A2(\pc_target[6][25] ), .B1(n2291), .B2(
        \pc_target[7][25] ), .ZN(n3389) );
  NAND2_X1 U5436 ( .A1(n3390), .A2(n3391), .ZN(N101) );
  NOR4_X1 U5437 ( .A1(n3392), .A2(n3393), .A3(n3394), .A4(n3395), .ZN(n3391)
         );
  OAI221_X1 U5438 ( .B1(n286), .B2(n2248), .C1(n252), .C2(n2249), .A(n3396), 
        .ZN(n3395) );
  AOI22_X1 U5439 ( .A1(n2251), .A2(\pc_target[26][26] ), .B1(n2252), .B2(
        \pc_target[27][26] ), .ZN(n3396) );
  OAI221_X1 U5442 ( .B1(n146), .B2(n2253), .C1(n82), .C2(n2254), .A(n3397), 
        .ZN(n3394) );
  AOI22_X1 U5443 ( .A1(n2256), .A2(\pc_target[30][26] ), .B1(n2257), .B2(
        \pc_target[31][26] ), .ZN(n3397) );
  OAI221_X1 U5446 ( .B1(n562), .B2(n2258), .C1(n528), .C2(n2259), .A(n3398), 
        .ZN(n3393) );
  AOI22_X1 U5447 ( .A1(n2261), .A2(\pc_target[18][26] ), .B1(n2262), .B2(
        \pc_target[19][26] ), .ZN(n3398) );
  OAI221_X1 U5450 ( .B1(n356), .B2(n2263), .C1(n321), .C2(n2264), .A(n3399), 
        .ZN(n3392) );
  AOI22_X1 U5451 ( .A1(n2266), .A2(\pc_target[20][26] ), .B1(n2267), .B2(
        \pc_target[21][26] ), .ZN(n3399) );
  NOR4_X1 U5454 ( .A1(n3400), .A2(n3401), .A3(n3402), .A4(n3403), .ZN(n3390)
         );
  OAI221_X1 U5455 ( .B1(n839), .B2(n2272), .C1(n805), .C2(n2273), .A(n3404), 
        .ZN(n3403) );
  AOI22_X1 U5456 ( .A1(n2275), .A2(\pc_target[10][26] ), .B1(n2276), .B2(
        \pc_target[11][26] ), .ZN(n3404) );
  OAI221_X1 U5459 ( .B1(n701), .B2(n2277), .C1(n667), .C2(n2278), .A(n3405), 
        .ZN(n3402) );
  AOI22_X1 U5460 ( .A1(n2280), .A2(\pc_target[14][26] ), .B1(n2281), .B2(
        \pc_target[15][26] ), .ZN(n3405) );
  OAI221_X1 U5463 ( .B1(n1113), .B2(n2282), .C1(n1079), .C2(n2283), .A(n3406), 
        .ZN(n3401) );
  AOI22_X1 U5464 ( .A1(n2285), .A2(\pc_target[2][26] ), .B1(n2286), .B2(
        \pc_target[3][26] ), .ZN(n3406) );
  OAI221_X1 U5467 ( .B1(n976), .B2(n2287), .C1(n942), .C2(n2288), .A(n3407), 
        .ZN(n3400) );
  AOI22_X1 U5468 ( .A1(n2290), .A2(\pc_target[6][26] ), .B1(n2291), .B2(
        \pc_target[7][26] ), .ZN(n3407) );
  NAND2_X1 U5471 ( .A1(n3408), .A2(n3409), .ZN(N100) );
  NOR4_X1 U5472 ( .A1(n3410), .A2(n3411), .A3(n3412), .A4(n3413), .ZN(n3409)
         );
  OAI221_X1 U5473 ( .B1(n313), .B2(n2248), .C1(n279), .C2(n2249), .A(n3414), 
        .ZN(n3413) );
  AOI22_X1 U5474 ( .A1(n2251), .A2(\pc_target[26][27] ), .B1(n2252), .B2(
        \pc_target[27][27] ), .ZN(n3414) );
  OAI221_X1 U5481 ( .B1(n173), .B2(n2253), .C1(n136), .C2(n2254), .A(n3419), 
        .ZN(n3412) );
  AOI22_X1 U5482 ( .A1(n2256), .A2(\pc_target[30][27] ), .B1(n2257), .B2(
        \pc_target[31][27] ), .ZN(n3419) );
  AND3_X1 U5486 ( .A1(PC_read[0]), .A2(PC_read[4]), .A3(PC_read[3]), .ZN(n3415) );
  AND3_X1 U5489 ( .A1(PC_read[4]), .A2(n3422), .A3(PC_read[3]), .ZN(n3417) );
  OAI221_X1 U5491 ( .B1(n589), .B2(n2258), .C1(n555), .C2(n2259), .A(n3423), 
        .ZN(n3411) );
  AOI22_X1 U5492 ( .A1(n2261), .A2(\pc_target[18][27] ), .B1(n2262), .B2(
        \pc_target[19][27] ), .ZN(n3423) );
  OAI221_X1 U5499 ( .B1(n383), .B2(n2263), .C1(n348), .C2(n2264), .A(n3426), 
        .ZN(n3410) );
  AOI22_X1 U5500 ( .A1(n2266), .A2(\pc_target[20][27] ), .B1(n2267), .B2(
        \pc_target[21][27] ), .ZN(n3426) );
  AND3_X1 U5504 ( .A1(PC_read[4]), .A2(n3427), .A3(PC_read[0]), .ZN(n3424) );
  AND3_X1 U5507 ( .A1(n3422), .A2(n3427), .A3(PC_read[4]), .ZN(n3425) );
  NOR4_X1 U5509 ( .A1(n3428), .A2(n3429), .A3(n3430), .A4(n3431), .ZN(n3408)
         );
  OAI221_X1 U5510 ( .B1(n866), .B2(n2272), .C1(n832), .C2(n2273), .A(n3432), 
        .ZN(n3431) );
  AOI22_X1 U5511 ( .A1(n2275), .A2(\pc_target[10][27] ), .B1(n2276), .B2(
        \pc_target[11][27] ), .ZN(n3432) );
  OAI221_X1 U5518 ( .B1(n728), .B2(n2277), .C1(n694), .C2(n2278), .A(n3435), 
        .ZN(n3430) );
  AOI22_X1 U5519 ( .A1(n2280), .A2(\pc_target[14][27] ), .B1(n2281), .B2(
        \pc_target[15][27] ), .ZN(n3435) );
  INV_X1 U5527 ( .A(PC_read[3]), .ZN(n3427) );
  OAI221_X1 U5529 ( .B1(n1140), .B2(n2282), .C1(n1106), .C2(n2283), .A(n3436), 
        .ZN(n3429) );
  AOI22_X1 U5530 ( .A1(n2285), .A2(\pc_target[2][27] ), .B1(n2286), .B2(
        \pc_target[3][27] ), .ZN(n3436) );
  OAI221_X1 U5539 ( .B1(n1003), .B2(n2287), .C1(n969), .C2(n2288), .A(n3440), 
        .ZN(n3428) );
  AOI22_X1 U5540 ( .A1(n2290), .A2(\pc_target[6][27] ), .B1(n2291), .B2(
        \pc_target[7][27] ), .ZN(n3440) );
  INV_X1 U5544 ( .A(PC_read[1]), .ZN(n3439) );
  INV_X1 U5547 ( .A(PC_read[0]), .ZN(n3422) );
  INV_X1 U5551 ( .A(PC_read[2]), .ZN(n3441) );
  DFFR_X2 \pc_target_reg[6][30]  ( .D(n6290), .CK(Clk), .RN(n3824), .Q(
        \pc_target[6][30] ) );
  DFFR_X2 \pc_target_reg[6][28]  ( .D(n6291), .CK(Clk), .RN(n3825), .Q(
        \pc_target[6][28] ) );
  DFFR_X2 \pc_target_reg[6][26]  ( .D(n6292), .CK(Clk), .RN(n3824), .Q(
        \pc_target[6][26] ) );
  DFFR_X2 \pc_target_reg[6][24]  ( .D(n6293), .CK(Clk), .RN(n3823), .Q(
        \pc_target[6][24] ) );
  DFFR_X2 \pc_target_reg[6][22]  ( .D(n6294), .CK(Clk), .RN(n3825), .Q(
        \pc_target[6][22] ) );
  DFFR_X2 \pc_target_reg[6][20]  ( .D(n6295), .CK(Clk), .RN(n3825), .Q(
        \pc_target[6][20] ) );
  DFFR_X2 \pc_target_reg[6][18]  ( .D(n6296), .CK(Clk), .RN(n3825), .Q(
        \pc_target[6][18] ) );
  DFFR_X2 \pc_target_reg[6][16]  ( .D(n6297), .CK(Clk), .RN(n3824), .Q(
        \pc_target[6][16] ) );
  DFFR_X2 \pc_target_reg[6][14]  ( .D(n6298), .CK(Clk), .RN(n3825), .Q(
        \pc_target[6][14] ) );
  DFFR_X2 \pc_target_reg[6][12]  ( .D(n6299), .CK(Clk), .RN(n3825), .Q(
        \pc_target[6][12] ) );
  DFFR_X2 \pc_target_reg[6][10]  ( .D(n6300), .CK(Clk), .RN(n3824), .Q(
        \pc_target[6][10] ) );
  DFFR_X2 \pc_target_reg[6][8]  ( .D(n6301), .CK(Clk), .RN(n3825), .Q(
        \pc_target[6][8] ) );
  DFFR_X2 \pc_target_reg[6][6]  ( .D(n6302), .CK(Clk), .RN(n3823), .Q(
        \pc_target[6][6] ) );
  DFFR_X2 \pc_target_reg[6][4]  ( .D(n6303), .CK(Clk), .RN(n3824), .Q(
        \pc_target[6][4] ) );
  DFFR_X2 \pc_target_reg[6][2]  ( .D(n6304), .CK(Clk), .RN(n3825), .Q(
        \pc_target[6][2] ) );
  DFFR_X2 \pc_target_reg[6][0]  ( .D(n6305), .CK(Clk), .RN(n3824), .Q(
        \pc_target[6][0] ) );
  DFFR_X2 \pc_target_reg[6][1]  ( .D(n6306), .CK(Clk), .RN(n3824), .Q(
        \pc_target[6][1] ) );
  DFFR_X2 \pc_target_reg[6][3]  ( .D(n6307), .CK(Clk), .RN(n3824), .Q(
        \pc_target[6][3] ) );
  DFFR_X2 \pc_target_reg[6][5]  ( .D(n6308), .CK(Clk), .RN(n3825), .Q(
        \pc_target[6][5] ) );
  DFFR_X2 \pc_target_reg[6][7]  ( .D(n6309), .CK(Clk), .RN(n3826), .Q(
        \pc_target[6][7] ) );
  DFFR_X2 \pc_target_reg[6][9]  ( .D(n6310), .CK(Clk), .RN(n3824), .Q(
        \pc_target[6][9] ) );
  DFFR_X2 \pc_target_reg[6][11]  ( .D(n6311), .CK(Clk), .RN(n3826), .Q(
        \pc_target[6][11] ) );
  DFFR_X2 \pc_target_reg[6][13]  ( .D(n6312), .CK(Clk), .RN(n3826), .Q(
        \pc_target[6][13] ) );
  DFFR_X2 \pc_target_reg[6][15]  ( .D(n6313), .CK(Clk), .RN(n3824), .Q(
        \pc_target[6][15] ) );
  DFFR_X2 \pc_target_reg[6][17]  ( .D(n6314), .CK(Clk), .RN(n3824), .Q(
        \pc_target[6][17] ) );
  DFFR_X2 \pc_target_reg[6][19]  ( .D(n6315), .CK(Clk), .RN(n3826), .Q(
        \pc_target[6][19] ) );
  DFFR_X2 \pc_target_reg[6][21]  ( .D(n6316), .CK(Clk), .RN(n3825), .Q(
        \pc_target[6][21] ) );
  DFFR_X2 \pc_target_reg[6][23]  ( .D(n6317), .CK(Clk), .RN(n3826), .Q(
        \pc_target[6][23] ) );
  DFFR_X2 \pc_target_reg[6][25]  ( .D(n6318), .CK(Clk), .RN(n3826), .Q(
        \pc_target[6][25] ) );
  DFFR_X2 \pc_target_reg[6][27]  ( .D(n6319), .CK(Clk), .RN(n3825), .Q(
        \pc_target[6][27] ) );
  DFFR_X2 \pc_target_reg[6][29]  ( .D(n6320), .CK(Clk), .RN(n3825), .Q(
        \pc_target[6][29] ) );
  DFFR_X2 \pc_target_reg[6][31]  ( .D(n6321), .CK(Clk), .RN(n3822), .Q(
        \pc_target[6][31] ) );
  DFFR_X2 \pc_target_reg[2][30]  ( .D(n6418), .CK(Clk), .RN(n3822), .Q(
        \pc_target[2][30] ) );
  DFFR_X2 \pc_target_reg[2][28]  ( .D(n6419), .CK(Clk), .RN(n3822), .Q(
        \pc_target[2][28] ) );
  DFFR_X2 \pc_target_reg[2][26]  ( .D(n6420), .CK(Clk), .RN(n3822), .Q(
        \pc_target[2][26] ) );
  DFFR_X2 \pc_target_reg[2][24]  ( .D(n6421), .CK(Clk), .RN(n3822), .Q(
        \pc_target[2][24] ) );
  DFFR_X2 \pc_target_reg[2][22]  ( .D(n6422), .CK(Clk), .RN(n3822), .Q(
        \pc_target[2][22] ) );
  DFFR_X2 \pc_target_reg[2][20]  ( .D(n6423), .CK(Clk), .RN(n3822), .Q(
        \pc_target[2][20] ) );
  DFFR_X2 \pc_target_reg[2][18]  ( .D(n6424), .CK(Clk), .RN(n3822), .Q(
        \pc_target[2][18] ) );
  DFFR_X2 \pc_target_reg[2][16]  ( .D(n6425), .CK(Clk), .RN(n3822), .Q(
        \pc_target[2][16] ) );
  DFFR_X2 \pc_target_reg[2][14]  ( .D(n6426), .CK(Clk), .RN(n3822), .Q(
        \pc_target[2][14] ) );
  DFFR_X2 \pc_target_reg[2][12]  ( .D(n6427), .CK(Clk), .RN(n3822), .Q(
        \pc_target[2][12] ) );
  DFFR_X2 \pc_target_reg[2][7]  ( .D(n6437), .CK(Clk), .RN(n3823), .Q(
        \pc_target[2][7] ) );
  DFFR_X2 \pc_target_reg[2][11]  ( .D(n6439), .CK(Clk), .RN(n3823), .Q(
        \pc_target[2][11] ) );
  DFFR_X2 \pc_target_reg[2][13]  ( .D(n6440), .CK(Clk), .RN(n3823), .Q(
        \pc_target[2][13] ) );
  DFFR_X2 \pc_target_reg[2][15]  ( .D(n6441), .CK(Clk), .RN(n3822), .Q(
        \pc_target[2][15] ) );
  DFFR_X2 \pc_target_reg[2][17]  ( .D(n6442), .CK(Clk), .RN(n3823), .Q(
        \pc_target[2][17] ) );
  DFFR_X2 \pc_target_reg[2][19]  ( .D(n6443), .CK(Clk), .RN(n3823), .Q(
        \pc_target[2][19] ) );
  DFFR_X2 \pc_target_reg[2][21]  ( .D(n6444), .CK(Clk), .RN(n3823), .Q(
        \pc_target[2][21] ) );
  DFFR_X2 \pc_target_reg[2][23]  ( .D(n6445), .CK(Clk), .RN(n3823), .Q(
        \pc_target[2][23] ) );
  DFFR_X2 \pc_target_reg[2][25]  ( .D(n6446), .CK(Clk), .RN(n3823), .Q(
        \pc_target[2][25] ) );
  DFFR_X2 \pc_target_reg[2][27]  ( .D(n6447), .CK(Clk), .RN(n3823), .Q(
        \pc_target[2][27] ) );
  DFFR_X2 \pc_target_reg[2][29]  ( .D(n6448), .CK(Clk), .RN(n3824), .Q(
        \pc_target[2][29] ) );
  DFFR_X2 \pc_target_reg[2][31]  ( .D(n6449), .CK(Clk), .RN(n3823), .Q(
        \pc_target[2][31] ) );
  DFFR_X1 \pc_target_reg[2][6]  ( .D(n6430), .CK(Clk), .RN(n3910), .Q(
        \pc_target[2][6] ) );
  DFFR_X1 \pc_target_reg[2][5]  ( .D(n6436), .CK(Clk), .RN(n3910), .Q(
        \pc_target[2][5] ) );
  DFFR_X1 \pc_target_reg[2][4]  ( .D(n6431), .CK(Clk), .RN(n3910), .Q(
        \pc_target[2][4] ) );
  DFFR_X1 \pc_target_reg[2][2]  ( .D(n6432), .CK(Clk), .RN(n3910), .Q(
        \pc_target[2][2] ) );
  DFFR_X1 \pc_target_reg[2][1]  ( .D(n6434), .CK(Clk), .RN(n3910), .Q(
        \pc_target[2][1] ) );
  DFFR_X1 \pc_target_reg[2][0]  ( .D(n6433), .CK(Clk), .RN(n3827), .Q(
        \pc_target[2][0] ) );
  DFFR_X1 \pc_lut_reg[14][3]  ( .D(n7075), .CK(Clk), .RN(n3911), .Q(
        \pc_lut[14][3] ) );
  DFFR_X1 \pc_lut_reg[14][2]  ( .D(n7072), .CK(Clk), .RN(n3911), .Q(
        \pc_lut[14][2] ) );
  DFFR_X1 \pc_lut_reg[14][1]  ( .D(n7074), .CK(Clk), .RN(n3911), .Q(
        \pc_lut[14][1] ) );
  DFFR_X1 \pc_lut_reg[15][3]  ( .D(n7043), .CK(Clk), .RN(n3911), .Q(
        \pc_lut[15][3] ) );
  DFFR_X1 \pc_lut_reg[15][2]  ( .D(n7040), .CK(Clk), .RN(n3912), .Q(
        \pc_lut[15][2] ) );
  DFFR_X1 \pc_lut_reg[15][1]  ( .D(n7042), .CK(Clk), .RN(n3911), .Q(
        \pc_lut[15][1] ) );
  DFFR_X1 \pc_lut_reg[15][0]  ( .D(n7041), .CK(Clk), .RN(n3912), .Q(
        \pc_lut[15][0] ) );
  DFFR_X1 \pc_lut_reg[26][4]  ( .D(n6687), .CK(Clk), .RN(n3912), .Q(
        \pc_lut[26][4] ) );
  DFFR_X1 \pc_lut_reg[26][3]  ( .D(n6691), .CK(Clk), .RN(n3912), .Q(
        \pc_lut[26][3] ) );
  DFFR_X1 \pc_lut_reg[26][1]  ( .D(n6690), .CK(Clk), .RN(n3912), .Q(
        \pc_lut[26][1] ) );
  DFFR_X1 \pc_lut_reg[28][4]  ( .D(n6623), .CK(Clk), .RN(n3912), .QN(n1290) );
  DFFR_X1 \pc_lut_reg[28][3]  ( .D(n6627), .CK(Clk), .RN(n3912), .QN(n1294) );
  DFFR_X1 \pc_lut_reg[28][2]  ( .D(n6624), .CK(Clk), .RN(n3912), .QN(n1291) );
  DFFR_X1 \pc_lut_reg[29][4]  ( .D(n6591), .CK(Clk), .RN(n3912), .QN(n1255) );
  DFFR_X1 \pc_lut_reg[29][3]  ( .D(n6595), .CK(Clk), .RN(n3912), .QN(n1260) );
  DFFR_X1 \pc_lut_reg[29][2]  ( .D(n6592), .CK(Clk), .RN(n3912), .QN(n1257) );
  DFFR_X1 \pc_lut_reg[29][0]  ( .D(n6593), .CK(Clk), .RN(n3912), .QN(n1258) );
  DFFR_X1 \pc_target_reg[24][5]  ( .D(n5732), .CK(Clk), .RN(n3910), .QN(n302)
         );
  DFFR_X1 \pc_target_reg[24][4]  ( .D(n5727), .CK(Clk), .RN(n3911), .QN(n297)
         );
  DFFR_X1 \pc_target_reg[17][5]  ( .D(n5956), .CK(Clk), .RN(n3911), .QN(n544)
         );
  DFFR_X1 \pc_target_reg[17][4]  ( .D(n5951), .CK(Clk), .RN(n3911), .QN(n539)
         );
  DFFR_X1 \pc_target_reg[9][5]  ( .D(n6212), .CK(Clk), .RN(n3908), .QN(n821)
         );
  DFFR_X1 \pc_target_reg[9][4]  ( .D(n6207), .CK(Clk), .RN(n3908), .QN(n816)
         );
  DFFR_X1 \pc_target_reg[4][5]  ( .D(n6372), .CK(Clk), .RN(n3909), .QN(n992)
         );
  DFFR_X1 \pc_target_reg[4][4]  ( .D(n6367), .CK(Clk), .RN(n3909), .QN(n987)
         );
  DFFR_X1 \pc_target_reg[2][10]  ( .D(n6428), .CK(Clk), .RN(n3910), .Q(
        \pc_target[2][10] ) );
  DFFR_X1 \pc_target_reg[2][9]  ( .D(n6438), .CK(Clk), .RN(n3910), .Q(
        \pc_target[2][9] ) );
  DFFR_X1 \pc_target_reg[2][8]  ( .D(n6429), .CK(Clk), .RN(n3910), .Q(
        \pc_target[2][8] ) );
  DFFR_X1 \pc_target_reg[10][10]  ( .D(n6172), .CK(Clk), .RN(n3908), .Q(
        \pc_target[10][10] ) );
  DFFR_X1 \pc_target_reg[10][9]  ( .D(n6182), .CK(Clk), .RN(n3908), .Q(
        \pc_target[10][9] ) );
  DFFR_X1 \pc_target_reg[10][8]  ( .D(n6173), .CK(Clk), .RN(n3908), .Q(
        \pc_target[10][8] ) );
  DFFR_X1 \pc_target_reg[10][3]  ( .D(n6179), .CK(Clk), .RN(n3908), .Q(
        \pc_target[10][3] ) );
  DFFR_X1 \pc_target_reg[15][10]  ( .D(n6012), .CK(Clk), .RN(n3909), .Q(
        \pc_target[15][10] ) );
  DFFR_X1 \pc_target_reg[15][9]  ( .D(n6022), .CK(Clk), .RN(n3909), .Q(
        \pc_target[15][9] ) );
  DFFR_X1 \pc_target_reg[15][8]  ( .D(n6013), .CK(Clk), .RN(n3909), .Q(
        \pc_target[15][8] ) );
  DFFR_X1 \pc_target_reg[15][6]  ( .D(n6014), .CK(Clk), .RN(n3909), .Q(
        \pc_target[15][6] ) );
  DFFR_X1 \pc_target_reg[15][5]  ( .D(n6020), .CK(Clk), .RN(n3909), .Q(
        \pc_target[15][5] ) );
  DFFR_X1 \pc_target_reg[15][4]  ( .D(n6015), .CK(Clk), .RN(n3909), .Q(
        \pc_target[15][4] ) );
  DFFR_X1 \pc_target_reg[15][2]  ( .D(n6016), .CK(Clk), .RN(n3909), .Q(
        \pc_target[15][2] ) );
  DFFR_X1 \pc_target_reg[15][1]  ( .D(n6018), .CK(Clk), .RN(n3909), .Q(
        \pc_target[15][1] ) );
  DFFR_X1 \pc_target_reg[15][0]  ( .D(n6017), .CK(Clk), .RN(n3912), .Q(
        \pc_target[15][0] ) );
  DFFR_X1 \pc_target_reg[15][3]  ( .D(n6019), .CK(Clk), .RN(n3909), .Q(
        \pc_target[15][3] ) );
  DFFR_X1 \pc_target_reg[2][3]  ( .D(n6435), .CK(Clk), .RN(n3910), .Q(
        \pc_target[2][3] ) );
  DFFR_X1 \pc_target_reg[3][10]  ( .D(n6396), .CK(Clk), .RN(n3910), .Q(
        \pc_target[3][10] ) );
  DFFR_X1 \pc_target_reg[3][9]  ( .D(n6406), .CK(Clk), .RN(n3909), .Q(
        \pc_target[3][9] ) );
  DFFR_X1 \pc_target_reg[3][8]  ( .D(n6397), .CK(Clk), .RN(n3910), .Q(
        \pc_target[3][8] ) );
  DFFR_X1 \pc_target_reg[3][6]  ( .D(n6398), .CK(Clk), .RN(n3910), .Q(
        \pc_target[3][6] ) );
  DFFR_X1 \pc_target_reg[3][5]  ( .D(n6404), .CK(Clk), .RN(n3909), .Q(
        \pc_target[3][5] ) );
  DFFR_X1 \pc_target_reg[3][4]  ( .D(n6399), .CK(Clk), .RN(n3910), .Q(
        \pc_target[3][4] ) );
  DFFR_X1 \pc_target_reg[3][3]  ( .D(n6403), .CK(Clk), .RN(n3909), .Q(
        \pc_target[3][3] ) );
  DFFR_X1 \pc_target_reg[3][2]  ( .D(n6400), .CK(Clk), .RN(n3910), .Q(
        \pc_target[3][2] ) );
  DFFR_X1 \pc_target_reg[3][1]  ( .D(n6402), .CK(Clk), .RN(n3909), .Q(
        \pc_target[3][1] ) );
  DFFR_X1 \pc_target_reg[3][0]  ( .D(n6401), .CK(Clk), .RN(n3921), .Q(
        \pc_target[3][0] ) );
  DFFR_X1 \pc_target_reg[21][10]  ( .D(n5820), .CK(Clk), .RN(n3911), .Q(
        \pc_target[21][10] ) );
  DFFR_X1 \pc_target_reg[21][9]  ( .D(n5830), .CK(Clk), .RN(n3911), .Q(
        \pc_target[21][9] ) );
  DFFR_X1 \pc_target_reg[21][8]  ( .D(n5821), .CK(Clk), .RN(n3911), .Q(
        \pc_target[21][8] ) );
  DFFR_X1 \pc_target_reg[21][6]  ( .D(n5822), .CK(Clk), .RN(n3911), .Q(
        \pc_target[21][6] ) );
  DFFR_X1 \pc_target_reg[21][5]  ( .D(n5828), .CK(Clk), .RN(n3911), .Q(
        \pc_target[21][5] ) );
  DFFR_X1 \pc_target_reg[21][4]  ( .D(n5823), .CK(Clk), .RN(n3911), .Q(
        \pc_target[21][4] ) );
  DFFR_X1 \pc_target_reg[24][30]  ( .D(n5714), .CK(Clk), .RN(n3911), .QN(n284)
         );
  NOR2_X1 U68 ( .A1(n2404), .A2(n2405), .ZN(n2401) );
  NOR2_X1 U69 ( .A1(n2412), .A2(n2413), .ZN(n2400) );
  INV_X1 U134 ( .A(n2419), .ZN(N215) );
  OAI21_X1 U135 ( .B1(n1393), .B2(n2249), .A(n2352), .ZN(n2351) );
  NAND2_X1 U168 ( .A1(n2252), .A2(\pc_lut[27][0] ), .ZN(n2352) );
  OAI21_X1 U169 ( .B1(n1258), .B2(n2254), .A(n2353), .ZN(n2350) );
  NAND2_X1 U202 ( .A1(n2257), .A2(\pc_lut[31][0] ), .ZN(n2353) );
  OAI21_X1 U203 ( .B1(n1657), .B2(n2259), .A(n2354), .ZN(n2349) );
  NAND2_X1 U204 ( .A1(n2262), .A2(\pc_lut[19][0] ), .ZN(n2354) );
  OAI21_X1 U269 ( .B1(n1461), .B2(n2264), .A(n2355), .ZN(n2348) );
  NAND2_X1 U270 ( .A1(n2267), .A2(\pc_lut[21][0] ), .ZN(n2355) );
  OAI21_X1 U335 ( .B1(n1927), .B2(n2273), .A(n2360), .ZN(n2359) );
  NAND2_X1 U336 ( .A1(n2276), .A2(\pc_lut[11][0] ), .ZN(n2360) );
  OAI21_X1 U369 ( .B1(n1792), .B2(n2278), .A(n2361), .ZN(n2358) );
  NAND2_X1 U370 ( .A1(n2281), .A2(\pc_lut[15][0] ), .ZN(n2361) );
  OAI21_X1 U403 ( .B1(n2191), .B2(n2283), .A(n2362), .ZN(n2357) );
  NAND2_X1 U404 ( .A1(n2286), .A2(\pc_lut[3][0] ), .ZN(n2362) );
  OAI21_X1 U405 ( .B1(n2059), .B2(n2288), .A(n2363), .ZN(n2356) );
  NAND2_X1 U438 ( .A1(n2291), .A2(\pc_lut[7][0] ), .ZN(n2363) );
  INV_X1 U439 ( .A(n2370), .ZN(n2369) );
  INV_X1 U472 ( .A(n2371), .ZN(n2368) );
  INV_X1 U473 ( .A(n2372), .ZN(n2367) );
  OAI22_X1 U538 ( .A1(n1497), .A2(n2263), .B1(n1462), .B2(n2264), .ZN(n2366)
         );
  INV_X1 U539 ( .A(n2378), .ZN(n2377) );
  INV_X1 U604 ( .A(n2379), .ZN(n2376) );
  INV_X1 U605 ( .A(n2380), .ZN(n2375) );
  INV_X1 U606 ( .A(n2381), .ZN(n2374) );
  NOR2_X1 U671 ( .A1(n2384), .A2(n2386), .ZN(n2383) );
  NOR2_X1 U672 ( .A1(n2392), .A2(n2394), .ZN(n2382) );
  INV_X2 U737 ( .A(Set_target[15]), .ZN(n123) );
  INV_X2 U738 ( .A(Set_target[13]), .ZN(n121) );
  INV_X2 U771 ( .A(Set_target[12]), .ZN(n95) );
  INV_X2 U772 ( .A(Set_target[14]), .ZN(n93) );
  INV_X2 U777 ( .A(n2210), .ZN(n2208) );
  NAND2_X4 U805 ( .A1(n2141), .A2(n176), .ZN(n2210) );
  INV_X2 U806 ( .A(n1946), .ZN(n1944) );
  INV_X2 U808 ( .A(n1676), .ZN(n1674) );
  INV_X2 U873 ( .A(n2078), .ZN(n2076) );
  INV_X2 U874 ( .A(n2176), .ZN(n2174) );
  NAND2_X4 U939 ( .A1(n2141), .A2(n141), .ZN(n2176) );
  AND2_X1 U940 ( .A1(n2141), .A2(n74), .ZN(n2) );
  INV_X1 U973 ( .A(n2), .ZN(n3) );
  INV_X1 U974 ( .A(n2), .ZN(n283) );
  NAND2_X4 U1007 ( .A1(n2010), .A2(n141), .ZN(n2044) );
  NAND2_X4 U1008 ( .A1(n1608), .A2(n141), .ZN(n1642) );
  NAND2_X4 U1009 ( .A1(n1878), .A2(n141), .ZN(n1912) );
  NAND2_X4 U1074 ( .A1(n2010), .A2(n176), .ZN(n2078) );
  NAND2_X4 U1075 ( .A1(n1878), .A2(n176), .ZN(n1946) );
  NAND2_X4 U1140 ( .A1(n1608), .A2(n176), .ZN(n1676) );
  NAND2_X4 U1174 ( .A1(n1742), .A2(n176), .ZN(n1811) );
  NOR2_X4 U1175 ( .A1(PC_write[0]), .A2(PC_write[1]), .ZN(n176) );
  AND2_X1 U1209 ( .A1(n1608), .A2(n74), .ZN(n525) );
  INV_X1 U1210 ( .A(n525), .ZN(n558) );
  INV_X1 U1275 ( .A(n525), .ZN(n768) );
  AND2_X1 U1276 ( .A1(n2141), .A2(n38), .ZN(n802) );
  INV_X1 U1341 ( .A(n802), .ZN(n871) );
  INV_X1 U1342 ( .A(n802), .ZN(n973) );
  AND2_X1 U1375 ( .A1(n1878), .A2(n74), .ZN(n1240) );
  INV_X1 U1376 ( .A(n1240), .ZN(n1256) );
  INV_X1 U1409 ( .A(n1240), .ZN(n1259) );
  AND2_X1 U1410 ( .A1(n2010), .A2(n74), .ZN(n1275) );
  INV_X1 U1411 ( .A(n1275), .ZN(n1292) );
  INV_X1 U1476 ( .A(n1275), .ZN(n1293) );
  NAND2_X4 U1543 ( .A1(n1742), .A2(n141), .ZN(n1777) );
  AND2_X1 U1576 ( .A1(n1478), .A2(n74), .ZN(n1344) );
  INV_X1 U1577 ( .A(n1344), .ZN(n1392) );
  INV_X1 U1579 ( .A(n1344), .ZN(n1394) );
  INV_X2 U1591 ( .A(n697), .ZN(n698) );
  NAND2_X2 U1593 ( .A1(n628), .A2(n176), .ZN(n697) );
  INV_X2 U1595 ( .A(n1109), .ZN(n1110) );
  INV_X2 U1621 ( .A(n1075), .ZN(n1076) );
  INV_X2 U1623 ( .A(n317), .ZN(n318) );
  INV_X2 U1625 ( .A(n352), .ZN(n353) );
  INV_X2 U1627 ( .A(n76), .ZN(n77) );
  NOR2_X4 U1629 ( .A1(n2143), .A2(PC_write[1]), .ZN(n141) );
  INV_X2 U1631 ( .A(n663), .ZN(n664) );
  NOR2_X4 U1633 ( .A1(n2142), .A2(n2143), .ZN(n38) );
  INV_X2 U1635 ( .A(n631), .ZN(n630) );
  NAND2_X2 U1637 ( .A1(PC_write[23]), .A2(n3521), .ZN(n1197) );
  NAND2_X2 U1639 ( .A1(PC_write[25]), .A2(n3521), .ZN(n1199) );
  NAND2_X2 U1641 ( .A1(PC_write[27]), .A2(n3521), .ZN(n1201) );
  NAND2_X2 U1642 ( .A1(PC_write[21]), .A2(n3521), .ZN(n1195) );
  NAND2_X2 U1643 ( .A1(PC_write[19]), .A2(n3521), .ZN(n1193) );
  NAND2_X2 U1644 ( .A1(PC_write[29]), .A2(n3521), .ZN(n1203) );
  NAND2_X2 U1645 ( .A1(PC_write[31]), .A2(n3521), .ZN(n1205) );
  NAND2_X2 U1648 ( .A1(PC_write[17]), .A2(n3521), .ZN(n1191) );
  NAND2_X2 U1650 ( .A1(PC_write[15]), .A2(n3521), .ZN(n1189) );
  NAND2_X2 U1652 ( .A1(PC_write[28]), .A2(n3521), .ZN(n1150) );
  NAND2_X2 U1654 ( .A1(PC_write[26]), .A2(n3521), .ZN(n1152) );
  NAND2_X2 U1656 ( .A1(PC_write[13]), .A2(n3521), .ZN(n1187) );
  NAND2_X2 U1658 ( .A1(PC_write[11]), .A2(n3521), .ZN(n1185) );
  NAND2_X2 U1660 ( .A1(PC_write[24]), .A2(n3521), .ZN(n1154) );
  NAND2_X2 U1662 ( .A1(PC_write[22]), .A2(n3521), .ZN(n1156) );
  NAND2_X2 U1664 ( .A1(PC_write[9]), .A2(n3521), .ZN(n1183) );
  NAND2_X2 U1666 ( .A1(PC_write[7]), .A2(n3521), .ZN(n1181) );
  NAND2_X2 U1668 ( .A1(PC_write[20]), .A2(n3521), .ZN(n1158) );
  NAND2_X2 U1670 ( .A1(PC_write[18]), .A2(n3521), .ZN(n1160) );
  NAND2_X2 U1672 ( .A1(PC_write[5]), .A2(n3521), .ZN(n1179) );
  NAND2_X2 U1684 ( .A1(PC_write[6]), .A2(n3521), .ZN(n1172) );
  NAND2_X2 U1686 ( .A1(PC_write[16]), .A2(n3521), .ZN(n1162) );
  NAND2_X2 U1688 ( .A1(PC_write[14]), .A2(n3521), .ZN(n1164) );
  NAND2_X2 U1690 ( .A1(PC_write[8]), .A2(n3521), .ZN(n1170) );
  NAND2_X2 U1692 ( .A1(PC_write[10]), .A2(n3521), .ZN(n1168) );
  NAND2_X2 U1694 ( .A1(PC_write[12]), .A2(n3521), .ZN(n1166) );
  NAND2_X2 U1696 ( .A1(PC_write[30]), .A2(n3521), .ZN(n1147) );
  AND2_X1 U1698 ( .A1(n1478), .A2(n38), .ZN(n1426) );
  INV_X1 U1700 ( .A(n1426), .ZN(n1427) );
  INV_X1 U1702 ( .A(n1426), .ZN(n1428) );
  NOR2_X4 U1706 ( .A1(n2142), .A2(PC_write[0]), .ZN(n74) );
  AND2_X2 U1710 ( .A1(n316), .A2(n177), .ZN(n213) );
  AND2_X1 U1712 ( .A1(n489), .A2(n176), .ZN(n1446) );
  INV_X1 U1714 ( .A(n1446), .ZN(n1463) );
  INV_X1 U1716 ( .A(n1446), .ZN(n1481) );
  INV_X1 U1720 ( .A(n3521), .ZN(n1496) );
  BUF_X8 U1722 ( .A(n3518), .Z(n3521) );
  INV_X2 U1724 ( .A(n906), .ZN(n905) );
  AND2_X1 U1728 ( .A1(n903), .A2(n38), .ZN(n1498) );
  INV_X1 U1730 ( .A(n1498), .ZN(n1611) );
  INV_X1 U1732 ( .A(n1498), .ZN(n1656) );
  INV_X2 U1734 ( .A(n734), .ZN(n733) );
  INV_X2 U1738 ( .A(n248), .ZN(n249) );
  INV_X2 U1749 ( .A(n835), .ZN(n836) );
  NAND2_X2 U1751 ( .A1(n766), .A2(n176), .ZN(n835) );
  AND2_X2 U1755 ( .A1(n731), .A2(n454), .ZN(n903) );
  AND2_X4 U1757 ( .A1(n3437), .A2(n3420), .ZN(n2291) );
  AND2_X4 U1759 ( .A1(n3415), .A2(n3416), .ZN(n2252) );
  AND2_X4 U1761 ( .A1(n3415), .A2(n3420), .ZN(n2257) );
  AND2_X4 U1763 ( .A1(n3421), .A2(n3424), .ZN(n2267) );
  AND2_X4 U1765 ( .A1(n3433), .A2(n3416), .ZN(n2276) );
  NOR3_X2 U1767 ( .A1(n3422), .A2(PC_read[4]), .A3(n3427), .ZN(n3433) );
  AND2_X4 U1769 ( .A1(n3437), .A2(n3416), .ZN(n2286) );
  NOR2_X2 U1771 ( .A1(n3439), .A2(PC_read[2]), .ZN(n3416) );
  NOR3_X2 U1773 ( .A1(PC_read[3]), .A2(PC_read[4]), .A3(n3422), .ZN(n3437) );
  AND2_X4 U1775 ( .A1(n3433), .A2(n3420), .ZN(n2281) );
  AND2_X4 U1776 ( .A1(n3416), .A2(n3424), .ZN(n2262) );
  NAND2_X4 U1777 ( .A1(n3415), .A2(n3421), .ZN(n2254) );
  NAND2_X4 U1794 ( .A1(n3424), .A2(n3420), .ZN(n2264) );
  NOR2_X2 U1810 ( .A1(n3441), .A2(n3439), .ZN(n3420) );
  NAND2_X4 U1811 ( .A1(n3433), .A2(n3418), .ZN(n2273) );
  NAND2_X4 U1827 ( .A1(n3437), .A2(n3418), .ZN(n2283) );
  NAND2_X4 U1828 ( .A1(n3415), .A2(n3418), .ZN(n2249) );
  NAND2_X4 U1844 ( .A1(n3437), .A2(n3421), .ZN(n2288) );
  NAND2_X4 U1845 ( .A1(n3433), .A2(n3421), .ZN(n2278) );
  NAND2_X4 U1848 ( .A1(n3418), .A2(n3424), .ZN(n2259) );
  NAND2_X4 U1850 ( .A1(n3434), .A2(n3418), .ZN(n2272) );
  NOR2_X2 U1852 ( .A1(PC_read[1]), .A2(PC_read[2]), .ZN(n3418) );
  NOR3_X2 U1854 ( .A1(PC_read[0]), .A2(PC_read[4]), .A3(n3427), .ZN(n3434) );
  NAND2_X4 U1856 ( .A1(n3417), .A2(n3421), .ZN(n2253) );
  NAND2_X4 U1858 ( .A1(n3420), .A2(n3425), .ZN(n2263) );
  NAND2_X4 U1860 ( .A1(n3438), .A2(n3418), .ZN(n2282) );
  NOR3_X2 U1862 ( .A1(PC_read[3]), .A2(PC_read[4]), .A3(PC_read[0]), .ZN(n3438) );
  NAND2_X4 U1864 ( .A1(n3418), .A2(n3425), .ZN(n2258) );
  NAND2_X4 U1866 ( .A1(n3434), .A2(n3421), .ZN(n2277) );
  NAND2_X4 U1868 ( .A1(n3438), .A2(n3421), .ZN(n2287) );
  NOR2_X2 U1870 ( .A1(n3441), .A2(PC_read[1]), .ZN(n3421) );
  NAND2_X4 U1872 ( .A1(n3417), .A2(n3418), .ZN(n2248) );
  AND2_X4 U1875 ( .A1(n3421), .A2(n3425), .ZN(n2266) );
  AND2_X4 U1883 ( .A1(n3434), .A2(n3416), .ZN(n2275) );
  AND2_X4 U1885 ( .A1(n3416), .A2(n3425), .ZN(n2261) );
  AND2_X4 U1887 ( .A1(n3434), .A2(n3420), .ZN(n2280) );
  AND2_X4 U1889 ( .A1(n3417), .A2(n3420), .ZN(n2256) );
  AND2_X4 U1891 ( .A1(n3438), .A2(n3420), .ZN(n2290) );
  AND2_X4 U1893 ( .A1(n3438), .A2(n3416), .ZN(n2285) );
  AND2_X4 U1895 ( .A1(n3417), .A2(n3416), .ZN(n2251) );
  NAND2_X4 U1897 ( .A1(n628), .A2(n141), .ZN(n663) );
  AND2_X4 U1901 ( .A1(n766), .A2(n141), .ZN(n3442) );
  INV_X4 U1903 ( .A(n3442), .ZN(n801) );
  NAND2_X4 U1905 ( .A1(n1040), .A2(n141), .ZN(n1075) );
  AND2_X4 U1909 ( .A1(n731), .A2(n592), .ZN(n1040) );
  AND2_X4 U1910 ( .A1(n903), .A2(n176), .ZN(n3443) );
  INV_X4 U1911 ( .A(n3443), .ZN(n972) );
  INV_X2 U1940 ( .A(Set_target[22]), .ZN(n85) );
  INV_X2 U1974 ( .A(Set_target[17]), .ZN(n125) );
  INV_X2 U1975 ( .A(Set_target[16]), .ZN(n91) );
  INV_X2 U1990 ( .A(Set_target[18]), .ZN(n89) );
  NAND2_X4 U1992 ( .A1(n141), .A2(n39), .ZN(n76) );
  AND2_X4 U2009 ( .A1(n177), .A2(n178), .ZN(n39) );
  AND2_X4 U2024 ( .A1(n213), .A2(n176), .ZN(n3444) );
  INV_X4 U2025 ( .A(n3444), .ZN(n282) );
  NAND2_X4 U2026 ( .A1(n351), .A2(n74), .ZN(n352) );
  NAND2_X4 U2042 ( .A1(n351), .A2(n38), .ZN(n317) );
  AND2_X4 U2077 ( .A1(n489), .A2(n141), .ZN(n3445) );
  INV_X4 U2078 ( .A(n3445), .ZN(n524) );
  AND2_X4 U2094 ( .A1(n766), .A2(n74), .ZN(n3446) );
  INV_X4 U2096 ( .A(n3446), .ZN(n769) );
  OR2_X4 U2111 ( .A1(n3447), .A2(n3448), .ZN(n631) );
  INV_X1 U2112 ( .A(n628), .ZN(n3447) );
  INV_X1 U2114 ( .A(n74), .ZN(n3448) );
  MUX2_X1 U2116 ( .A(Set_target[22]), .B(\pc_target[16][22] ), .S(n1463), .Z(
        n5974) );
  INV_X2 U2118 ( .A(n1043), .ZN(n1042) );
  NAND2_X4 U2120 ( .A1(n1040), .A2(n74), .ZN(n1043) );
  INV_X2 U2122 ( .A(Set_target[30]), .ZN(n75) );
  INV_X2 U2158 ( .A(Set_target[11]), .ZN(n119) );
  CLKBUF_X1 U2160 ( .A(SetT_NT), .Z(n3518) );
  INV_X2 U2162 ( .A(Set_target[21]), .ZN(n129) );
  INV_X2 U2164 ( .A(Set_target[25]), .ZN(n133) );
  INV_X2 U2166 ( .A(Set_target[24]), .ZN(n83) );
  INV_X2 U2168 ( .A(Set_target[26]), .ZN(n81) );
  INV_X2 U2170 ( .A(Set_target[29]), .ZN(n137) );
  AND2_X2 U2172 ( .A1(n3519), .A2(n316), .ZN(n766) );
  AND2_X1 U2174 ( .A1(n3520), .A2(n1143), .ZN(n3519) );
  AND2_X1 U2175 ( .A1(n3520), .A2(n1143), .ZN(n731) );
  INV_X2 U2180 ( .A(n422), .ZN(n421) );
  AND4_X1 U2186 ( .A1(WR), .A2(SetT_NT), .A3(Enable), .A4(n1144), .ZN(n593) );
  AND2_X2 U2188 ( .A1(n3519), .A2(n178), .ZN(n628) );
  INV_X4 U2192 ( .A(n1611), .ZN(n870) );
  AND2_X2 U2196 ( .A1(n593), .A2(PC_write[4]), .ZN(n177) );
  INV_X2 U2198 ( .A(Set_target[19]), .ZN(n127) );
  INV_X1 U2200 ( .A(n3518), .ZN(n3529) );
  INV_X2 U2202 ( .A(Set_target[23]), .ZN(n131) );
  INV_X2 U2207 ( .A(Set_target[20]), .ZN(n87) );
  INV_X2 U2208 ( .A(Set_target[28]), .ZN(n79) );
  INV_X2 U2209 ( .A(Set_target[27]), .ZN(n135) );
  INV_X1 U2211 ( .A(n1980), .ZN(n3522) );
  INV_X1 U2213 ( .A(n3522), .ZN(n3523) );
  INV_X2 U2215 ( .A(n3522), .ZN(n3524) );
  INV_X1 U2217 ( .A(n1848), .ZN(n3525) );
  INV_X1 U2219 ( .A(n3525), .ZN(n3526) );
  INV_X2 U2221 ( .A(n3525), .ZN(n3527) );
  INV_X2 U2223 ( .A(n1463), .ZN(n559) );
  INV_X2 U2227 ( .A(n216), .ZN(n215) );
  INV_X2 U2229 ( .A(n457), .ZN(n456) );
  INV_X2 U2233 ( .A(n6), .ZN(n5) );
  INV_X1 U2237 ( .A(SetT_NT), .ZN(n3528) );
  INV_X1 U2238 ( .A(n1578), .ZN(n3530) );
  INV_X1 U2239 ( .A(n3530), .ZN(n3531) );
  INV_X1 U2269 ( .A(n3530), .ZN(n3533) );
  INV_X1 U2274 ( .A(n3530), .ZN(n3532) );
  AND2_X4 U2303 ( .A1(n1206), .A2(n176), .ZN(n3534) );
  INV_X4 U2306 ( .A(n3534), .ZN(n1277) );
  AND2_X4 U2308 ( .A1(n1742), .A2(n74), .ZN(n3535) );
  INV_X4 U2310 ( .A(n3535), .ZN(n1745) );
  AND2_X4 U2312 ( .A1(n1206), .A2(n141), .ZN(n3536) );
  INV_X4 U2314 ( .A(n3536), .ZN(n1242) );
  AND2_X4 U2316 ( .A1(n1742), .A2(n38), .ZN(n3537) );
  INV_X4 U2318 ( .A(n3537), .ZN(n1711) );
  AND2_X4 U2320 ( .A1(n1343), .A2(n74), .ZN(n3538) );
  INV_X2 U2324 ( .A(n2044), .ZN(n2042) );
  INV_X2 U2326 ( .A(n1912), .ZN(n1910) );
  INV_X2 U2328 ( .A(n1811), .ZN(n1809) );
  INV_X2 U2330 ( .A(n1642), .ZN(n1640) );
  INV_X2 U2333 ( .A(n1777), .ZN(n1775) );
  INV_X2 U2334 ( .A(n1412), .ZN(n1410) );
  INV_X2 U2337 ( .A(n1392), .ZN(n1479) );
  INV_X2 U2339 ( .A(n3), .ZN(n2144) );
  INV_X2 U2341 ( .A(n1378), .ZN(n1376) );
  INV_X2 U2343 ( .A(n1427), .ZN(n1444) );
  INV_X2 U2347 ( .A(n1292), .ZN(n2011) );
  INV_X2 U2349 ( .A(n1256), .ZN(n1879) );
  INV_X2 U2351 ( .A(n558), .ZN(n1609) );
  INV_X2 U2353 ( .A(n871), .ZN(n2110) );
  INV_X2 U2357 ( .A(n3523), .ZN(n1978) );
  INV_X2 U2359 ( .A(n3526), .ZN(n1846) );
  INV_X2 U2361 ( .A(n3531), .ZN(n1576) );
  BTB_PC_SIZE32_BTBSIZE5_DW01_cmp6_0 eq_43 ( .A({N188, N189, N190, N191, N192, 
        N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, 
        N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, 
        N217, N218, N219}), .B(PC_read), .TC(1'b0), .EQ(N220) );
  DFFR_X1 \pc_target_reg[16][30]  ( .D(n5970), .CK(Clk), .RN(Reset), .QN(n560)
         );
  DFFR_X1 \pc_target_reg[9][30]  ( .D(n6194), .CK(Clk), .RN(Reset), .QN(n803)
         );
  DFFR_X1 \pc_target_reg[4][30]  ( .D(n6354), .CK(Clk), .RN(Reset), .QN(n974)
         );
  DFFR_X1 \pc_target_reg[17][30]  ( .D(n5938), .CK(Clk), .RN(Reset), .QN(n526)
         );
  DFFR_X1 \pc_target_reg[13][30]  ( .D(n6066), .CK(Clk), .RN(Reset), .QN(n665)
         );
  DFFR_X1 \pc_target_reg[5][30]  ( .D(n6322), .CK(Clk), .RN(Reset), .QN(n940)
         );
  DFFR_X1 \pc_target_reg[0][30]  ( .D(n6482), .CK(Clk), .RN(Reset), .QN(n1111)
         );
  DFFR_X1 \pc_target_reg[1][30]  ( .D(n6450), .CK(Clk), .RN(Reset), .QN(n1077)
         );
  DFFR_X1 \pc_target_reg[23][30]  ( .D(n5746), .CK(Clk), .RN(Reset), .QN(n319)
         );
  DFFR_X1 \pc_target_reg[22][30]  ( .D(n5778), .CK(Clk), .RN(Reset), .QN(n354)
         );
  DFFR_X1 \pc_target_reg[25][30]  ( .D(n5682), .CK(Clk), .RN(Reset), .QN(n250)
         );
  DFFR_X1 \pc_target_reg[28][30]  ( .D(n5586), .CK(Clk), .RN(Reset), .QN(n144)
         );
  DFFR_X1 \pc_target_reg[29][30]  ( .D(n5554), .CK(Clk), .RN(Reset), .QN(n78)
         );
  DFFR_X1 \pc_target_reg[8][30]  ( .D(n6226), .CK(Clk), .RN(Reset), .QN(n837)
         );
  DFFR_X1 \pc_target_reg[12][30]  ( .D(n6098), .CK(Clk), .RN(Reset), .QN(n699)
         );
  DFFR_X1 \pc_target_reg[16][22]  ( .D(n5974), .CK(Clk), .RN(Reset), .Q(
        \pc_target[16][22] ), .QN(n564) );
  DFFR_X1 \pc_lut_reg[31][3]  ( .D(n6531), .CK(Clk), .RN(Reset), .Q(
        \pc_lut[31][3] ) );
  DFFR_X1 \pc_lut_reg[31][2]  ( .D(n6528), .CK(Clk), .RN(Reset), .Q(
        \pc_lut[31][2] ) );
  DFFR_X1 \pc_lut_reg[31][1]  ( .D(n6530), .CK(Clk), .RN(Reset), .Q(
        \pc_lut[31][1] ) );
  DFFR_X1 \pc_lut_reg[31][0]  ( .D(n6529), .CK(Clk), .RN(Reset), .Q(
        \pc_lut[31][0] ) );
  DFFR_X1 \pc_lut_reg[27][3]  ( .D(n6659), .CK(Clk), .RN(Reset), .Q(
        \pc_lut[27][3] ) );
  DFFR_X1 \pc_lut_reg[27][1]  ( .D(n6658), .CK(Clk), .RN(Reset), .Q(
        \pc_lut[27][1] ) );
  DFFR_X1 \pc_lut_reg[27][0]  ( .D(n6657), .CK(Clk), .RN(Reset), .Q(
        \pc_lut[27][0] ) );
  DFFR_X1 \pc_lut_reg[31][4]  ( .D(n6527), .CK(Clk), .RN(Reset), .Q(
        \pc_lut[31][4] ) );
  DFFR_X1 \pc_lut_reg[27][4]  ( .D(n6655), .CK(Clk), .RN(Reset), .Q(
        \pc_lut[27][4] ) );
  DFFR_X1 \pc_target_reg[7][31]  ( .D(n6289), .CK(Clk), .RN(Reset), .Q(
        \pc_target[7][31] ) );
  DFFR_X1 \pc_target_reg[7][23]  ( .D(n6285), .CK(Clk), .RN(Reset), .Q(
        \pc_target[7][23] ) );
  DFFR_X1 \pc_target_reg[7][26]  ( .D(n6260), .CK(Clk), .RN(Reset), .Q(
        \pc_target[7][26] ) );
  DFFR_X1 \pc_target_reg[7][19]  ( .D(n6283), .CK(Clk), .RN(Reset), .Q(
        \pc_target[7][19] ) );
  DFFR_X1 \pc_target_reg[7][14]  ( .D(n6266), .CK(Clk), .RN(Reset), .Q(
        \pc_target[7][14] ) );
  DFFR_X1 \pc_target_reg[7][11]  ( .D(n6279), .CK(Clk), .RN(Reset), .Q(
        \pc_target[7][11] ) );
  DFFR_X1 \pc_target_reg[7][30]  ( .D(n6258), .CK(Clk), .RN(Reset), .Q(
        \pc_target[7][30] ) );
  DFFR_X1 \pc_target_reg[7][29]  ( .D(n6288), .CK(Clk), .RN(Reset), .Q(
        \pc_target[7][29] ) );
  DFFR_X1 \pc_target_reg[7][28]  ( .D(n6259), .CK(Clk), .RN(Reset), .Q(
        \pc_target[7][28] ) );
  DFFR_X1 \pc_target_reg[7][27]  ( .D(n6287), .CK(Clk), .RN(Reset), .Q(
        \pc_target[7][27] ) );
  DFFR_X1 \pc_target_reg[7][25]  ( .D(n6286), .CK(Clk), .RN(Reset), .Q(
        \pc_target[7][25] ) );
  DFFR_X1 \pc_target_reg[7][24]  ( .D(n6261), .CK(Clk), .RN(Reset), .Q(
        \pc_target[7][24] ) );
  DFFR_X1 \pc_target_reg[7][22]  ( .D(n6262), .CK(Clk), .RN(Reset), .Q(
        \pc_target[7][22] ) );
  DFFR_X1 \pc_target_reg[7][21]  ( .D(n6284), .CK(Clk), .RN(Reset), .Q(
        \pc_target[7][21] ) );
  DFFR_X1 \pc_target_reg[7][20]  ( .D(n6263), .CK(Clk), .RN(Reset), .Q(
        \pc_target[7][20] ) );
  DFFR_X1 \pc_target_reg[7][18]  ( .D(n6264), .CK(Clk), .RN(Reset), .Q(
        \pc_target[7][18] ) );
  DFFR_X1 \pc_target_reg[7][17]  ( .D(n6282), .CK(Clk), .RN(Reset), .Q(
        \pc_target[7][17] ) );
  DFFR_X1 \pc_target_reg[7][16]  ( .D(n6265), .CK(Clk), .RN(Reset), .Q(
        \pc_target[7][16] ) );
  DFFR_X1 \pc_target_reg[7][15]  ( .D(n6281), .CK(Clk), .RN(Reset), .Q(
        \pc_target[7][15] ) );
  DFFR_X1 \pc_target_reg[7][13]  ( .D(n6280), .CK(Clk), .RN(Reset), .Q(
        \pc_target[7][13] ) );
  DFFR_X1 \pc_target_reg[7][12]  ( .D(n6267), .CK(Clk), .RN(Reset), .Q(
        \pc_target[7][12] ) );
  DFFR_X1 \pc_target_reg[7][10]  ( .D(n6268), .CK(Clk), .RN(Reset), .Q(
        \pc_target[7][10] ) );
  DFFR_X1 \pc_target_reg[7][9]  ( .D(n6278), .CK(Clk), .RN(Reset), .Q(
        \pc_target[7][9] ) );
  DFFR_X1 \pc_target_reg[7][8]  ( .D(n6269), .CK(Clk), .RN(Reset), .Q(
        \pc_target[7][8] ) );
  DFFR_X1 \pc_target_reg[7][7]  ( .D(n6277), .CK(Clk), .RN(Reset), .Q(
        \pc_target[7][7] ) );
  INV_X2 U807 ( .A(n938), .ZN(n939) );
  NAND2_X4 U1141 ( .A1(n903), .A2(n141), .ZN(n938) );
  INV_X2 U1208 ( .A(n3810), .ZN(n1515) );
  NAND2_X4 U1477 ( .A1(n1040), .A2(n176), .ZN(n1109) );
  NAND2_X4 U1542 ( .A1(n766), .A2(n38), .ZN(n734) );
  OAI211_X1 U1581 ( .C1(n3528), .C2(n1144), .A(Enable), .B(WR), .ZN(n3793) );
  NOR2_X1 U1583 ( .A1(n1708), .A2(PC_write[4]), .ZN(n3794) );
  NAND2_X4 U1585 ( .A1(n903), .A2(n74), .ZN(n906) );
  NAND2_X4 U1587 ( .A1(n213), .A2(n141), .ZN(n248) );
  INV_X2 U1589 ( .A(n3538), .ZN(n1346) );
  INV_X2 U1597 ( .A(n596), .ZN(n595) );
  NAND2_X4 U1704 ( .A1(n628), .A2(n38), .ZN(n596) );
  AND2_X1 U1708 ( .A1(n1206), .A2(n38), .ZN(n3795) );
  INV_X4 U1711 ( .A(n3795), .ZN(n1148) );
  AND4_X1 U1718 ( .A1(WR), .A2(SetT_NT), .A3(Enable), .A4(n1144), .ZN(n3520)
         );
  INV_X2 U1726 ( .A(n3805), .ZN(n1209) );
  AND2_X2 U1736 ( .A1(n1309), .A2(n592), .ZN(n1608) );
  AND2_X1 U1743 ( .A1(n1343), .A2(n38), .ZN(n3796) );
  INV_X4 U1753 ( .A(n3796), .ZN(n1312) );
  INV_X2 U1846 ( .A(n1008), .ZN(n1007) );
  NAND2_X4 U1899 ( .A1(n1040), .A2(n38), .ZN(n1008) );
  INV_X2 U1907 ( .A(n142), .ZN(n143) );
  NAND2_X4 U1913 ( .A1(n176), .A2(n39), .ZN(n142) );
  NAND2_X4 U1915 ( .A1(n213), .A2(n74), .ZN(n216) );
  AND2_X4 U1917 ( .A1(n213), .A2(n38), .ZN(n3797) );
  INV_X4 U1919 ( .A(n3797), .ZN(n181) );
  NAND2_X4 U1921 ( .A1(n489), .A2(n38), .ZN(n457) );
  NAND2_X4 U1923 ( .A1(n38), .A2(n39), .ZN(n6) );
  AND2_X4 U1925 ( .A1(n74), .A2(n39), .ZN(n3798) );
  INV_X4 U1927 ( .A(n3798), .ZN(n42) );
  NAND2_X4 U1929 ( .A1(n351), .A2(n176), .ZN(n422) );
  AND2_X4 U1931 ( .A1(n454), .A2(n177), .ZN(n351) );
  NAND2_X4 U1933 ( .A1(n1343), .A2(n176), .ZN(n1412) );
  AND2_X4 U1935 ( .A1(n351), .A2(n141), .ZN(n3799) );
  INV_X4 U1937 ( .A(n3799), .ZN(n388) );
  INV_X2 U1941 ( .A(n492), .ZN(n491) );
  NAND2_X4 U1947 ( .A1(n489), .A2(n74), .ZN(n492) );
  AND2_X2 U1949 ( .A1(n592), .A2(n177), .ZN(n489) );
  AND2_X4 U1951 ( .A1(n1478), .A2(n176), .ZN(n3800) );
  INV_X4 U1953 ( .A(n3800), .ZN(n1547) );
  AND2_X2 U1955 ( .A1(n1843), .A2(n178), .ZN(n1742) );
  INV_X1 U1957 ( .A(n3796), .ZN(n3801) );
  INV_X1 U1959 ( .A(n3801), .ZN(n3802) );
  INV_X2 U1961 ( .A(n3801), .ZN(n3804) );
  INV_X2 U1963 ( .A(n3801), .ZN(n3803) );
  AND2_X4 U1965 ( .A1(n1206), .A2(n74), .ZN(n3805) );
  INV_X1 U1967 ( .A(n3795), .ZN(n3806) );
  INV_X1 U1969 ( .A(n3806), .ZN(n3807) );
  INV_X2 U1971 ( .A(n3806), .ZN(n3809) );
  INV_X2 U1973 ( .A(n3806), .ZN(n3808) );
  AND2_X4 U2008 ( .A1(n1478), .A2(n141), .ZN(n3810) );
  NAND2_X4 U2043 ( .A1(n1343), .A2(n141), .ZN(n1378) );
  AND2_X2 U2044 ( .A1(n1309), .A2(n316), .ZN(n1343) );
  AND2_X2 U2062 ( .A1(n1309), .A2(n178), .ZN(n1206) );
  CLKBUF_X3 U2124 ( .A(n3821), .Z(n3811) );
  CLKBUF_X3 U2126 ( .A(n3821), .Z(n3812) );
  CLKBUF_X3 U2128 ( .A(n3820), .Z(n3813) );
  CLKBUF_X3 U2130 ( .A(n3820), .Z(n3814) );
  CLKBUF_X3 U2132 ( .A(n3820), .Z(n3815) );
  CLKBUF_X3 U2134 ( .A(n3819), .Z(n3816) );
  CLKBUF_X3 U2136 ( .A(n3819), .Z(n3817) );
  CLKBUF_X3 U2138 ( .A(n3819), .Z(n3818) );
  CLKBUF_X3 U2145 ( .A(Reset), .Z(n3819) );
  CLKBUF_X3 U2146 ( .A(Reset), .Z(n3820) );
  CLKBUF_X3 U2148 ( .A(Reset), .Z(n3821) );
  CLKBUF_X1 U2150 ( .A(n3976), .Z(n3822) );
  CLKBUF_X1 U2152 ( .A(n3975), .Z(n3823) );
  CLKBUF_X1 U2154 ( .A(n3975), .Z(n3824) );
  CLKBUF_X1 U2156 ( .A(n3975), .Z(n3825) );
  CLKBUF_X1 U2176 ( .A(n3975), .Z(n3826) );
  CLKBUF_X1 U2178 ( .A(n3975), .Z(n3827) );
  CLKBUF_X1 U2182 ( .A(n3975), .Z(n3828) );
  CLKBUF_X1 U2184 ( .A(n3974), .Z(n3829) );
  CLKBUF_X1 U2190 ( .A(n3974), .Z(n3830) );
  CLKBUF_X1 U2194 ( .A(n3974), .Z(n3831) );
  CLKBUF_X1 U2225 ( .A(n3974), .Z(n3832) );
  CLKBUF_X1 U2231 ( .A(n3974), .Z(n3833) );
  CLKBUF_X1 U2235 ( .A(n3974), .Z(n3834) );
  CLKBUF_X1 U2242 ( .A(n3973), .Z(n3835) );
  CLKBUF_X1 U2244 ( .A(n3973), .Z(n3836) );
  CLKBUF_X1 U2246 ( .A(n3973), .Z(n3837) );
  CLKBUF_X1 U2248 ( .A(n3973), .Z(n3838) );
  CLKBUF_X1 U2250 ( .A(n3973), .Z(n3839) );
  CLKBUF_X1 U2252 ( .A(n3973), .Z(n3840) );
  CLKBUF_X1 U2254 ( .A(n3972), .Z(n3841) );
  CLKBUF_X1 U2256 ( .A(n3972), .Z(n3842) );
  CLKBUF_X1 U2258 ( .A(n3972), .Z(n3843) );
  CLKBUF_X1 U2260 ( .A(n3972), .Z(n3844) );
  CLKBUF_X1 U2262 ( .A(n3972), .Z(n3845) );
  CLKBUF_X1 U2264 ( .A(n3972), .Z(n3846) );
  CLKBUF_X1 U2266 ( .A(n3971), .Z(n3847) );
  CLKBUF_X1 U2276 ( .A(n3971), .Z(n3848) );
  CLKBUF_X1 U2278 ( .A(n3971), .Z(n3849) );
  CLKBUF_X1 U2280 ( .A(n3971), .Z(n3850) );
  CLKBUF_X1 U2282 ( .A(n3971), .Z(n3851) );
  CLKBUF_X1 U2284 ( .A(n3971), .Z(n3852) );
  CLKBUF_X1 U2286 ( .A(n3970), .Z(n3853) );
  CLKBUF_X1 U2288 ( .A(n3970), .Z(n3854) );
  CLKBUF_X1 U2290 ( .A(n3970), .Z(n3855) );
  CLKBUF_X1 U2292 ( .A(n3970), .Z(n3856) );
  CLKBUF_X1 U2294 ( .A(n3970), .Z(n3857) );
  CLKBUF_X1 U2296 ( .A(n3970), .Z(n3858) );
  CLKBUF_X1 U2298 ( .A(n3969), .Z(n3859) );
  CLKBUF_X1 U2300 ( .A(n3969), .Z(n3860) );
  CLKBUF_X1 U2302 ( .A(n3969), .Z(n3861) );
  CLKBUF_X1 U2322 ( .A(n3969), .Z(n3862) );
  CLKBUF_X1 U2345 ( .A(n3969), .Z(n3863) );
  CLKBUF_X1 U2355 ( .A(n3969), .Z(n3864) );
  CLKBUF_X1 U2363 ( .A(n3968), .Z(n3865) );
  CLKBUF_X1 U2365 ( .A(n3968), .Z(n3866) );
  CLKBUF_X1 U2366 ( .A(n3968), .Z(n3867) );
  CLKBUF_X1 U2367 ( .A(n3968), .Z(n3868) );
  CLKBUF_X1 U2382 ( .A(n3968), .Z(n3869) );
  CLKBUF_X1 U2384 ( .A(n3968), .Z(n3870) );
  CLKBUF_X1 U2385 ( .A(n3967), .Z(n3871) );
  CLKBUF_X1 U2400 ( .A(n3967), .Z(n3872) );
  CLKBUF_X1 U2401 ( .A(n3967), .Z(n3873) );
  CLKBUF_X1 U2416 ( .A(n3967), .Z(n3874) );
  CLKBUF_X1 U2417 ( .A(n3967), .Z(n3875) );
  CLKBUF_X1 U2418 ( .A(n3967), .Z(n3876) );
  CLKBUF_X1 U2419 ( .A(n3966), .Z(n3877) );
  CLKBUF_X1 U2434 ( .A(n3966), .Z(n3878) );
  CLKBUF_X1 U2435 ( .A(n3966), .Z(n3879) );
  CLKBUF_X1 U2436 ( .A(n3966), .Z(n3880) );
  CLKBUF_X1 U2440 ( .A(n3966), .Z(n3881) );
  CLKBUF_X1 U2442 ( .A(n3966), .Z(n3882) );
  CLKBUF_X1 U2444 ( .A(n3965), .Z(n3883) );
  CLKBUF_X1 U2446 ( .A(n3965), .Z(n3884) );
  CLKBUF_X1 U2448 ( .A(n3965), .Z(n3885) );
  CLKBUF_X1 U2450 ( .A(n3965), .Z(n3886) );
  CLKBUF_X1 U2452 ( .A(n3965), .Z(n3887) );
  CLKBUF_X1 U2454 ( .A(n3965), .Z(n3888) );
  CLKBUF_X1 U2456 ( .A(n3964), .Z(n3889) );
  CLKBUF_X1 U2458 ( .A(n3964), .Z(n3890) );
  CLKBUF_X1 U2460 ( .A(n3964), .Z(n3891) );
  CLKBUF_X1 U2462 ( .A(n3964), .Z(n3892) );
  CLKBUF_X1 U2464 ( .A(n3964), .Z(n3893) );
  CLKBUF_X1 U2465 ( .A(n3964), .Z(n3894) );
  CLKBUF_X1 U2475 ( .A(n3963), .Z(n3895) );
  CLKBUF_X1 U2477 ( .A(n3963), .Z(n3896) );
  CLKBUF_X1 U2479 ( .A(n3963), .Z(n3897) );
  CLKBUF_X1 U2481 ( .A(n3963), .Z(n3898) );
  CLKBUF_X1 U2483 ( .A(n3963), .Z(n3899) );
  CLKBUF_X1 U2485 ( .A(n3963), .Z(n3900) );
  CLKBUF_X1 U2487 ( .A(n3962), .Z(n3901) );
  CLKBUF_X1 U2489 ( .A(n3962), .Z(n3902) );
  CLKBUF_X1 U2491 ( .A(n3962), .Z(n3903) );
  CLKBUF_X1 U2493 ( .A(n3962), .Z(n3904) );
  CLKBUF_X1 U2495 ( .A(n3962), .Z(n3905) );
  CLKBUF_X1 U2497 ( .A(n3962), .Z(n3906) );
  CLKBUF_X1 U2499 ( .A(n3961), .Z(n3907) );
  CLKBUF_X1 U2501 ( .A(n3961), .Z(n3908) );
  CLKBUF_X1 U2502 ( .A(n3961), .Z(n3909) );
  CLKBUF_X1 U2503 ( .A(n3961), .Z(n3910) );
  CLKBUF_X1 U2505 ( .A(n3961), .Z(n3911) );
  CLKBUF_X1 U2507 ( .A(n3961), .Z(n3912) );
  CLKBUF_X1 U2509 ( .A(n3960), .Z(n3913) );
  CLKBUF_X1 U2511 ( .A(n3960), .Z(n3914) );
  CLKBUF_X1 U2513 ( .A(n3960), .Z(n3915) );
  CLKBUF_X1 U2515 ( .A(n3960), .Z(n3916) );
  CLKBUF_X1 U2517 ( .A(n3960), .Z(n3917) );
  CLKBUF_X1 U2519 ( .A(n3960), .Z(n3918) );
  CLKBUF_X1 U2521 ( .A(n3959), .Z(n3919) );
  CLKBUF_X1 U2523 ( .A(n3959), .Z(n3920) );
  CLKBUF_X1 U2525 ( .A(n3959), .Z(n3921) );
  CLKBUF_X1 U2527 ( .A(n3959), .Z(n3922) );
  CLKBUF_X1 U2529 ( .A(n3959), .Z(n3923) );
  CLKBUF_X1 U2530 ( .A(n3959), .Z(n3924) );
  CLKBUF_X1 U2533 ( .A(n3958), .Z(n3925) );
  CLKBUF_X1 U2539 ( .A(n3958), .Z(n3926) );
  CLKBUF_X1 U2541 ( .A(n3958), .Z(n3927) );
  CLKBUF_X1 U2543 ( .A(n3958), .Z(n3928) );
  CLKBUF_X1 U2545 ( .A(n3958), .Z(n3929) );
  CLKBUF_X1 U2547 ( .A(n3958), .Z(n3930) );
  CLKBUF_X1 U2549 ( .A(n3957), .Z(n3931) );
  CLKBUF_X1 U2551 ( .A(n3957), .Z(n3932) );
  CLKBUF_X1 U2553 ( .A(n3957), .Z(n3933) );
  CLKBUF_X1 U2555 ( .A(n3957), .Z(n3934) );
  CLKBUF_X1 U2557 ( .A(n3957), .Z(n3935) );
  CLKBUF_X1 U2559 ( .A(n3957), .Z(n3936) );
  CLKBUF_X1 U2561 ( .A(n3956), .Z(n3937) );
  CLKBUF_X1 U2563 ( .A(n3956), .Z(n3938) );
  CLKBUF_X1 U2565 ( .A(n3956), .Z(n3939) );
  CLKBUF_X1 U2566 ( .A(n3956), .Z(n3940) );
  CLKBUF_X1 U2567 ( .A(n3956), .Z(n3941) );
  CLKBUF_X1 U2581 ( .A(n3956), .Z(n3942) );
  CLKBUF_X1 U2584 ( .A(n3955), .Z(n3943) );
  CLKBUF_X1 U2600 ( .A(n3955), .Z(n3944) );
  CLKBUF_X1 U2601 ( .A(n3955), .Z(n3945) );
  CLKBUF_X1 U2615 ( .A(n3955), .Z(n3946) );
  CLKBUF_X1 U2617 ( .A(n3955), .Z(n3947) );
  CLKBUF_X1 U2618 ( .A(n3955), .Z(n3948) );
  CLKBUF_X1 U2634 ( .A(n3954), .Z(n3949) );
  CLKBUF_X1 U2635 ( .A(n3954), .Z(n3950) );
  CLKBUF_X1 U2636 ( .A(n3954), .Z(n3951) );
  CLKBUF_X1 U2639 ( .A(n3954), .Z(n3952) );
  CLKBUF_X1 U2641 ( .A(n3954), .Z(n3953) );
  CLKBUF_X3 U2643 ( .A(n3811), .Z(n3954) );
  CLKBUF_X3 U2645 ( .A(n3811), .Z(n3955) );
  CLKBUF_X3 U2647 ( .A(n3811), .Z(n3956) );
  CLKBUF_X3 U2649 ( .A(n3812), .Z(n3957) );
  CLKBUF_X3 U2651 ( .A(n3812), .Z(n3958) );
  CLKBUF_X3 U2653 ( .A(n3812), .Z(n3959) );
  CLKBUF_X3 U2655 ( .A(n3813), .Z(n3960) );
  CLKBUF_X3 U2657 ( .A(n3813), .Z(n3961) );
  CLKBUF_X3 U2659 ( .A(n3813), .Z(n3962) );
  CLKBUF_X3 U2661 ( .A(n3814), .Z(n3963) );
  CLKBUF_X3 U2663 ( .A(n3814), .Z(n3964) );
  CLKBUF_X3 U2664 ( .A(n3814), .Z(n3965) );
  CLKBUF_X3 U2665 ( .A(n3815), .Z(n3966) );
  CLKBUF_X3 U2673 ( .A(n3815), .Z(n3967) );
  CLKBUF_X3 U2675 ( .A(n3815), .Z(n3968) );
  CLKBUF_X3 U2677 ( .A(n3816), .Z(n3969) );
  CLKBUF_X3 U2679 ( .A(n3816), .Z(n3970) );
  CLKBUF_X3 U2681 ( .A(n3816), .Z(n3971) );
  CLKBUF_X3 U2683 ( .A(n3817), .Z(n3972) );
  CLKBUF_X3 U2685 ( .A(n3817), .Z(n3973) );
  CLKBUF_X3 U2687 ( .A(n3817), .Z(n3974) );
  CLKBUF_X3 U2689 ( .A(n3818), .Z(n3975) );
  CLKBUF_X3 U2691 ( .A(n3818), .Z(n3976) );
endmodule


module datapath_NUMBIT32_ADDRESS_WIDTH_RF5_ADDRESS_WIDTH_DM32 ( CLK, RST, INP1, 
        INP2, IMM26, RS1, RS2, RD, REGF_LATCH_EN, RegA_LATCH_EN, RegB_LATCH_EN, 
        RegIMM_LATCH_EN, RegRD1_LATCH_EN, SIGN_UNSIGN, RFR1_EN, RFR2_EN, 
        MUX_IMM_SEL, JUMP, JUMP_EN, EQ_COND, MUXA_SEL, MUXB_SEL, 
        RALUOUT_LATCH_EN, REGME_LATCH_EN, RegRD2_LATCH_EN, .ALU_OPCODE({
        \ALU_OPCODE[4] , \ALU_OPCODE[3] , \ALU_OPCODE[2] , \ALU_OPCODE[1] , 
        \ALU_OPCODE[0] }), ADDR_DRAM, DATAIN_DRAM, DATAOUT_DRAM, LMD_LATCH_EN, 
        RALUOUT2_LATCH_EN, RegRD3_LATCH_EN, RPCplus8_LATCH_EN, WB_MUX_SEL, 
        RF_WE, ROUT_LATCH_EN, JandL, BRANCH_CTRL_SIG, BRANCH_ALU_OUT, Data_out, 
        REGWRITE_XM, REGWRITE_MW );
  input [31:0] INP1;
  input [15:0] INP2;
  input [25:0] IMM26;
  input [4:0] RS1;
  input [4:0] RS2;
  input [4:0] RD;
  output [31:0] ADDR_DRAM;
  output [31:0] DATAIN_DRAM;
  input [31:0] DATAOUT_DRAM;
  output [31:0] BRANCH_ALU_OUT;
  output [31:0] Data_out;
  input CLK, RST, REGF_LATCH_EN, RegA_LATCH_EN, RegB_LATCH_EN, RegIMM_LATCH_EN,
         RegRD1_LATCH_EN, SIGN_UNSIGN, RFR1_EN, RFR2_EN, MUX_IMM_SEL, JUMP,
         JUMP_EN, EQ_COND, MUXA_SEL, MUXB_SEL, RALUOUT_LATCH_EN,
         REGME_LATCH_EN, RegRD2_LATCH_EN, \ALU_OPCODE[4] , \ALU_OPCODE[3] ,
         \ALU_OPCODE[2] , \ALU_OPCODE[1] , \ALU_OPCODE[0] , LMD_LATCH_EN,
         RALUOUT2_LATCH_EN, RegRD3_LATCH_EN, RPCplus8_LATCH_EN, WB_MUX_SEL,
         RF_WE, ROUT_LATCH_EN, JandL, REGWRITE_XM, REGWRITE_MW;
  output BRANCH_CTRL_SIG;
  wire   n214, n215, n216, BRANCH_T_NT, ForwardC, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n99, n100, n101, n104, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, net92960, net92959,
         net92958, net94217, net94215, net94214, net95253, net95252, net95311,
         net95310, net95343, net95342, net95411, net95416, net95415, net95422,
         net95434, net95433, net95551, net95521, n98, n137, n136, n1, n102,
         n103, n105, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n208, n209, n210, \RPCplus8_OUT[9] , \RPCplus8_OUT[8] ,
         \RPCplus8_OUT[7] , \RPCplus8_OUT[6] , \RPCplus8_OUT[5] ,
         \RPCplus8_OUT[4] , \RPCplus8_OUT[3] , \RPCplus8_OUT[31] ,
         \RPCplus8_OUT[30] , \RPCplus8_OUT[2] , \RPCplus8_OUT[29] ,
         \RPCplus8_OUT[28] , \RPCplus8_OUT[27] , \RPCplus8_OUT[26] ,
         \RPCplus8_OUT[25] , \RPCplus8_OUT[24] , \RPCplus8_OUT[23] ,
         \RPCplus8_OUT[22] , \RPCplus8_OUT[21] , \RPCplus8_OUT[20] ,
         \RPCplus8_OUT[1] , \RPCplus8_OUT[19] , \RPCplus8_OUT[18] ,
         \RPCplus8_OUT[17] , \RPCplus8_OUT[16] , \RPCplus8_OUT[15] ,
         \RPCplus8_OUT[14] , \RPCplus8_OUT[13] , \RPCplus8_OUT[12] ,
         \RPCplus8_OUT[11] , \RPCplus8_OUT[10] , \RPCplus8_OUT[0] ,
         \RME_OUT[9] , \RME_OUT[8] , \RME_OUT[7] , \RME_OUT[6] , \RME_OUT[5] ,
         \RME_OUT[4] , \RME_OUT[3] , \RME_OUT[31] , \RME_OUT[30] ,
         \RME_OUT[2] , \RME_OUT[29] , \RME_OUT[28] , \RME_OUT[27] ,
         \RME_OUT[26] , \RME_OUT[25] , \RME_OUT[24] , \RME_OUT[23] ,
         \RME_OUT[22] , \RME_OUT[21] , \RME_OUT[20] , \RME_OUT[1] ,
         \RME_OUT[19] , \RME_OUT[18] , \RME_OUT[17] , \RME_OUT[16] ,
         \RME_OUT[15] , \RME_OUT[14] , \RME_OUT[13] , \RME_OUT[12] ,
         \RME_OUT[11] , \RME_OUT[10] , \RME_OUT[0] , \RIMM2_OUT[9] ,
         \RIMM2_OUT[8] , \RIMM2_OUT[7] , \RIMM2_OUT[6] , \RIMM2_OUT[5] ,
         \RIMM2_OUT[4] , \RIMM2_OUT[3] , \RIMM2_OUT[31] , \RIMM2_OUT[30] ,
         \RIMM2_OUT[2] , \RIMM2_OUT[29] , \RIMM2_OUT[28] , \RIMM2_OUT[27] ,
         \RIMM2_OUT[26] , \RIMM2_OUT[25] , \RIMM2_OUT[24] , \RIMM2_OUT[23] ,
         \RIMM2_OUT[22] , \RIMM2_OUT[21] , \RIMM2_OUT[20] , \RIMM2_OUT[1] ,
         \RIMM2_OUT[19] , \RIMM2_OUT[18] , \RIMM2_OUT[17] , \RIMM2_OUT[16] ,
         \RIMM2_OUT[15] , \RIMM2_OUT[14] , \RIMM2_OUT[13] , \RIMM2_OUT[12] ,
         \RIMM2_OUT[11] , \RIMM2_OUT[10] , \RIMM2_OUT[0] , \RIMM1_OUT[9] ,
         \RIMM1_OUT[8] , \RIMM1_OUT[7] , \RIMM1_OUT[6] , \RIMM1_OUT[5] ,
         \RIMM1_OUT[4] , \RIMM1_OUT[3] , \RIMM1_OUT[31] , \RIMM1_OUT[30] ,
         \RIMM1_OUT[2] , \RIMM1_OUT[29] , \RIMM1_OUT[28] , \RIMM1_OUT[27] ,
         \RIMM1_OUT[26] , \RIMM1_OUT[25] , \RIMM1_OUT[24] , \RIMM1_OUT[23] ,
         \RIMM1_OUT[22] , \RIMM1_OUT[21] , \RIMM1_OUT[20] , \RIMM1_OUT[1] ,
         \RIMM1_OUT[19] , \RIMM1_OUT[18] , \RIMM1_OUT[17] , \RIMM1_OUT[16] ,
         \RIMM1_OUT[15] , \RIMM1_OUT[14] , \RIMM1_OUT[13] , \RIMM1_OUT[12] ,
         \RIMM1_OUT[11] , \RIMM1_OUT[10] , \RIMM1_OUT[0] , \RD1_OUT[4] ,
         \RD1_OUT[3] , \RD1_OUT[2] , \RD1_OUT[1] , \RD1_OUT[0] ,
         \RALUOUT2_OUT[9] , \RALUOUT2_OUT[8] , \RALUOUT2_OUT[7] ,
         \RALUOUT2_OUT[6] , \RALUOUT2_OUT[5] , \RALUOUT2_OUT[4] ,
         \RALUOUT2_OUT[3] , \RALUOUT2_OUT[31] , \RALUOUT2_OUT[30] ,
         \RALUOUT2_OUT[2] , \RALUOUT2_OUT[29] , \RALUOUT2_OUT[28] ,
         \RALUOUT2_OUT[27] , \RALUOUT2_OUT[26] , \RALUOUT2_OUT[25] ,
         \RALUOUT2_OUT[24] , \RALUOUT2_OUT[23] , \RALUOUT2_OUT[22] ,
         \RALUOUT2_OUT[21] , \RALUOUT2_OUT[20] , \RALUOUT2_OUT[1] ,
         \RALUOUT2_OUT[19] , \RALUOUT2_OUT[18] , \RALUOUT2_OUT[17] ,
         \RALUOUT2_OUT[16] , \RALUOUT2_OUT[15] , \RALUOUT2_OUT[14] ,
         \RALUOUT2_OUT[13] , \RALUOUT2_OUT[12] , \RALUOUT2_OUT[11] ,
         \RALUOUT2_OUT[10] , \RALUOUT2_OUT[0] , \MUX_IMM_OUT[1] ,
         \MUX_IMM_OUT[0] , \LMD_OUT[9] , \LMD_OUT[8] , \LMD_OUT[7] ,
         \LMD_OUT[6] , \LMD_OUT[5] , \LMD_OUT[4] , \LMD_OUT[3] , \LMD_OUT[31] ,
         \LMD_OUT[30] , \LMD_OUT[2] , \LMD_OUT[29] , \LMD_OUT[28] ,
         \LMD_OUT[27] , \LMD_OUT[26] , \LMD_OUT[25] , \LMD_OUT[24] ,
         \LMD_OUT[23] , \LMD_OUT[22] , \LMD_OUT[21] , \LMD_OUT[20] ,
         \LMD_OUT[1] , \LMD_OUT[19] , \LMD_OUT[18] , \LMD_OUT[17] ,
         \LMD_OUT[16] , \LMD_OUT[15] , \LMD_OUT[14] , \LMD_OUT[13] ,
         \LMD_OUT[12] , \LMD_OUT[11] , \LMD_OUT[10] , \LMD_OUT[0] , n217;
  wire   [4:0] MUX_WRaddr_OUT;
  wire   [31:0] MUX_WRdata_OUT;
  wire   [31:0] RA_IN;
  wire   [31:0] RB_IN;
  wire   [31:0] SIGNEXT_IMP2;
  wire   [31:0] SIGNEXT_IMM26;
  wire   [31:0] MUX_IMM_OUT;
  wire   [31:0] RA_OUT;
  wire   [31:0] RB_OUT;
  wire   [31:0] MUX_FORWARDING_BRANCH_OUT;
  wire   [31:0] MUXA_OUT;
  wire   [1:0] ForwardD;
  wire   [31:0] MUXC_OUT;
  wire   [31:0] ALU_inputB;
  wire   [31:0] MUXB_OUT;
  wire   [31:0] ALU_inputA;
  wire   [31:0] ALU_OUT;
  wire   [4:0] RD2_OUT;
  wire   [1:0] ForwardA;
  wire   [1:0] forwardB;
  wire   [4:0] RD3_OUT;

  P4addersub_N32 P4adder_branching ( .A(MUXA_OUT), .B({MUX_IMM_OUT[31], 
        MUX_IMM_OUT[31], MUX_IMM_OUT[31:2]}), .sub_add(1'b0), .Y({
        BRANCH_ALU_OUT[31], n214, BRANCH_ALU_OUT[29:26], n215, 
        BRANCH_ALU_OUT[24], n216, BRANCH_ALU_OUT[22:0]}) );
  alu_NUMBIT32 alu_0 ( .DATA1({ALU_inputA[31], n186, ALU_inputA[29:0]}), 
        .DATA2(MUXB_OUT), .FUNC({\ALU_OPCODE[4] , \ALU_OPCODE[3] , 
        \ALU_OPCODE[2] , \ALU_OPCODE[1] , \ALU_OPCODE[0] }), .OUTALU(ALU_OUT)
         );
  OAI221_X1 U3 ( .B1(net94215), .B2(n3), .C1(net92960), .C2(n5), .A(n6), .ZN(
        MUX_FORWARDING_BRANCH_OUT[9]) );
  NAND2_X1 U4 ( .A1(RA_IN[9]), .A2(n208), .ZN(n6) );
  OAI221_X1 U5 ( .B1(net94215), .B2(n8), .C1(net95433), .C2(n9), .A(n10), .ZN(
        MUX_FORWARDING_BRANCH_OUT[8]) );
  NAND2_X1 U6 ( .A1(RA_IN[8]), .A2(n209), .ZN(n10) );
  OAI221_X1 U7 ( .B1(net95422), .B2(n11), .C1(net95411), .C2(n12), .A(n13), 
        .ZN(MUX_FORWARDING_BRANCH_OUT[7]) );
  NAND2_X1 U8 ( .A1(RA_IN[7]), .A2(n208), .ZN(n13) );
  OAI221_X1 U9 ( .B1(net94217), .B2(n14), .C1(net95433), .C2(n15), .A(n16), 
        .ZN(MUX_FORWARDING_BRANCH_OUT[6]) );
  NAND2_X1 U10 ( .A1(RA_IN[6]), .A2(n208), .ZN(n16) );
  NAND2_X1 U12 ( .A1(RA_IN[5]), .A2(n209), .ZN(n19) );
  OAI221_X1 U13 ( .B1(net95422), .B2(n20), .C1(net95411), .C2(n21), .A(n22), 
        .ZN(MUX_FORWARDING_BRANCH_OUT[4]) );
  NAND2_X1 U14 ( .A1(RA_IN[4]), .A2(n208), .ZN(n22) );
  OAI221_X1 U15 ( .B1(net95422), .B2(n23), .C1(net95411), .C2(n24), .A(n25), 
        .ZN(MUX_FORWARDING_BRANCH_OUT[3]) );
  NAND2_X1 U16 ( .A1(RA_IN[3]), .A2(n208), .ZN(n25) );
  OAI221_X1 U17 ( .B1(net94217), .B2(n26), .C1(net95434), .C2(n27), .A(n28), 
        .ZN(MUX_FORWARDING_BRANCH_OUT[31]) );
  NAND2_X1 U18 ( .A1(RA_IN[31]), .A2(n209), .ZN(n28) );
  OAI221_X1 U19 ( .B1(net95422), .B2(n29), .C1(net95434), .C2(n30), .A(n31), 
        .ZN(MUX_FORWARDING_BRANCH_OUT[30]) );
  NAND2_X1 U20 ( .A1(RA_IN[30]), .A2(n209), .ZN(n31) );
  OAI221_X1 U21 ( .B1(net94215), .B2(n32), .C1(net95434), .C2(n33), .A(n34), 
        .ZN(MUX_FORWARDING_BRANCH_OUT[2]) );
  NAND2_X1 U22 ( .A1(RA_IN[2]), .A2(n209), .ZN(n34) );
  OAI221_X1 U23 ( .B1(net94217), .B2(n35), .C1(net95433), .C2(n36), .A(n37), 
        .ZN(MUX_FORWARDING_BRANCH_OUT[29]) );
  NAND2_X1 U24 ( .A1(RA_IN[29]), .A2(n209), .ZN(n37) );
  OAI221_X1 U25 ( .B1(net94217), .B2(n38), .C1(net92959), .C2(n39), .A(n40), 
        .ZN(MUX_FORWARDING_BRANCH_OUT[28]) );
  NAND2_X1 U26 ( .A1(RA_IN[28]), .A2(n7), .ZN(n40) );
  NAND2_X1 U28 ( .A1(RA_IN[27]), .A2(n208), .ZN(n43) );
  OAI221_X1 U29 ( .B1(net95422), .B2(n44), .C1(net95411), .C2(n45), .A(n46), 
        .ZN(MUX_FORWARDING_BRANCH_OUT[26]) );
  NAND2_X1 U30 ( .A1(RA_IN[26]), .A2(n7), .ZN(n46) );
  OAI221_X1 U31 ( .B1(net95422), .B2(n47), .C1(net95411), .C2(n48), .A(n49), 
        .ZN(MUX_FORWARDING_BRANCH_OUT[25]) );
  NAND2_X1 U32 ( .A1(RA_IN[25]), .A2(n7), .ZN(n49) );
  OAI221_X1 U33 ( .B1(net94215), .B2(n50), .C1(net95411), .C2(n51), .A(n52), 
        .ZN(MUX_FORWARDING_BRANCH_OUT[24]) );
  NAND2_X1 U34 ( .A1(RA_IN[24]), .A2(n7), .ZN(n52) );
  OAI221_X1 U35 ( .B1(net94215), .B2(n53), .C1(net95411), .C2(n54), .A(n55), 
        .ZN(MUX_FORWARDING_BRANCH_OUT[23]) );
  NAND2_X1 U36 ( .A1(RA_IN[23]), .A2(n208), .ZN(n55) );
  OAI221_X1 U37 ( .B1(net94215), .B2(n56), .C1(net95411), .C2(n57), .A(n58), 
        .ZN(MUX_FORWARDING_BRANCH_OUT[22]) );
  NAND2_X1 U38 ( .A1(RA_IN[22]), .A2(n7), .ZN(n58) );
  OAI221_X1 U39 ( .B1(net94217), .B2(n59), .C1(net92960), .C2(n60), .A(n61), 
        .ZN(MUX_FORWARDING_BRANCH_OUT[21]) );
  NAND2_X1 U40 ( .A1(RA_IN[21]), .A2(n7), .ZN(n61) );
  OAI221_X1 U41 ( .B1(net94217), .B2(n62), .C1(net92959), .C2(n63), .A(n64), 
        .ZN(MUX_FORWARDING_BRANCH_OUT[20]) );
  NAND2_X1 U42 ( .A1(RA_IN[20]), .A2(n209), .ZN(n64) );
  NAND2_X1 U44 ( .A1(RA_IN[1]), .A2(n7), .ZN(n67) );
  OAI221_X1 U45 ( .B1(net95422), .B2(n68), .C1(net92960), .C2(n69), .A(n70), 
        .ZN(MUX_FORWARDING_BRANCH_OUT[19]) );
  NAND2_X1 U46 ( .A1(RA_IN[19]), .A2(n208), .ZN(n70) );
  OAI221_X1 U47 ( .B1(net94217), .B2(n71), .C1(net92960), .C2(n72), .A(n73), 
        .ZN(MUX_FORWARDING_BRANCH_OUT[18]) );
  NAND2_X1 U48 ( .A1(RA_IN[18]), .A2(n7), .ZN(n73) );
  OAI221_X1 U49 ( .B1(net94217), .B2(n74), .C1(net92959), .C2(n75), .A(n76), 
        .ZN(MUX_FORWARDING_BRANCH_OUT[17]) );
  NAND2_X1 U50 ( .A1(RA_IN[17]), .A2(n208), .ZN(n76) );
  NAND2_X1 U52 ( .A1(RA_IN[16]), .A2(n7), .ZN(n79) );
  OAI221_X1 U53 ( .B1(net95422), .B2(n80), .C1(net95411), .C2(n81), .A(n82), 
        .ZN(MUX_FORWARDING_BRANCH_OUT[15]) );
  NAND2_X1 U54 ( .A1(RA_IN[15]), .A2(n209), .ZN(n82) );
  OAI221_X1 U55 ( .B1(net94217), .B2(n83), .C1(net95433), .C2(n84), .A(n85), 
        .ZN(MUX_FORWARDING_BRANCH_OUT[14]) );
  NAND2_X1 U56 ( .A1(RA_IN[14]), .A2(n208), .ZN(n85) );
  OAI221_X1 U57 ( .B1(net94217), .B2(n86), .C1(net92959), .C2(n87), .A(n88), 
        .ZN(MUX_FORWARDING_BRANCH_OUT[13]) );
  NAND2_X1 U58 ( .A1(RA_IN[13]), .A2(n7), .ZN(n88) );
  NAND2_X1 U60 ( .A1(RA_IN[12]), .A2(n209), .ZN(n91) );
  OAI221_X1 U61 ( .B1(net95422), .B2(n92), .C1(net95411), .C2(n93), .A(n94), 
        .ZN(MUX_FORWARDING_BRANCH_OUT[11]) );
  NAND2_X1 U62 ( .A1(RA_IN[11]), .A2(n7), .ZN(n94) );
  OAI221_X1 U63 ( .B1(net95422), .B2(n95), .C1(net95434), .C2(n96), .A(n97), 
        .ZN(MUX_FORWARDING_BRANCH_OUT[10]) );
  NAND2_X1 U64 ( .A1(RA_IN[10]), .A2(n209), .ZN(n97) );
  NAND2_X1 U66 ( .A1(RA_IN[0]), .A2(n209), .ZN(n100) );
  NAND2_X1 U68 ( .A1(n210), .A2(n101), .ZN(n4) );
  INV_X1 U70 ( .A(ForwardD[1]), .ZN(n101) );
  OAI221_X1 U71 ( .B1(n3), .B2(net95343), .C1(n5), .C2(net95310), .A(n104), 
        .ZN(ALU_inputB[9]) );
  NAND2_X1 U72 ( .A1(RB_OUT[9]), .A2(n103), .ZN(n104) );
  OAI221_X1 U73 ( .B1(n8), .B2(n185), .C1(n9), .C2(net95310), .A(n106), .ZN(
        ALU_inputB[8]) );
  NAND2_X1 U74 ( .A1(RB_OUT[8]), .A2(n103), .ZN(n106) );
  OAI221_X1 U75 ( .B1(n11), .B2(n184), .C1(n12), .C2(net95310), .A(n107), .ZN(
        ALU_inputB[7]) );
  NAND2_X1 U76 ( .A1(RB_OUT[7]), .A2(n175), .ZN(n107) );
  OAI221_X1 U77 ( .B1(n14), .B2(n184), .C1(n15), .C2(net95310), .A(n108), .ZN(
        ALU_inputB[6]) );
  NAND2_X1 U78 ( .A1(RB_OUT[6]), .A2(n176), .ZN(n108) );
  OAI221_X1 U79 ( .B1(n17), .B2(n184), .C1(n18), .C2(net95310), .A(n109), .ZN(
        ALU_inputB[5]) );
  NAND2_X1 U80 ( .A1(RB_OUT[5]), .A2(n181), .ZN(n109) );
  OAI221_X1 U81 ( .B1(n20), .B2(net95343), .C1(n21), .C2(net95310), .A(n110), 
        .ZN(ALU_inputB[4]) );
  NAND2_X1 U82 ( .A1(RB_OUT[4]), .A2(n181), .ZN(n110) );
  OAI221_X1 U83 ( .B1(n23), .B2(n183), .C1(n24), .C2(net95311), .A(n111), .ZN(
        ALU_inputB[3]) );
  NAND2_X1 U84 ( .A1(RB_OUT[3]), .A2(n102), .ZN(n111) );
  OAI221_X1 U85 ( .B1(n26), .B2(net95343), .C1(n27), .C2(net95310), .A(n112), 
        .ZN(ALU_inputB[31]) );
  NAND2_X1 U86 ( .A1(RB_OUT[31]), .A2(n178), .ZN(n112) );
  OAI221_X1 U87 ( .B1(n29), .B2(n184), .C1(n30), .C2(net95311), .A(n113), .ZN(
        ALU_inputB[30]) );
  NAND2_X1 U88 ( .A1(RB_OUT[30]), .A2(n179), .ZN(n113) );
  OAI221_X1 U89 ( .B1(n32), .B2(net95343), .C1(n33), .C2(net95310), .A(n114), 
        .ZN(ALU_inputB[2]) );
  NAND2_X1 U90 ( .A1(RB_OUT[2]), .A2(n179), .ZN(n114) );
  OAI221_X1 U91 ( .B1(n35), .B2(n185), .C1(n36), .C2(net95311), .A(n115), .ZN(
        ALU_inputB[29]) );
  NAND2_X1 U92 ( .A1(RB_OUT[29]), .A2(n177), .ZN(n115) );
  OAI221_X1 U93 ( .B1(n38), .B2(n184), .C1(n39), .C2(net95311), .A(n116), .ZN(
        ALU_inputB[28]) );
  NAND2_X1 U94 ( .A1(RB_OUT[28]), .A2(n177), .ZN(n116) );
  OAI221_X1 U95 ( .B1(n41), .B2(net95343), .C1(n42), .C2(net95310), .A(n117), 
        .ZN(ALU_inputB[27]) );
  NAND2_X1 U96 ( .A1(RB_OUT[27]), .A2(n105), .ZN(n117) );
  OAI221_X1 U97 ( .B1(n44), .B2(net95343), .C1(n45), .C2(net95310), .A(n118), 
        .ZN(ALU_inputB[26]) );
  NAND2_X1 U98 ( .A1(RB_OUT[26]), .A2(n176), .ZN(n118) );
  OAI221_X1 U99 ( .B1(n47), .B2(n184), .C1(n48), .C2(net95311), .A(n119), .ZN(
        ALU_inputB[25]) );
  NAND2_X1 U100 ( .A1(RB_OUT[25]), .A2(n175), .ZN(n119) );
  OAI221_X1 U101 ( .B1(n50), .B2(n185), .C1(n51), .C2(net95310), .A(n120), 
        .ZN(ALU_inputB[24]) );
  NAND2_X1 U102 ( .A1(RB_OUT[24]), .A2(n177), .ZN(n120) );
  OAI221_X1 U103 ( .B1(n53), .B2(net95343), .C1(n54), .C2(net95311), .A(n121), 
        .ZN(ALU_inputB[23]) );
  NAND2_X1 U104 ( .A1(RB_OUT[23]), .A2(n180), .ZN(n121) );
  OAI221_X1 U105 ( .B1(n56), .B2(n184), .C1(n57), .C2(net95311), .A(n122), 
        .ZN(ALU_inputB[22]) );
  NAND2_X1 U106 ( .A1(RB_OUT[22]), .A2(n180), .ZN(n122) );
  OAI221_X1 U107 ( .B1(n59), .B2(net95343), .C1(n60), .C2(net95310), .A(n123), 
        .ZN(ALU_inputB[21]) );
  NAND2_X1 U108 ( .A1(RB_OUT[21]), .A2(n174), .ZN(n123) );
  OAI221_X1 U109 ( .B1(n62), .B2(n184), .C1(n63), .C2(net95310), .A(n124), 
        .ZN(ALU_inputB[20]) );
  NAND2_X1 U110 ( .A1(RB_OUT[20]), .A2(n103), .ZN(n124) );
  OAI221_X1 U111 ( .B1(n65), .B2(net95343), .C1(n66), .C2(net95311), .A(n125), 
        .ZN(ALU_inputB[1]) );
  NAND2_X1 U112 ( .A1(RB_OUT[1]), .A2(n175), .ZN(n125) );
  OAI221_X1 U113 ( .B1(n68), .B2(net95343), .C1(n69), .C2(net95310), .A(n126), 
        .ZN(ALU_inputB[19]) );
  NAND2_X1 U114 ( .A1(RB_OUT[19]), .A2(n102), .ZN(n126) );
  OAI221_X1 U115 ( .B1(n71), .B2(n185), .C1(n72), .C2(net95310), .A(n127), 
        .ZN(ALU_inputB[18]) );
  NAND2_X1 U116 ( .A1(RB_OUT[18]), .A2(n174), .ZN(n127) );
  OAI221_X1 U117 ( .B1(n74), .B2(n185), .C1(n75), .C2(net95310), .A(n128), 
        .ZN(ALU_inputB[17]) );
  NAND2_X1 U118 ( .A1(RB_OUT[17]), .A2(n105), .ZN(n128) );
  OAI221_X1 U119 ( .B1(n77), .B2(n185), .C1(n78), .C2(net95310), .A(n129), 
        .ZN(ALU_inputB[16]) );
  NAND2_X1 U120 ( .A1(RB_OUT[16]), .A2(n176), .ZN(n129) );
  OAI221_X1 U121 ( .B1(n80), .B2(net95343), .C1(n81), .C2(net95310), .A(n130), 
        .ZN(ALU_inputB[15]) );
  NAND2_X1 U122 ( .A1(RB_OUT[15]), .A2(n102), .ZN(n130) );
  OAI221_X1 U123 ( .B1(n83), .B2(net95343), .C1(n84), .C2(net95310), .A(n131), 
        .ZN(ALU_inputB[14]) );
  NAND2_X1 U124 ( .A1(RB_OUT[14]), .A2(n179), .ZN(n131) );
  OAI221_X1 U125 ( .B1(n86), .B2(net95343), .C1(n87), .C2(net95311), .A(n132), 
        .ZN(ALU_inputB[13]) );
  NAND2_X1 U126 ( .A1(RB_OUT[13]), .A2(n174), .ZN(n132) );
  OAI221_X1 U127 ( .B1(n89), .B2(net95343), .C1(n90), .C2(net95310), .A(n133), 
        .ZN(ALU_inputB[12]) );
  NAND2_X1 U128 ( .A1(RB_OUT[12]), .A2(n105), .ZN(n133) );
  OAI221_X1 U129 ( .B1(n92), .B2(net95343), .C1(n93), .C2(net95310), .A(n134), 
        .ZN(ALU_inputB[11]) );
  NAND2_X1 U130 ( .A1(RB_OUT[11]), .A2(n178), .ZN(n134) );
  OAI221_X1 U131 ( .B1(n95), .B2(n185), .C1(n96), .C2(net95311), .A(n135), 
        .ZN(ALU_inputB[10]) );
  NAND2_X1 U132 ( .A1(RB_OUT[10]), .A2(n178), .ZN(n135) );
  NAND2_X1 U140 ( .A1(RA_OUT[9]), .A2(n141), .ZN(n140) );
  INV_X1 U141 ( .A(MUXC_OUT[9]), .ZN(n5) );
  INV_X1 U142 ( .A(ADDR_DRAM[9]), .ZN(n3) );
  NAND2_X1 U144 ( .A1(RA_OUT[8]), .A2(n141), .ZN(n142) );
  INV_X1 U145 ( .A(MUXC_OUT[8]), .ZN(n9) );
  INV_X1 U146 ( .A(ADDR_DRAM[8]), .ZN(n8) );
  NAND2_X1 U148 ( .A1(RA_OUT[7]), .A2(n141), .ZN(n143) );
  INV_X1 U149 ( .A(MUXC_OUT[7]), .ZN(n12) );
  INV_X1 U150 ( .A(ADDR_DRAM[7]), .ZN(n11) );
  NAND2_X1 U152 ( .A1(RA_OUT[6]), .A2(n141), .ZN(n144) );
  INV_X1 U153 ( .A(MUXC_OUT[6]), .ZN(n15) );
  INV_X1 U154 ( .A(ADDR_DRAM[6]), .ZN(n14) );
  NAND2_X1 U156 ( .A1(RA_OUT[5]), .A2(n141), .ZN(n145) );
  INV_X1 U157 ( .A(MUXC_OUT[5]), .ZN(n18) );
  INV_X1 U158 ( .A(ADDR_DRAM[5]), .ZN(n17) );
  NAND2_X1 U160 ( .A1(RA_OUT[4]), .A2(n141), .ZN(n146) );
  INV_X1 U161 ( .A(MUXC_OUT[4]), .ZN(n21) );
  INV_X1 U162 ( .A(ADDR_DRAM[4]), .ZN(n20) );
  NAND2_X1 U164 ( .A1(RA_OUT[3]), .A2(n141), .ZN(n147) );
  INV_X1 U165 ( .A(MUXC_OUT[3]), .ZN(n24) );
  INV_X1 U166 ( .A(ADDR_DRAM[3]), .ZN(n23) );
  NAND2_X1 U168 ( .A1(RA_OUT[31]), .A2(n141), .ZN(n148) );
  INV_X1 U169 ( .A(MUXC_OUT[31]), .ZN(n27) );
  INV_X1 U170 ( .A(ADDR_DRAM[31]), .ZN(n26) );
  OAI221_X1 U171 ( .B1(n29), .B2(n138), .C1(n30), .C2(n139), .A(n149), .ZN(
        ALU_inputA[30]) );
  NAND2_X1 U172 ( .A1(RA_OUT[30]), .A2(n141), .ZN(n149) );
  INV_X1 U173 ( .A(MUXC_OUT[30]), .ZN(n30) );
  INV_X1 U174 ( .A(ADDR_DRAM[30]), .ZN(n29) );
  NAND2_X1 U176 ( .A1(RA_OUT[2]), .A2(n141), .ZN(n150) );
  INV_X1 U177 ( .A(MUXC_OUT[2]), .ZN(n33) );
  INV_X1 U178 ( .A(ADDR_DRAM[2]), .ZN(n32) );
  NAND2_X1 U180 ( .A1(RA_OUT[29]), .A2(n141), .ZN(n151) );
  INV_X1 U181 ( .A(MUXC_OUT[29]), .ZN(n36) );
  INV_X1 U182 ( .A(ADDR_DRAM[29]), .ZN(n35) );
  OAI221_X1 U183 ( .B1(n38), .B2(n138), .C1(n39), .C2(n139), .A(n152), .ZN(
        ALU_inputA[28]) );
  NAND2_X1 U184 ( .A1(RA_OUT[28]), .A2(n141), .ZN(n152) );
  INV_X1 U185 ( .A(MUXC_OUT[28]), .ZN(n39) );
  INV_X1 U186 ( .A(ADDR_DRAM[28]), .ZN(n38) );
  OAI221_X1 U187 ( .B1(n41), .B2(n138), .C1(n42), .C2(n139), .A(n153), .ZN(
        ALU_inputA[27]) );
  NAND2_X1 U188 ( .A1(RA_OUT[27]), .A2(n141), .ZN(n153) );
  INV_X1 U189 ( .A(MUXC_OUT[27]), .ZN(n42) );
  INV_X1 U190 ( .A(ADDR_DRAM[27]), .ZN(n41) );
  NAND2_X1 U192 ( .A1(RA_OUT[26]), .A2(n141), .ZN(n154) );
  INV_X1 U193 ( .A(MUXC_OUT[26]), .ZN(n45) );
  INV_X1 U194 ( .A(ADDR_DRAM[26]), .ZN(n44) );
  NAND2_X1 U196 ( .A1(RA_OUT[25]), .A2(n141), .ZN(n155) );
  INV_X1 U197 ( .A(MUXC_OUT[25]), .ZN(n48) );
  INV_X1 U198 ( .A(ADDR_DRAM[25]), .ZN(n47) );
  NAND2_X1 U200 ( .A1(RA_OUT[24]), .A2(n141), .ZN(n156) );
  INV_X1 U201 ( .A(MUXC_OUT[24]), .ZN(n51) );
  INV_X1 U202 ( .A(ADDR_DRAM[24]), .ZN(n50) );
  NAND2_X1 U204 ( .A1(RA_OUT[23]), .A2(n141), .ZN(n157) );
  INV_X1 U205 ( .A(MUXC_OUT[23]), .ZN(n54) );
  INV_X1 U206 ( .A(ADDR_DRAM[23]), .ZN(n53) );
  NAND2_X1 U208 ( .A1(RA_OUT[22]), .A2(n141), .ZN(n158) );
  INV_X1 U209 ( .A(MUXC_OUT[22]), .ZN(n57) );
  INV_X1 U210 ( .A(ADDR_DRAM[22]), .ZN(n56) );
  NAND2_X1 U212 ( .A1(RA_OUT[21]), .A2(n141), .ZN(n159) );
  INV_X1 U213 ( .A(MUXC_OUT[21]), .ZN(n60) );
  INV_X1 U214 ( .A(ADDR_DRAM[21]), .ZN(n59) );
  NAND2_X1 U216 ( .A1(RA_OUT[20]), .A2(n141), .ZN(n160) );
  INV_X1 U217 ( .A(MUXC_OUT[20]), .ZN(n63) );
  INV_X1 U218 ( .A(ADDR_DRAM[20]), .ZN(n62) );
  NAND2_X1 U220 ( .A1(RA_OUT[1]), .A2(n141), .ZN(n161) );
  INV_X1 U221 ( .A(MUXC_OUT[1]), .ZN(n66) );
  INV_X1 U222 ( .A(ADDR_DRAM[1]), .ZN(n65) );
  NAND2_X1 U224 ( .A1(RA_OUT[19]), .A2(n141), .ZN(n162) );
  INV_X1 U225 ( .A(MUXC_OUT[19]), .ZN(n69) );
  INV_X1 U226 ( .A(ADDR_DRAM[19]), .ZN(n68) );
  NAND2_X1 U228 ( .A1(RA_OUT[18]), .A2(n141), .ZN(n163) );
  INV_X1 U229 ( .A(MUXC_OUT[18]), .ZN(n72) );
  INV_X1 U230 ( .A(ADDR_DRAM[18]), .ZN(n71) );
  NAND2_X1 U232 ( .A1(RA_OUT[17]), .A2(n141), .ZN(n164) );
  INV_X1 U233 ( .A(MUXC_OUT[17]), .ZN(n75) );
  INV_X1 U234 ( .A(ADDR_DRAM[17]), .ZN(n74) );
  NAND2_X1 U236 ( .A1(RA_OUT[16]), .A2(n141), .ZN(n165) );
  INV_X1 U237 ( .A(MUXC_OUT[16]), .ZN(n78) );
  INV_X1 U238 ( .A(ADDR_DRAM[16]), .ZN(n77) );
  NAND2_X1 U240 ( .A1(RA_OUT[15]), .A2(n141), .ZN(n166) );
  INV_X1 U241 ( .A(MUXC_OUT[15]), .ZN(n81) );
  INV_X1 U242 ( .A(ADDR_DRAM[15]), .ZN(n80) );
  NAND2_X1 U244 ( .A1(RA_OUT[14]), .A2(n141), .ZN(n167) );
  INV_X1 U245 ( .A(MUXC_OUT[14]), .ZN(n84) );
  INV_X1 U246 ( .A(ADDR_DRAM[14]), .ZN(n83) );
  NAND2_X1 U248 ( .A1(RA_OUT[13]), .A2(n141), .ZN(n168) );
  INV_X1 U249 ( .A(MUXC_OUT[13]), .ZN(n87) );
  INV_X1 U250 ( .A(ADDR_DRAM[13]), .ZN(n86) );
  NAND2_X1 U252 ( .A1(RA_OUT[12]), .A2(n141), .ZN(n169) );
  INV_X1 U253 ( .A(MUXC_OUT[12]), .ZN(n90) );
  INV_X1 U254 ( .A(ADDR_DRAM[12]), .ZN(n89) );
  NAND2_X1 U256 ( .A1(RA_OUT[11]), .A2(n141), .ZN(n170) );
  INV_X1 U257 ( .A(MUXC_OUT[11]), .ZN(n93) );
  INV_X1 U258 ( .A(ADDR_DRAM[11]), .ZN(n92) );
  NAND2_X1 U260 ( .A1(RA_OUT[10]), .A2(n141), .ZN(n171) );
  INV_X1 U261 ( .A(MUXC_OUT[10]), .ZN(n96) );
  INV_X1 U262 ( .A(ADDR_DRAM[10]), .ZN(n95) );
  NAND2_X1 U264 ( .A1(RA_OUT[0]), .A2(n141), .ZN(n172) );
  INV_X1 U267 ( .A(MUXC_OUT[0]), .ZN(n99) );
  INV_X1 U269 ( .A(ForwardA[1]), .ZN(n173) );
  OAI221_X1 U65 ( .B1(net94217), .B2(n98), .C1(net95434), .C2(n99), .A(n100), 
        .ZN(MUX_FORWARDING_BRANCH_OUT[0]) );
  INV_X1 U270 ( .A(ADDR_DRAM[0]), .ZN(n98) );
  INV_X1 U138 ( .A(forwardB[1]), .ZN(n137) );
  BUF_X1 U11 ( .A(forwardB[1]), .Z(n1) );
  INV_X1 U27 ( .A(net95415), .ZN(n102) );
  INV_X1 U43 ( .A(net95415), .ZN(n103) );
  INV_X1 U51 ( .A(net95415), .ZN(n105) );
  INV_X1 U59 ( .A(net95415), .ZN(n174) );
  INV_X1 U67 ( .A(net95415), .ZN(n175) );
  INV_X1 U69 ( .A(net95415), .ZN(n176) );
  INV_X1 U133 ( .A(net95415), .ZN(n177) );
  INV_X1 U134 ( .A(net95415), .ZN(n178) );
  BUF_X1 U135 ( .A(net95551), .Z(n179) );
  BUF_X1 U136 ( .A(net95252), .Z(n180) );
  BUF_X1 U137 ( .A(net95253), .Z(n181) );
  INV_X1 U139 ( .A(net95415), .ZN(net95252) );
  INV_X1 U143 ( .A(net95342), .ZN(n182) );
  INV_X1 U147 ( .A(n182), .ZN(n183) );
  INV_X1 U151 ( .A(n182), .ZN(n185) );
  INV_X1 U155 ( .A(n182), .ZN(n184) );
  CLKBUF_X1 U159 ( .A(ALU_inputA[30]), .Z(n186) );
  OAI221_X4 U163 ( .B1(n35), .B2(n138), .C1(n36), .C2(n139), .A(n151), .ZN(
        ALU_inputA[29]) );
  OAI221_X4 U167 ( .B1(n65), .B2(n138), .C1(n66), .C2(n139), .A(n161), .ZN(
        ALU_inputA[1]) );
  OAI221_X4 U175 ( .B1(n17), .B2(n138), .C1(n18), .C2(n139), .A(n145), .ZN(
        ALU_inputA[5]) );
  OAI221_X4 U179 ( .B1(n26), .B2(n138), .C1(n27), .C2(n139), .A(n148), .ZN(
        ALU_inputA[31]) );
  OAI221_X4 U203 ( .B1(n53), .B2(n138), .C1(n54), .C2(n139), .A(n157), .ZN(
        ALU_inputA[23]) );
  OAI221_X4 U207 ( .B1(n71), .B2(n138), .C1(n72), .C2(n139), .A(n163), .ZN(
        ALU_inputA[18]) );
  OAI221_X4 U211 ( .B1(n74), .B2(n138), .C1(n75), .C2(n139), .A(n164), .ZN(
        ALU_inputA[17]) );
  OAI221_X4 U215 ( .B1(n68), .B2(n138), .C1(n69), .C2(n139), .A(n162), .ZN(
        ALU_inputA[19]) );
  OAI221_X4 U219 ( .B1(n62), .B2(n138), .C1(n63), .C2(n139), .A(n160), .ZN(
        ALU_inputA[20]) );
  OAI221_X4 U223 ( .B1(n3), .B2(n138), .C1(n5), .C2(n139), .A(n140), .ZN(
        ALU_inputA[9]) );
  OAI221_X4 U227 ( .B1(n89), .B2(n138), .C1(n90), .C2(n139), .A(n169), .ZN(
        ALU_inputA[12]) );
  OAI221_X4 U231 ( .B1(n8), .B2(n138), .C1(n9), .C2(n139), .A(n142), .ZN(
        ALU_inputA[8]) );
  OAI221_X4 U235 ( .B1(n95), .B2(n138), .C1(n96), .C2(n139), .A(n171), .ZN(
        ALU_inputA[10]) );
  OAI221_X4 U239 ( .B1(n14), .B2(n138), .C1(n15), .C2(n139), .A(n144), .ZN(
        ALU_inputA[6]) );
  OAI221_X4 U243 ( .B1(n83), .B2(n138), .C1(n84), .C2(n139), .A(n167), .ZN(
        ALU_inputA[14]) );
  OAI221_X4 U247 ( .B1(n20), .B2(n138), .C1(n21), .C2(n139), .A(n146), .ZN(
        ALU_inputA[4]) );
  OAI221_X4 U251 ( .B1(n32), .B2(n138), .C1(n33), .C2(n139), .A(n150), .ZN(
        ALU_inputA[2]) );
  OAI221_X4 U255 ( .B1(n59), .B2(n138), .C1(n60), .C2(n139), .A(n159), .ZN(
        ALU_inputA[21]) );
  OAI221_X4 U259 ( .B1(n77), .B2(n138), .C1(n78), .C2(n139), .A(n165), .ZN(
        ALU_inputA[16]) );
  OAI221_X4 U263 ( .B1(n56), .B2(n138), .C1(n57), .C2(n139), .A(n158), .ZN(
        ALU_inputA[22]) );
  OAI221_X4 U265 ( .B1(n11), .B2(n138), .C1(n12), .C2(n139), .A(n143), .ZN(
        ALU_inputA[7]) );
  OAI221_X4 U266 ( .B1(n86), .B2(n138), .C1(n87), .C2(n139), .A(n168), .ZN(
        ALU_inputA[13]) );
  OR2_X2 U268 ( .A1(n1), .A2(forwardB[0]), .ZN(net95415) );
  INV_X1 U271 ( .A(net95521), .ZN(n187) );
  INV_X1 U272 ( .A(n98), .ZN(n188) );
  NAND2_X1 U273 ( .A1(n187), .A2(n191), .ZN(n189) );
  NAND2_X1 U274 ( .A1(n193), .A2(n188), .ZN(n190) );
  AND2_X1 U275 ( .A1(forwardB[0]), .A2(n137), .ZN(n191) );
  NAND2_X1 U276 ( .A1(n192), .A2(n189), .ZN(ALU_inputB[0]) );
  AND2_X1 U277 ( .A1(n190), .A2(n136), .ZN(n192) );
  NOR2_X1 U278 ( .A1(n137), .A2(forwardB[0]), .ZN(n193) );
  OR3_X1 U279 ( .A1(forwardB[0]), .A2(n1), .A3(n194), .ZN(n136) );
  INV_X1 U280 ( .A(RB_OUT[0]), .ZN(n194) );
  INV_X1 U281 ( .A(MUXC_OUT[0]), .ZN(net95521) );
  OR2_X1 U282 ( .A1(n137), .A2(forwardB[0]), .ZN(net95342) );
  OR2_X1 U283 ( .A1(n137), .A2(net95416), .ZN(net95343) );
  OAI221_X4 U284 ( .B1(n98), .B2(n138), .C1(n99), .C2(n139), .A(n172), .ZN(
        ALU_inputA[0]) );
  INV_X2 U285 ( .A(n191), .ZN(net95310) );
  INV_X1 U286 ( .A(n191), .ZN(net95311) );
  CLKBUF_X2 U287 ( .A(n4), .Z(net95411) );
  OAI221_X4 U288 ( .B1(n23), .B2(n138), .C1(n24), .C2(n139), .A(n147), .ZN(
        ALU_inputA[3]) );
  OAI221_X4 U289 ( .B1(net94215), .B2(n17), .C1(net95433), .C2(n18), .A(n19), 
        .ZN(MUX_FORWARDING_BRANCH_OUT[5]) );
  OAI221_X4 U290 ( .B1(n80), .B2(n138), .C1(n81), .C2(n139), .A(n166), .ZN(
        ALU_inputA[15]) );
  CLKBUF_X1 U291 ( .A(MUX_IMM_OUT[16]), .Z(n195) );
  INV_X1 U292 ( .A(net95415), .ZN(net95551) );
  CLKBUF_X1 U293 ( .A(RD2_OUT[4]), .Z(n196) );
  CLKBUF_X1 U294 ( .A(RD2_OUT[2]), .Z(n197) );
  CLKBUF_X1 U295 ( .A(RD2_OUT[1]), .Z(n198) );
  CLKBUF_X1 U296 ( .A(RD2_OUT[0]), .Z(n199) );
  CLKBUF_X1 U297 ( .A(RD3_OUT[4]), .Z(n200) );
  CLKBUF_X1 U298 ( .A(RD3_OUT[3]), .Z(n201) );
  CLKBUF_X1 U299 ( .A(RD3_OUT[0]), .Z(n202) );
  CLKBUF_X1 U300 ( .A(RD2_OUT[3]), .Z(n203) );
  INV_X2 U301 ( .A(net94214), .ZN(net94215) );
  INV_X1 U302 ( .A(net92958), .ZN(net95434) );
  INV_X1 U303 ( .A(net92958), .ZN(net95433) );
  INV_X1 U304 ( .A(net92958), .ZN(net92960) );
  CLKBUF_X3 U305 ( .A(n2), .Z(net95422) );
  CLKBUF_X1 U306 ( .A(MUX_FORWARDING_BRANCH_OUT[10]), .Z(n204) );
  OAI221_X1 U307 ( .B1(net94215), .B2(n89), .C1(net95411), .C2(n90), .A(n91), 
        .ZN(MUX_FORWARDING_BRANCH_OUT[12]) );
  OAI221_X1 U308 ( .B1(net95422), .B2(n41), .C1(net95411), .C2(n42), .A(n43), 
        .ZN(MUX_FORWARDING_BRANCH_OUT[27]) );
  OAI221_X1 U309 ( .B1(net95422), .B2(n65), .C1(net95411), .C2(n66), .A(n67), 
        .ZN(MUX_FORWARDING_BRANCH_OUT[1]) );
  CLKBUF_X1 U310 ( .A(forwardB[0]), .Z(net95416) );
  BUF_X4 U311 ( .A(n214), .Z(BRANCH_ALU_OUT[30]) );
  BUF_X4 U312 ( .A(n215), .Z(BRANCH_ALU_OUT[25]) );
  BUF_X1 U313 ( .A(MUX_FORWARDING_BRANCH_OUT[3]), .Z(n205) );
  OR2_X4 U315 ( .A1(n173), .A2(ForwardA[0]), .ZN(n138) );
  OAI221_X4 U316 ( .B1(n92), .B2(n138), .C1(n93), .C2(n139), .A(n170), .ZN(
        ALU_inputA[11]) );
  NAND2_X4 U317 ( .A1(ForwardA[0]), .A2(n173), .ZN(n139) );
  BUF_X2 U318 ( .A(n216), .Z(BRANCH_ALU_OUT[23]) );
  NOR2_X1 U319 ( .A1(ForwardD[0]), .A2(n217), .ZN(n208) );
  NOR2_X1 U320 ( .A1(ForwardD[0]), .A2(n217), .ZN(n209) );
  NOR2_X1 U321 ( .A1(ForwardD[0]), .A2(ForwardD[1]), .ZN(n7) );
  NOR2_X4 U322 ( .A1(ForwardA[0]), .A2(ForwardA[1]), .ZN(n141) );
  CLKBUF_X1 U323 ( .A(ForwardD[0]), .Z(n210) );
  OR2_X1 U324 ( .A1(n101), .A2(ForwardD[0]), .ZN(n2) );
  INV_X1 U325 ( .A(net95415), .ZN(net95253) );
  INV_X1 U326 ( .A(n2), .ZN(net94214) );
  INV_X2 U327 ( .A(net94214), .ZN(net94217) );
  OAI221_X1 U328 ( .B1(net95422), .B2(n77), .C1(net92960), .C2(n78), .A(n79), 
        .ZN(MUX_FORWARDING_BRANCH_OUT[16]) );
  INV_X1 U329 ( .A(n4), .ZN(net92958) );
  INV_X1 U330 ( .A(net92958), .ZN(net92959) );
  register_file_NUMBIT32_BITADDR5 reg_file_0 ( .CLK(CLK), .RESET(RST), 
        .ENABLE(REGF_LATCH_EN), .RD1(RFR1_EN), .RD2(RFR2_EN), .WR(RF_WE), 
        .ADD_WR(MUX_WRaddr_OUT), .ADD_RD1(RS1), .ADD_RD2(RS2), .DATAIN(
        MUX_WRdata_OUT), .OUT1(RA_IN), .OUT2(RB_IN) );
  signExtend_NUMBIT_in16_NUMBIT_out32 signExtend_0 ( .in_s(INP2), 
        .sign_unsign(SIGN_UNSIGN), .out_s(SIGNEXT_IMP2) );
  signExtend_NUMBIT_in26_NUMBIT_out32 signExtend_1 ( .in_s(IMM26), 
        .sign_unsign(1'b1), .out_s(SIGNEXT_IMM26) );
  MUX21_GENERIC_N32_0 mux_IMM ( .A(SIGNEXT_IMP2), .B(SIGNEXT_IMM26), .SEL(
        MUX_IMM_SEL), .Y({MUX_IMM_OUT[31:2], \MUX_IMM_OUT[1] , 
        \MUX_IMM_OUT[0] }) );
  reg_NUMBIT32_0 reg_in1 ( .clk(CLK), .en(RegIMM_LATCH_EN), .rst(RST), .d(INP1), .q({\RIMM1_OUT[31] , \RIMM1_OUT[30] , \RIMM1_OUT[29] , \RIMM1_OUT[28] , 
        \RIMM1_OUT[27] , \RIMM1_OUT[26] , \RIMM1_OUT[25] , \RIMM1_OUT[24] , 
        \RIMM1_OUT[23] , \RIMM1_OUT[22] , \RIMM1_OUT[21] , \RIMM1_OUT[20] , 
        \RIMM1_OUT[19] , \RIMM1_OUT[18] , \RIMM1_OUT[17] , \RIMM1_OUT[16] , 
        \RIMM1_OUT[15] , \RIMM1_OUT[14] , \RIMM1_OUT[13] , \RIMM1_OUT[12] , 
        \RIMM1_OUT[11] , \RIMM1_OUT[10] , \RIMM1_OUT[9] , \RIMM1_OUT[8] , 
        \RIMM1_OUT[7] , \RIMM1_OUT[6] , \RIMM1_OUT[5] , \RIMM1_OUT[4] , 
        \RIMM1_OUT[3] , \RIMM1_OUT[2] , \RIMM1_OUT[1] , \RIMM1_OUT[0] }) );
  reg_NUMBIT32_9 reg_A ( .clk(CLK), .en(RegA_LATCH_EN), .rst(RST), .d(RA_IN), 
        .q(RA_OUT) );
  reg_NUMBIT32_8 reg_B ( .clk(CLK), .en(RegB_LATCH_EN), .rst(RST), .d(RB_IN), 
        .q(RB_OUT) );
  reg_NUMBIT32_7 reg_in2 ( .clk(CLK), .en(RegIMM_LATCH_EN), .rst(RST), .d({
        MUX_IMM_OUT[31:17], n195, MUX_IMM_OUT[15:2], \MUX_IMM_OUT[1] , 
        \MUX_IMM_OUT[0] }), .q({\RIMM2_OUT[31] , \RIMM2_OUT[30] , 
        \RIMM2_OUT[29] , \RIMM2_OUT[28] , \RIMM2_OUT[27] , \RIMM2_OUT[26] , 
        \RIMM2_OUT[25] , \RIMM2_OUT[24] , \RIMM2_OUT[23] , \RIMM2_OUT[22] , 
        \RIMM2_OUT[21] , \RIMM2_OUT[20] , \RIMM2_OUT[19] , \RIMM2_OUT[18] , 
        \RIMM2_OUT[17] , \RIMM2_OUT[16] , \RIMM2_OUT[15] , \RIMM2_OUT[14] , 
        \RIMM2_OUT[13] , \RIMM2_OUT[12] , \RIMM2_OUT[11] , \RIMM2_OUT[10] , 
        \RIMM2_OUT[9] , \RIMM2_OUT[8] , \RIMM2_OUT[7] , \RIMM2_OUT[6] , 
        \RIMM2_OUT[5] , \RIMM2_OUT[4] , \RIMM2_OUT[3] , \RIMM2_OUT[2] , 
        \RIMM2_OUT[1] , \RIMM2_OUT[0] }) );
  reg_NUMBIT5_0 reg_RD1 ( .clk(CLK), .en(RegRD1_LATCH_EN), .rst(RST), .d(RD), 
        .q({\RD1_OUT[4] , \RD1_OUT[3] , \RD1_OUT[2] , \RD1_OUT[1] , 
        \RD1_OUT[0] }) );
  BranchMgmt_NUMBIT32 BranchMgmt_0 ( .Rin(MUX_FORWARDING_BRANCH_OUT), .Cond(
        EQ_COND), .Jump(JUMP), .Branch(BRANCH_T_NT) );
  MUX21 mux_BRANCH ( .A(BRANCH_T_NT), .B(1'b0), .SEL(JUMP_EN), .Y(
        BRANCH_CTRL_SIG) );
  MUX21_GENERIC_N32_5 mux_A ( .A(INP1), .B({MUX_FORWARDING_BRANCH_OUT[31:11], 
        n204, MUX_FORWARDING_BRANCH_OUT[9:4], n205, 
        MUX_FORWARDING_BRANCH_OUT[2:0]}), .SEL(MUXA_SEL), .Y(MUXA_OUT) );
  MUX21_GENERIC_N32_4 mux_B ( .A(ALU_inputB), .B({\RIMM2_OUT[31] , 
        \RIMM2_OUT[30] , \RIMM2_OUT[29] , \RIMM2_OUT[28] , \RIMM2_OUT[27] , 
        \RIMM2_OUT[26] , \RIMM2_OUT[25] , \RIMM2_OUT[24] , \RIMM2_OUT[23] , 
        \RIMM2_OUT[22] , \RIMM2_OUT[21] , \RIMM2_OUT[20] , \RIMM2_OUT[19] , 
        \RIMM2_OUT[18] , \RIMM2_OUT[17] , \RIMM2_OUT[16] , \RIMM2_OUT[15] , 
        \RIMM2_OUT[14] , \RIMM2_OUT[13] , \RIMM2_OUT[12] , \RIMM2_OUT[11] , 
        \RIMM2_OUT[10] , \RIMM2_OUT[9] , \RIMM2_OUT[8] , \RIMM2_OUT[7] , 
        \RIMM2_OUT[6] , \RIMM2_OUT[5] , \RIMM2_OUT[4] , \RIMM2_OUT[3] , 
        \RIMM2_OUT[2] , \RIMM2_OUT[1] , \RIMM2_OUT[0] }), .SEL(MUXB_SEL), .Y(
        MUXB_OUT) );
  reg_NUMBIT32_6 reg_ALUOUT ( .clk(CLK), .en(RALUOUT_LATCH_EN), .rst(RST), .d(
        ALU_OUT), .q(ADDR_DRAM) );
  reg_NUMBIT32_5 reg_ME ( .clk(CLK), .en(REGME_LATCH_EN), .rst(RST), .d(RB_OUT), .q({\RME_OUT[31] , \RME_OUT[30] , \RME_OUT[29] , \RME_OUT[28] , 
        \RME_OUT[27] , \RME_OUT[26] , \RME_OUT[25] , \RME_OUT[24] , 
        \RME_OUT[23] , \RME_OUT[22] , \RME_OUT[21] , \RME_OUT[20] , 
        \RME_OUT[19] , \RME_OUT[18] , \RME_OUT[17] , \RME_OUT[16] , 
        \RME_OUT[15] , \RME_OUT[14] , \RME_OUT[13] , \RME_OUT[12] , 
        \RME_OUT[11] , \RME_OUT[10] , \RME_OUT[9] , \RME_OUT[8] , \RME_OUT[7] , 
        \RME_OUT[6] , \RME_OUT[5] , \RME_OUT[4] , \RME_OUT[3] , \RME_OUT[2] , 
        \RME_OUT[1] , \RME_OUT[0] }) );
  reg_NUMBIT5_2 reg_RD2 ( .clk(CLK), .en(RegRD2_LATCH_EN), .rst(RST), .d({
        \RD1_OUT[4] , \RD1_OUT[3] , \RD1_OUT[2] , \RD1_OUT[1] , \RD1_OUT[0] }), 
        .q(RD2_OUT) );
  reg_NUMBIT32_4 reg_LMD ( .clk(CLK), .en(LMD_LATCH_EN), .rst(RST), .d(
        DATAOUT_DRAM), .q({\LMD_OUT[31] , \LMD_OUT[30] , \LMD_OUT[29] , 
        \LMD_OUT[28] , \LMD_OUT[27] , \LMD_OUT[26] , \LMD_OUT[25] , 
        \LMD_OUT[24] , \LMD_OUT[23] , \LMD_OUT[22] , \LMD_OUT[21] , 
        \LMD_OUT[20] , \LMD_OUT[19] , \LMD_OUT[18] , \LMD_OUT[17] , 
        \LMD_OUT[16] , \LMD_OUT[15] , \LMD_OUT[14] , \LMD_OUT[13] , 
        \LMD_OUT[12] , \LMD_OUT[11] , \LMD_OUT[10] , \LMD_OUT[9] , 
        \LMD_OUT[8] , \LMD_OUT[7] , \LMD_OUT[6] , \LMD_OUT[5] , \LMD_OUT[4] , 
        \LMD_OUT[3] , \LMD_OUT[2] , \LMD_OUT[1] , \LMD_OUT[0] }) );
  reg_NUMBIT32_3 reg_ALUOUT2 ( .clk(CLK), .en(RALUOUT2_LATCH_EN), .rst(RST), 
        .d(ADDR_DRAM), .q({\RALUOUT2_OUT[31] , \RALUOUT2_OUT[30] , 
        \RALUOUT2_OUT[29] , \RALUOUT2_OUT[28] , \RALUOUT2_OUT[27] , 
        \RALUOUT2_OUT[26] , \RALUOUT2_OUT[25] , \RALUOUT2_OUT[24] , 
        \RALUOUT2_OUT[23] , \RALUOUT2_OUT[22] , \RALUOUT2_OUT[21] , 
        \RALUOUT2_OUT[20] , \RALUOUT2_OUT[19] , \RALUOUT2_OUT[18] , 
        \RALUOUT2_OUT[17] , \RALUOUT2_OUT[16] , \RALUOUT2_OUT[15] , 
        \RALUOUT2_OUT[14] , \RALUOUT2_OUT[13] , \RALUOUT2_OUT[12] , 
        \RALUOUT2_OUT[11] , \RALUOUT2_OUT[10] , \RALUOUT2_OUT[9] , 
        \RALUOUT2_OUT[8] , \RALUOUT2_OUT[7] , \RALUOUT2_OUT[6] , 
        \RALUOUT2_OUT[5] , \RALUOUT2_OUT[4] , \RALUOUT2_OUT[3] , 
        \RALUOUT2_OUT[2] , \RALUOUT2_OUT[1] , \RALUOUT2_OUT[0] }) );
  reg_NUMBIT5_1 reg_RD3 ( .clk(CLK), .en(RegRD3_LATCH_EN), .rst(RST), .d({n196, 
        n203, n197, n198, n199}), .q(RD3_OUT) );
  reg_NUMBIT32_2 PCplus8 ( .clk(CLK), .en(RPCplus8_LATCH_EN), .rst(RST), .d({
        \RIMM1_OUT[31] , \RIMM1_OUT[30] , \RIMM1_OUT[29] , \RIMM1_OUT[28] , 
        \RIMM1_OUT[27] , \RIMM1_OUT[26] , \RIMM1_OUT[25] , \RIMM1_OUT[24] , 
        \RIMM1_OUT[23] , \RIMM1_OUT[22] , \RIMM1_OUT[21] , \RIMM1_OUT[20] , 
        \RIMM1_OUT[19] , \RIMM1_OUT[18] , \RIMM1_OUT[17] , \RIMM1_OUT[16] , 
        \RIMM1_OUT[15] , \RIMM1_OUT[14] , \RIMM1_OUT[13] , \RIMM1_OUT[12] , 
        \RIMM1_OUT[11] , \RIMM1_OUT[10] , \RIMM1_OUT[9] , \RIMM1_OUT[8] , 
        \RIMM1_OUT[7] , \RIMM1_OUT[6] , \RIMM1_OUT[5] , \RIMM1_OUT[4] , 
        \RIMM1_OUT[3] , \RIMM1_OUT[2] , \RIMM1_OUT[1] , \RIMM1_OUT[0] }), .q({
        \RPCplus8_OUT[31] , \RPCplus8_OUT[30] , \RPCplus8_OUT[29] , 
        \RPCplus8_OUT[28] , \RPCplus8_OUT[27] , \RPCplus8_OUT[26] , 
        \RPCplus8_OUT[25] , \RPCplus8_OUT[24] , \RPCplus8_OUT[23] , 
        \RPCplus8_OUT[22] , \RPCplus8_OUT[21] , \RPCplus8_OUT[20] , 
        \RPCplus8_OUT[19] , \RPCplus8_OUT[18] , \RPCplus8_OUT[17] , 
        \RPCplus8_OUT[16] , \RPCplus8_OUT[15] , \RPCplus8_OUT[14] , 
        \RPCplus8_OUT[13] , \RPCplus8_OUT[12] , \RPCplus8_OUT[11] , 
        \RPCplus8_OUT[10] , \RPCplus8_OUT[9] , \RPCplus8_OUT[8] , 
        \RPCplus8_OUT[7] , \RPCplus8_OUT[6] , \RPCplus8_OUT[5] , 
        \RPCplus8_OUT[4] , \RPCplus8_OUT[3] , \RPCplus8_OUT[2] , 
        \RPCplus8_OUT[1] , \RPCplus8_OUT[0] }) );
  MUX21_GENERIC_N32_3 MUX_FORWARD_MEM ( .A(MUXC_OUT), .B({\RME_OUT[31] , 
        \RME_OUT[30] , \RME_OUT[29] , \RME_OUT[28] , \RME_OUT[27] , 
        \RME_OUT[26] , \RME_OUT[25] , \RME_OUT[24] , \RME_OUT[23] , 
        \RME_OUT[22] , \RME_OUT[21] , \RME_OUT[20] , \RME_OUT[19] , 
        \RME_OUT[18] , \RME_OUT[17] , \RME_OUT[16] , \RME_OUT[15] , 
        \RME_OUT[14] , \RME_OUT[13] , \RME_OUT[12] , \RME_OUT[11] , 
        \RME_OUT[10] , \RME_OUT[9] , \RME_OUT[8] , \RME_OUT[7] , \RME_OUT[6] , 
        \RME_OUT[5] , \RME_OUT[4] , \RME_OUT[3] , \RME_OUT[2] , \RME_OUT[1] , 
        \RME_OUT[0] }), .SEL(ForwardC), .Y(DATAIN_DRAM) );
  MUX21_GENERIC_N32_2 mux_C ( .A({\LMD_OUT[31] , \LMD_OUT[30] , \LMD_OUT[29] , 
        \LMD_OUT[28] , \LMD_OUT[27] , \LMD_OUT[26] , \LMD_OUT[25] , 
        \LMD_OUT[24] , \LMD_OUT[23] , \LMD_OUT[22] , \LMD_OUT[21] , 
        \LMD_OUT[20] , \LMD_OUT[19] , \LMD_OUT[18] , \LMD_OUT[17] , 
        \LMD_OUT[16] , \LMD_OUT[15] , \LMD_OUT[14] , \LMD_OUT[13] , 
        \LMD_OUT[12] , \LMD_OUT[11] , \LMD_OUT[10] , \LMD_OUT[9] , 
        \LMD_OUT[8] , \LMD_OUT[7] , \LMD_OUT[6] , \LMD_OUT[5] , \LMD_OUT[4] , 
        \LMD_OUT[3] , \LMD_OUT[2] , \LMD_OUT[1] , \LMD_OUT[0] }), .B({
        \RALUOUT2_OUT[31] , \RALUOUT2_OUT[30] , \RALUOUT2_OUT[29] , 
        \RALUOUT2_OUT[28] , \RALUOUT2_OUT[27] , \RALUOUT2_OUT[26] , 
        \RALUOUT2_OUT[25] , \RALUOUT2_OUT[24] , \RALUOUT2_OUT[23] , 
        \RALUOUT2_OUT[22] , \RALUOUT2_OUT[21] , \RALUOUT2_OUT[20] , 
        \RALUOUT2_OUT[19] , \RALUOUT2_OUT[18] , \RALUOUT2_OUT[17] , 
        \RALUOUT2_OUT[16] , \RALUOUT2_OUT[15] , \RALUOUT2_OUT[14] , 
        \RALUOUT2_OUT[13] , \RALUOUT2_OUT[12] , \RALUOUT2_OUT[11] , 
        \RALUOUT2_OUT[10] , \RALUOUT2_OUT[9] , \RALUOUT2_OUT[8] , 
        \RALUOUT2_OUT[7] , \RALUOUT2_OUT[6] , \RALUOUT2_OUT[5] , 
        \RALUOUT2_OUT[4] , \RALUOUT2_OUT[3] , \RALUOUT2_OUT[2] , 
        \RALUOUT2_OUT[1] , \RALUOUT2_OUT[0] }), .SEL(WB_MUX_SEL), .Y(MUXC_OUT)
         );
  reg_NUMBIT32_1 reg_OUT ( .clk(CLK), .en(ROUT_LATCH_EN), .rst(RST), .d(
        MUXC_OUT), .q(Data_out) );
  MUX21_GENERIC_N5 mux_WRaddr ( .A({1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .B({n200, 
        n201, RD3_OUT[2:1], n202}), .SEL(JandL), .Y(MUX_WRaddr_OUT) );
  MUX21_GENERIC_N32_1 mux_WRdata ( .A({\RPCplus8_OUT[31] , \RPCplus8_OUT[30] , 
        \RPCplus8_OUT[29] , \RPCplus8_OUT[28] , \RPCplus8_OUT[27] , 
        \RPCplus8_OUT[26] , \RPCplus8_OUT[25] , \RPCplus8_OUT[24] , 
        \RPCplus8_OUT[23] , \RPCplus8_OUT[22] , \RPCplus8_OUT[21] , 
        \RPCplus8_OUT[20] , \RPCplus8_OUT[19] , \RPCplus8_OUT[18] , 
        \RPCplus8_OUT[17] , \RPCplus8_OUT[16] , \RPCplus8_OUT[15] , 
        \RPCplus8_OUT[14] , \RPCplus8_OUT[13] , \RPCplus8_OUT[12] , 
        \RPCplus8_OUT[11] , \RPCplus8_OUT[10] , \RPCplus8_OUT[9] , 
        \RPCplus8_OUT[8] , \RPCplus8_OUT[7] , \RPCplus8_OUT[6] , 
        \RPCplus8_OUT[5] , \RPCplus8_OUT[4] , \RPCplus8_OUT[3] , 
        \RPCplus8_OUT[2] , \RPCplus8_OUT[1] , \RPCplus8_OUT[0] }), .B(MUXC_OUT), .SEL(JandL), .Y(MUX_WRdata_OUT) );
  ForwardingUnit_NUMBIT32_ADDRESS_WIDTH_RF5 FORWARDING_UNIT_0 ( .CLK(CLK), 
        .RST(RST), .RS1(RS1), .RS2(RS2), .RD_XM(RD2_OUT), .RD_MW(RD3_OUT), 
        .REGWRITE_XM(REGWRITE_XM), .REGWRITE_MW(REGWRITE_MW), .ForwardA(
        ForwardA), .forwardB(forwardB), .ForwardC(ForwardC), .ForwardD(
        ForwardD) );
  OAI221_X2 U191 ( .B1(n50), .B2(n138), .C1(n51), .C2(n139), .A(n156), .ZN(
        ALU_inputA[24]) );
  OAI221_X2 U195 ( .B1(n47), .B2(n138), .C1(n48), .C2(n139), .A(n155), .ZN(
        ALU_inputA[25]) );
  OAI221_X2 U199 ( .B1(n44), .B2(n138), .C1(n45), .C2(n139), .A(n154), .ZN(
        ALU_inputA[26]) );
  INV_X1 U314 ( .A(n101), .ZN(n217) );
endmodule


module dlx_cu_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE29 ( Clk, Rst, 
        Flush_BTB, STALL, IR_IN, IR_LATCH_EN, NPC_LATCH_EN, I_R_type, 
        REGF_LATCH_EN, RegA_LATCH_EN, RegB_LATCH_EN, RegIMM_LATCH_EN, 
        RegRD1_LATCH_EN, SIGN_UNSIGN, RFR1_EN, RFR2_EN, MUX_IMM_SEL, JUMP, 
        JUMP_EN, EQ_COND, MUXA_SEL, MUXB_SEL, ALU_OUTREG_EN, REGME_LATCH_EN, 
        RegRD2_LATCH_EN, .ALU_OPCODE({\ALU_OPCODE[4] , \ALU_OPCODE[3] , 
        \ALU_OPCODE[2] , \ALU_OPCODE[1] , \ALU_OPCODE[0] }), DRAM_EN, DRAM_RE, 
        DRAM_WE, LMD_LATCH_EN, RALUOUT2_LATCH_EN, RegRD3_LATCH_EN, PC_LATCH_EN, 
        RPCplus8_LATCH_EN, WB_MUX_SEL, RF_WE, ROUT_LATCH_EN, JandL, 
        REGWRITE_DX, REGWRITE_XM, REGWRITE_MW, MEMREAD_DX );
  input [31:0] IR_IN;
  input Clk, Rst, Flush_BTB, STALL;
  output IR_LATCH_EN, NPC_LATCH_EN, I_R_type, REGF_LATCH_EN, RegA_LATCH_EN,
         RegB_LATCH_EN, RegIMM_LATCH_EN, RegRD1_LATCH_EN, SIGN_UNSIGN, RFR1_EN,
         RFR2_EN, MUX_IMM_SEL, JUMP, JUMP_EN, EQ_COND, MUXA_SEL, MUXB_SEL,
         ALU_OUTREG_EN, REGME_LATCH_EN, RegRD2_LATCH_EN, \ALU_OPCODE[4] ,
         \ALU_OPCODE[3] , \ALU_OPCODE[2] , \ALU_OPCODE[1] , \ALU_OPCODE[0] ,
         DRAM_EN, DRAM_RE, DRAM_WE, LMD_LATCH_EN, RALUOUT2_LATCH_EN,
         RegRD3_LATCH_EN, PC_LATCH_EN, RPCplus8_LATCH_EN, WB_MUX_SEL, RF_WE,
         ROUT_LATCH_EN, JandL, REGWRITE_DX, REGWRITE_XM, REGWRITE_MW,
         MEMREAD_DX;
  wire   IR_IN_31, IR_IN_30, IR_IN_29, IR_IN_28, IR_IN_27, IR_IN_26,
         NPC_LATCH_EN, n205, RFR2_EN, n206, REGWRITE_MW, cw_3, cw_2, cw_0,
         cw3_11, cw3_10, cw3_3, cw3_0, cw4_3, \cw4[0] , n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n150, n151,
         n152, n153, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n178, n179, n180, n1, n2, n130, n149, n154, n167, n177, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n238, n239;
  wire   [15:5] cw;
  wire   [8:5] cw3;
  wire   [4:0] aluOpcode_i;
  assign IR_IN_31 = IR_IN[31];
  assign IR_IN_30 = IR_IN[30];
  assign IR_IN_29 = IR_IN[29];
  assign IR_IN_28 = IR_IN[28];
  assign IR_IN_27 = IR_IN[27];
  assign IR_IN_26 = IR_IN[26];
  assign IR_LATCH_EN = NPC_LATCH_EN;
  assign RegB_LATCH_EN = RFR2_EN;
  assign RF_WE = REGWRITE_MW;
  assign ROUT_LATCH_EN = 1'b0;
  assign RegRD1_LATCH_EN = cw[5];

  DFFS_X1 \aluOpcode3_reg[4]  ( .D(aluOpcode_i[4]), .CK(Clk), .SN(n238), .Q(
        ALU_OPCODE[4]) );
  DFFS_X1 \aluOpcode3_reg[1]  ( .D(aluOpcode_i[1]), .CK(Clk), .SN(n238), .Q(
        ALU_OPCODE[1]) );
  AND2_X1 U4 ( .A1(n34), .A2(n35), .ZN(cw_2) );
  NOR2_X1 U5 ( .A1(n36), .A2(n192), .ZN(cw[6]) );
  NOR2_X1 U6 ( .A1(n38), .A2(n192), .ZN(cw[13]) );
  OR2_X1 U7 ( .A1(cw_3), .A2(cw[8]), .ZN(cw[14]) );
  NOR2_X1 U8 ( .A1(n192), .A2(n39), .ZN(cw_3) );
  OAI211_X1 U9 ( .C1(n185), .C2(n40), .A(n41), .B(n42), .ZN(aluOpcode_i[4]) );
  OAI21_X1 U10 ( .B1(n43), .B2(n44), .A(n183), .ZN(n41) );
  NAND4_X1 U11 ( .A1(n46), .A2(n47), .A3(n48), .A4(n49), .ZN(aluOpcode_i[3])
         );
  OAI211_X1 U12 ( .C1(n50), .C2(n181), .A(n154), .B(IR_IN_29), .ZN(n48) );
  AND2_X1 U13 ( .A1(n194), .A2(n53), .ZN(n50) );
  OAI21_X1 U14 ( .B1(n54), .B2(n55), .A(n56), .ZN(n47) );
  INV_X1 U15 ( .A(n57), .ZN(n55) );
  NOR4_X1 U16 ( .A1(IR_IN[4]), .A2(IR_IN[2]), .A3(n58), .A4(n59), .ZN(n54) );
  INV_X1 U17 ( .A(n60), .ZN(n46) );
  NAND4_X1 U18 ( .A1(n61), .A2(n62), .A3(n63), .A4(n64), .ZN(aluOpcode_i[2])
         );
  AOI21_X1 U19 ( .B1(n56), .B2(n65), .A(n60), .ZN(n64) );
  OAI211_X1 U20 ( .C1(n66), .C2(n67), .A(n68), .B(n69), .ZN(n60) );
  NAND3_X1 U21 ( .A1(n70), .A2(n71), .A3(n57), .ZN(n65) );
  AOI22_X1 U22 ( .A1(IR_IN[5]), .A2(n72), .B1(IR_IN[2]), .B2(n73), .ZN(n57) );
  NAND4_X1 U23 ( .A1(n74), .A2(IR_IN[2]), .A3(n75), .A4(n76), .ZN(n70) );
  OAI211_X1 U24 ( .C1(n77), .C2(n181), .A(IR_IN_28), .B(n78), .ZN(n63) );
  NOR2_X1 U25 ( .A1(IR_IN_31), .A2(IR_IN_29), .ZN(n77) );
  NAND4_X1 U26 ( .A1(n42), .A2(n79), .A3(n80), .A4(n81), .ZN(aluOpcode_i[1])
         );
  NOR3_X1 U28 ( .A1(n86), .A2(n154), .A3(n194), .ZN(n85) );
  NOR2_X1 U29 ( .A1(IR_IN_28), .A2(n181), .ZN(n82) );
  OAI21_X1 U30 ( .B1(n44), .B2(n87), .A(n183), .ZN(n79) );
  NAND2_X1 U31 ( .A1(n88), .A2(n89), .ZN(n87) );
  OAI211_X1 U32 ( .C1(n90), .C2(n91), .A(IR_IN[2]), .B(n74), .ZN(n88) );
  NOR2_X1 U33 ( .A1(IR_IN[5]), .A2(n92), .ZN(n90) );
  OAI211_X1 U34 ( .C1(IR_IN[5]), .C2(n93), .A(n94), .B(n95), .ZN(n44) );
  AOI211_X1 U35 ( .C1(n96), .C2(IR_IN[2]), .A(n97), .B(n98), .ZN(n95) );
  NOR3_X1 U36 ( .A1(n99), .A2(IR_IN[2]), .A3(IR_IN[1]), .ZN(n97) );
  NOR2_X1 U37 ( .A1(n100), .A2(n92), .ZN(n96) );
  AOI21_X1 U38 ( .B1(IR_IN[5]), .B2(IR_IN[0]), .A(IR_IN[3]), .ZN(n100) );
  AOI211_X1 U39 ( .C1(IR_IN[0]), .C2(n92), .A(n101), .B(IR_IN[3]), .ZN(n93) );
  INV_X1 U40 ( .A(n102), .ZN(n42) );
  OAI222_X1 U41 ( .A1(n154), .A2(n103), .B1(n190), .B2(n105), .C1(n106), .C2(
        n40), .ZN(n102) );
  AOI21_X1 U43 ( .B1(n154), .B2(IR_IN_28), .A(IR_IN_27), .ZN(n110) );
  AOI22_X1 U44 ( .A1(n111), .A2(n2), .B1(n112), .B2(n185), .ZN(n105) );
  NAND2_X1 U45 ( .A1(n113), .A2(IR_IN_28), .ZN(n111) );
  AOI21_X1 U46 ( .B1(n114), .B2(n2), .A(n115), .ZN(n103) );
  NOR3_X1 U47 ( .A1(n184), .A2(n194), .A3(n53), .ZN(n115) );
  NOR2_X1 U48 ( .A1(IR_IN_31), .A2(IR_IN_26), .ZN(n53) );
  NAND3_X1 U49 ( .A1(n117), .A2(n113), .A3(n194), .ZN(n114) );
  INV_X1 U50 ( .A(n118), .ZN(n113) );
  OAI211_X1 U51 ( .C1(n119), .C2(n2), .A(n80), .B(n120), .ZN(aluOpcode_i[0])
         );
  AOI21_X1 U52 ( .B1(n56), .B2(n121), .A(n122), .ZN(n120) );
  NAND4_X1 U53 ( .A1(n71), .A2(n123), .A3(n124), .A4(n125), .ZN(n121) );
  AOI22_X1 U54 ( .A1(IR_IN[2]), .A2(n126), .B1(n73), .B2(IR_IN[0]), .ZN(n125)
         );
  NOR3_X1 U55 ( .A1(n59), .A2(IR_IN[4]), .A3(n75), .ZN(n73) );
  OAI33_X1 U56 ( .A1(n75), .A2(n98), .A3(n76), .B1(n127), .B2(IR_IN[0]), .B3(
        n128), .ZN(n126) );
  NAND2_X1 U57 ( .A1(n92), .A2(n58), .ZN(n127) );
  INV_X1 U58 ( .A(IR_IN[1]), .ZN(n92) );
  NOR2_X1 U59 ( .A1(n99), .A2(IR_IN[3]), .ZN(n98) );
  INV_X1 U60 ( .A(n91), .ZN(n75) );
  NOR2_X1 U61 ( .A1(n58), .A2(IR_IN[1]), .ZN(n91) );
  NAND4_X1 U62 ( .A1(n74), .A2(IR_IN[1]), .A3(IR_IN[5]), .A4(n101), .ZN(n124)
         );
  OR3_X1 U63 ( .A1(n58), .A2(n76), .A3(n89), .ZN(n123) );
  NAND4_X1 U64 ( .A1(n129), .A2(IR_IN[2]), .A3(IR_IN[1]), .A4(n58), .ZN(n71)
         );
  INV_X1 U65 ( .A(IR_IN[5]), .ZN(n58) );
  AND2_X1 U66 ( .A1(n94), .A2(n183), .ZN(n56) );
  AND3_X1 U67 ( .A1(n62), .A2(n49), .A3(n69), .ZN(n80) );
  AOI221_X1 U68 ( .B1(n167), .B2(n189), .C1(n118), .C2(n131), .A(n132), .ZN(
        n119) );
  NOR3_X1 U69 ( .A1(n194), .A2(n185), .A3(n66), .ZN(n132) );
  NOR2_X1 U70 ( .A1(n133), .A2(n109), .ZN(n118) );
  AOI21_X1 U71 ( .B1(n134), .B2(n135), .A(n187), .ZN(SIGN_UNSIGN) );
  INV_X1 U73 ( .A(n139), .ZN(n138) );
  OAI22_X1 U74 ( .A1(n140), .A2(n141), .B1(IR_IN_26), .B2(n86), .ZN(n137) );
  NAND3_X1 U75 ( .A1(IR_IN[5]), .A2(n142), .A3(n94), .ZN(n136) );
  NOR3_X1 U76 ( .A1(IR_IN[6]), .A2(IR_IN[10]), .A3(n143), .ZN(n94) );
  OR3_X1 U77 ( .A1(IR_IN[9]), .A2(IR_IN[8]), .A3(IR_IN[7]), .ZN(n143) );
  INV_X1 U78 ( .A(n144), .ZN(n142) );
  AOI211_X1 U79 ( .C1(n101), .C2(n129), .A(n72), .B(n43), .ZN(n144) );
  NOR4_X1 U80 ( .A1(n59), .A2(n101), .A3(n99), .A4(IR_IN[1]), .ZN(n43) );
  INV_X1 U81 ( .A(IR_IN[3]), .ZN(n59) );
  NOR2_X1 U82 ( .A1(n89), .A2(n99), .ZN(n72) );
  INV_X1 U83 ( .A(IR_IN[4]), .ZN(n99) );
  NAND3_X1 U84 ( .A1(IR_IN[1]), .A2(n101), .A3(IR_IN[3]), .ZN(n89) );
  NOR2_X1 U85 ( .A1(n128), .A2(n76), .ZN(n129) );
  INV_X1 U86 ( .A(IR_IN[0]), .ZN(n76) );
  INV_X1 U87 ( .A(n74), .ZN(n128) );
  NOR2_X1 U88 ( .A1(IR_IN[3]), .A2(IR_IN[4]), .ZN(n74) );
  INV_X1 U89 ( .A(IR_IN[2]), .ZN(n101) );
  NOR3_X1 U90 ( .A1(n145), .A2(n146), .A3(n196), .ZN(n134) );
  AOI21_X1 U91 ( .B1(n39), .B2(n36), .A(n192), .ZN(cw[5]) );
  AND2_X1 U92 ( .A1(n148), .A2(n177), .ZN(n36) );
  NOR2_X1 U93 ( .A1(n150), .A2(n192), .ZN(RegIMM_LATCH_EN) );
  OR2_X1 U94 ( .A1(cw[8]), .A2(cw[15]), .ZN(RFR2_EN) );
  AND2_X1 U95 ( .A1(n183), .A2(n35), .ZN(cw[15]) );
  NOR2_X1 U96 ( .A1(n139), .A2(n192), .ZN(cw[8]) );
  OR2_X1 U97 ( .A1(n151), .A2(n239), .ZN(n206) );
  AOI21_X1 U98 ( .B1(n152), .B2(n150), .A(STALL), .ZN(n151) );
  NOR2_X1 U99 ( .A1(n34), .A2(n153), .ZN(n150) );
  NAND3_X1 U100 ( .A1(n188), .A2(n155), .A3(n148), .ZN(n34) );
  NOR2_X1 U104 ( .A1(n159), .A2(n183), .ZN(n148) );
  NOR4_X1 U105 ( .A1(n133), .A2(n131), .A3(IR_IN_26), .A4(IR_IN_29), .ZN(n45)
         );
  OR2_X1 U106 ( .A1(n160), .A2(MUXA_SEL), .ZN(JUMP_EN) );
  NAND3_X1 U108 ( .A1(n161), .A2(n155), .A3(n156), .ZN(n145) );
  NAND4_X1 U109 ( .A1(n181), .A2(IR_IN_28), .A3(n2), .A4(n190), .ZN(n156) );
  INV_X1 U110 ( .A(n186), .ZN(n35) );
  AOI21_X1 U111 ( .B1(n162), .B2(n157), .A(n186), .ZN(n160) );
  OAI21_X1 U112 ( .B1(n163), .B2(n187), .A(n164), .ZN(JUMP) );
  INV_X1 U113 ( .A(cw_0), .ZN(n164) );
  AOI21_X1 U114 ( .B1(n162), .B2(n155), .A(n187), .ZN(cw_0) );
  NOR2_X1 U115 ( .A1(n165), .A2(n192), .ZN(I_R_type) );
  NOR4_X1 U116 ( .A1(n166), .A2(n159), .A3(n158), .A4(n153), .ZN(n165) );
  OAI211_X1 U117 ( .C1(n133), .C2(n193), .A(n139), .B(n163), .ZN(n153) );
  AND2_X1 U118 ( .A1(n161), .A2(n157), .ZN(n163) );
  NAND2_X1 U119 ( .A1(n78), .A2(n168), .ZN(n157) );
  NAND2_X1 U120 ( .A1(n169), .A2(n168), .ZN(n161) );
  NAND2_X1 U121 ( .A1(n170), .A2(n171), .ZN(n139) );
  INV_X1 U123 ( .A(n147), .ZN(n172) );
  OAI211_X1 U124 ( .C1(n140), .C2(n173), .A(n49), .B(n39), .ZN(n147) );
  NAND4_X1 U125 ( .A1(IR_IN_31), .A2(IR_IN_27), .A3(n171), .A4(n2), .ZN(n39)
         );
  NOR2_X1 U126 ( .A1(n109), .A2(n131), .ZN(n171) );
  INV_X1 U127 ( .A(n108), .ZN(n131) );
  NOR2_X1 U128 ( .A1(IR_IN_30), .A2(IR_IN_28), .ZN(n108) );
  NAND2_X1 U130 ( .A1(n168), .A2(n174), .ZN(n162) );
  NAND4_X1 U132 ( .A1(n191), .A2(n62), .A3(n68), .A4(n69), .ZN(n176) );
  NAND3_X1 U133 ( .A1(n174), .A2(n194), .A3(n170), .ZN(n69) );
  NAND3_X1 U134 ( .A1(n78), .A2(n194), .A3(n170), .ZN(n68) );
  INV_X1 U136 ( .A(IR_IN_31), .ZN(n40) );
  NAND3_X1 U137 ( .A1(n195), .A2(n174), .A3(n83), .ZN(n62) );
  OAI211_X1 U140 ( .C1(n66), .C2(n86), .A(n61), .B(n67), .ZN(n146) );
  NAND2_X1 U141 ( .A1(n112), .A2(n181), .ZN(n67) );
  NAND3_X1 U142 ( .A1(n112), .A2(n195), .A3(n169), .ZN(n61) );
  OAI22_X1 U143 ( .A1(n173), .A2(n178), .B1(n179), .B2(n66), .ZN(n175) );
  INV_X1 U144 ( .A(n174), .ZN(n66) );
  INV_X1 U146 ( .A(IR_IN_26), .ZN(n109) );
  AOI21_X1 U147 ( .B1(n195), .B2(n83), .A(n180), .ZN(n178) );
  INV_X1 U148 ( .A(n179), .ZN(n180) );
  NAND2_X1 U149 ( .A1(n112), .A2(n184), .ZN(n179) );
  INV_X1 U152 ( .A(n78), .ZN(n173) );
  NAND2_X1 U154 ( .A1(n140), .A2(n86), .ZN(n159) );
  NAND2_X1 U155 ( .A1(IR_IN_29), .A2(n51), .ZN(n86) );
  NAND2_X1 U156 ( .A1(IR_IN_29), .A2(n167), .ZN(n140) );
  INV_X1 U158 ( .A(n155), .ZN(n166) );
  NAND3_X1 U159 ( .A1(IR_IN_26), .A2(n104), .A3(n168), .ZN(n155) );
  NOR2_X1 U160 ( .A1(n117), .A2(IR_IN_29), .ZN(n168) );
  INV_X1 U163 ( .A(IR_IN_27), .ZN(n116) );
  INV_X1 U164 ( .A(IR_IN_30), .ZN(n104) );
  NOR4_X1 U165 ( .A1(n186), .A2(n133), .A3(n193), .A4(n141), .ZN(EQ_COND) );
  INV_X1 U166 ( .A(n169), .ZN(n141) );
  NOR2_X1 U167 ( .A1(IR_IN_30), .A2(IR_IN_26), .ZN(n169) );
  NOR2_X1 U169 ( .A1(n194), .A2(IR_IN_29), .ZN(n83) );
  INV_X1 U170 ( .A(IR_IN_28), .ZN(n52) );
  INV_X1 U171 ( .A(n51), .ZN(n133) );
  NOR2_X1 U172 ( .A1(IR_IN_31), .A2(IR_IN_27), .ZN(n51) );
  INV_X1 U174 ( .A(Flush_BTB), .ZN(n152) );
  INV_X1 U27 ( .A(n107), .ZN(n1) );
  INV_X1 U42 ( .A(n1), .ZN(n2) );
  AOI221_X1 U72 ( .B1(n154), .B2(n2), .C1(n108), .C2(n109), .A(n110), .ZN(n106) );
  CLKBUF_X3 U101 ( .A(n206), .Z(PC_LATCH_EN) );
  INV_X1 U102 ( .A(IR_IN_29), .ZN(n107) );
  AND2_X1 U103 ( .A1(IR_IN_30), .A2(n130), .ZN(n78) );
  INV_X1 U107 ( .A(IR_IN_26), .ZN(n130) );
  NOR3_X2 U122 ( .A1(n40), .A2(n184), .A3(n107), .ZN(n170) );
  NOR2_X2 U129 ( .A1(n109), .A2(n189), .ZN(n174) );
  INV_X1 U131 ( .A(IR_IN_30), .ZN(n149) );
  INV_X1 U135 ( .A(n149), .ZN(n154) );
  AND2_X2 U138 ( .A1(n84), .A2(n52), .ZN(n167) );
  INV_X4 U139 ( .A(n167), .ZN(n117) );
  AOI221_X1 U145 ( .B1(n82), .B2(n78), .C1(n83), .C2(n195), .A(n85), .ZN(n81)
         );
  NOR3_X1 U150 ( .A1(n175), .A2(n146), .A3(n176), .ZN(n177) );
  BUF_X1 U151 ( .A(n51), .Z(n181) );
  INV_X1 U153 ( .A(n45), .ZN(n182) );
  INV_X1 U157 ( .A(n182), .ZN(n183) );
  AOI211_X4 U161 ( .C1(n183), .C2(n136), .A(n137), .B(n138), .ZN(n135) );
  INV_X1 U162 ( .A(IR_IN_27), .ZN(n184) );
  INV_X1 U168 ( .A(n184), .ZN(n185) );
  NAND2_X1 U173 ( .A1(NPC_LATCH_EN), .A2(n152), .ZN(n187) );
  NAND2_X1 U175 ( .A1(NPC_LATCH_EN), .A2(n152), .ZN(n186) );
  NOR2_X4 U176 ( .A1(n239), .A2(STALL), .ZN(NPC_LATCH_EN) );
  NAND2_X1 U177 ( .A1(NPC_LATCH_EN), .A2(n152), .ZN(n37) );
  AND3_X2 U178 ( .A1(n177), .A2(n162), .A3(n172), .ZN(n188) );
  INV_X4 U179 ( .A(n188), .ZN(n158) );
  INV_X1 U180 ( .A(n154), .ZN(n190) );
  INV_X1 U181 ( .A(IR_IN_30), .ZN(n189) );
  AND2_X1 U182 ( .A1(IR_IN_29), .A2(IR_IN_28), .ZN(n112) );
  OR3_X2 U183 ( .A1(n173), .A2(n133), .A3(n193), .ZN(n191) );
  INV_X4 U184 ( .A(n191), .ZN(n122) );
  CLKBUF_X1 U185 ( .A(n186), .Z(n192) );
  OR2_X1 U186 ( .A1(n52), .A2(IR_IN_29), .ZN(n193) );
  INV_X1 U187 ( .A(IR_IN_28), .ZN(n194) );
  BUF_X1 U188 ( .A(n84), .Z(n195) );
  NOR2_X1 U189 ( .A1(n116), .A2(IR_IN_31), .ZN(n84) );
  CLKBUF_X1 U190 ( .A(n147), .Z(n196) );
  CLKBUF_X1 U191 ( .A(MUX_IMM_SEL), .Z(RegA_LATCH_EN) );
  OR2_X2 U192 ( .A1(n66), .A2(n140), .ZN(n49) );
  CLKBUF_X1 U193 ( .A(RegA_LATCH_EN), .Z(RFR1_EN) );
  BUF_X4 U194 ( .A(n205), .Z(MUX_IMM_SEL) );
  AOI21_X1 U195 ( .B1(n156), .B2(n38), .A(n37), .ZN(n205) );
  AND4_X2 U196 ( .A1(n148), .A2(n188), .A3(n157), .A4(n139), .ZN(n38) );
  AND2_X4 U197 ( .A1(n35), .A2(n145), .ZN(MUXA_SEL) );
  DFFR_X1 \cw5_reg[0]  ( .D(\cw4[0] ), .CK(Clk), .RN(Rst), .Q(JandL) );
  DFFR_X1 \cw5_reg[3]  ( .D(cw4_3), .CK(Clk), .RN(Rst), .Q(WB_MUX_SEL) );
  DFFR_X1 \cw4_reg[11]  ( .D(cw3_11), .CK(Clk), .RN(Rst), .Q(RPCplus8_LATCH_EN) );
  DFFR_X1 \cw4_reg[10]  ( .D(cw3_10), .CK(Clk), .RN(Rst), .Q(DRAM_EN) );
  DFFR_X1 \cw4_reg[8]  ( .D(cw3[8]), .CK(Clk), .RN(Rst), .Q(DRAM_WE) );
  DFFR_X1 \cw4_reg[7]  ( .D(cw3[7]), .CK(Clk), .RN(Rst), .Q(LMD_LATCH_EN) );
  DFFR_X1 \cw4_reg[6]  ( .D(cw3[6]), .CK(Clk), .RN(Rst), .Q(RALUOUT2_LATCH_EN)
         );
  DFFR_X1 \cw4_reg[5]  ( .D(cw3[5]), .CK(Clk), .RN(Rst), .Q(RegRD3_LATCH_EN)
         );
  DFFR_X1 \cw4_reg[3]  ( .D(cw3_3), .CK(Clk), .RN(Rst), .Q(cw4_3) );
  DFFR_X1 \cw4_reg[0]  ( .D(cw3_0), .CK(Clk), .RN(Rst), .Q(\cw4[0] ) );
  DFFR_X1 \cw4_reg[2]  ( .D(REGWRITE_DX), .CK(Clk), .RN(Rst), .Q(REGWRITE_XM)
         );
  DFFR_X1 \cw4_reg[9]  ( .D(MEMREAD_DX), .CK(Clk), .RN(Rst), .Q(DRAM_RE) );
  DFFR_X1 \cw5_reg[2]  ( .D(REGWRITE_XM), .CK(Clk), .RN(Rst), .Q(REGWRITE_MW)
         );
  DFFR_X1 \aluOpcode3_reg[3]  ( .D(aluOpcode_i[3]), .CK(Clk), .RN(Rst), .Q(
        ALU_OPCODE[3]) );
  DFFR_X1 \aluOpcode3_reg[0]  ( .D(aluOpcode_i[0]), .CK(Clk), .RN(Rst), .Q(
        ALU_OPCODE[0]) );
  DFFR_X1 \aluOpcode3_reg[2]  ( .D(aluOpcode_i[2]), .CK(Clk), .RN(Rst), .Q(
        ALU_OPCODE[2]) );
  DFFR_X1 \cw3_reg[11]  ( .D(cw_0), .CK(Clk), .RN(Rst), .Q(cw3_11) );
  DFFR_X1 \cw3_reg[0]  ( .D(cw_0), .CK(Clk), .RN(Rst), .Q(cw3_0) );
  DFFR_X1 \cw3_reg[2]  ( .D(cw_2), .CK(Clk), .RN(Rst), .Q(REGWRITE_DX) );
  DFFR_X1 \cw3_reg[15]  ( .D(cw[15]), .CK(Clk), .RN(Rst), .Q(MUXB_SEL) );
  DFFR_X1 \cw3_reg[13]  ( .D(cw[13]), .CK(Clk), .RN(Rst), .Q(ALU_OUTREG_EN) );
  DFFR_X1 \cw3_reg[6]  ( .D(cw[6]), .CK(Clk), .RN(Rst), .Q(cw3[6]) );
  DFFR_X1 \cw3_reg[8]  ( .D(cw[8]), .CK(Clk), .RN(Rst), .Q(cw3[8]) );
  DFFR_X1 \cw3_reg[12]  ( .D(cw[5]), .CK(Clk), .RN(Rst), .Q(RegRD2_LATCH_EN)
         );
  DFFR_X1 \cw3_reg[5]  ( .D(cw[5]), .CK(Clk), .RN(Rst), .Q(cw3[5]) );
  DFFR_X1 \cw3_reg[9]  ( .D(cw_3), .CK(Clk), .RN(Rst), .Q(MEMREAD_DX) );
  DFFR_X1 \cw3_reg[7]  ( .D(cw_3), .CK(Clk), .RN(Rst), .Q(cw3[7]) );
  DFFR_X1 \cw3_reg[3]  ( .D(cw_3), .CK(Clk), .RN(Rst), .Q(cw3_3) );
  DFFR_X1 \cw3_reg[14]  ( .D(cw[14]), .CK(Clk), .RN(Rst), .Q(REGME_LATCH_EN)
         );
  DFFR_X1 \cw3_reg[10]  ( .D(cw[14]), .CK(Clk), .RN(Rst), .Q(cw3_10) );
  INV_X1 U198 ( .A(n239), .ZN(REGF_LATCH_EN) );
  INV_X1 U199 ( .A(n239), .ZN(n238) );
  INV_X2 U200 ( .A(Rst), .ZN(n239) );
endmodule


module NPC_logic_PC_SIZE32 ( Flush_BTB, BRANCH_CTRL_SIG, OUTT_NT_i, PC_next, 
        BRANCH_ALU_OUT, OUT_PC_target_i, NPC, PC_BUS );
  input [31:0] PC_next;
  input [31:0] BRANCH_ALU_OUT;
  input [31:0] OUT_PC_target_i;
  input [31:0] NPC;
  output [31:0] PC_BUS;
  input Flush_BTB, BRANCH_CTRL_SIG, OUTT_NT_i;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n20, n1, n71,
         n72, n73;

  NAND2_X1 U1 ( .A1(n2), .A2(n3), .ZN(PC_BUS[9]) );
  AOI22_X1 U2 ( .A1(NPC[9]), .A2(n73), .B1(BRANCH_ALU_OUT[9]), .B2(n71), .ZN(
        n3) );
  AOI22_X1 U3 ( .A1(PC_next[9]), .A2(n6), .B1(OUT_PC_target_i[9]), .B2(n7), 
        .ZN(n2) );
  NAND2_X1 U4 ( .A1(n8), .A2(n9), .ZN(PC_BUS[8]) );
  AOI22_X1 U5 ( .A1(NPC[8]), .A2(n73), .B1(BRANCH_ALU_OUT[8]), .B2(n71), .ZN(
        n9) );
  AOI22_X1 U6 ( .A1(PC_next[8]), .A2(n6), .B1(OUT_PC_target_i[8]), .B2(n7), 
        .ZN(n8) );
  NAND2_X1 U7 ( .A1(n10), .A2(n11), .ZN(PC_BUS[7]) );
  AOI22_X1 U8 ( .A1(NPC[7]), .A2(n73), .B1(BRANCH_ALU_OUT[7]), .B2(n71), .ZN(
        n11) );
  AOI22_X1 U9 ( .A1(PC_next[7]), .A2(n6), .B1(OUT_PC_target_i[7]), .B2(n7), 
        .ZN(n10) );
  NAND2_X1 U10 ( .A1(n12), .A2(n13), .ZN(PC_BUS[6]) );
  AOI22_X1 U11 ( .A1(NPC[6]), .A2(n73), .B1(BRANCH_ALU_OUT[6]), .B2(n71), .ZN(
        n13) );
  AOI22_X1 U12 ( .A1(PC_next[6]), .A2(n6), .B1(OUT_PC_target_i[6]), .B2(n7), 
        .ZN(n12) );
  NAND2_X1 U13 ( .A1(n14), .A2(n15), .ZN(PC_BUS[5]) );
  AOI22_X1 U14 ( .A1(NPC[5]), .A2(n73), .B1(BRANCH_ALU_OUT[5]), .B2(n71), .ZN(
        n15) );
  AOI22_X1 U15 ( .A1(PC_next[5]), .A2(n6), .B1(OUT_PC_target_i[5]), .B2(n7), 
        .ZN(n14) );
  NAND2_X1 U16 ( .A1(n16), .A2(n17), .ZN(PC_BUS[4]) );
  AOI22_X1 U17 ( .A1(NPC[4]), .A2(n73), .B1(BRANCH_ALU_OUT[4]), .B2(n71), .ZN(
        n17) );
  AOI22_X1 U18 ( .A1(PC_next[4]), .A2(n6), .B1(OUT_PC_target_i[4]), .B2(n7), 
        .ZN(n16) );
  NAND2_X1 U19 ( .A1(n18), .A2(n19), .ZN(PC_BUS[3]) );
  AOI22_X1 U20 ( .A1(NPC[3]), .A2(n73), .B1(BRANCH_ALU_OUT[3]), .B2(n71), .ZN(
        n19) );
  AOI22_X1 U21 ( .A1(PC_next[3]), .A2(n6), .B1(OUT_PC_target_i[3]), .B2(n7), 
        .ZN(n18) );
  AOI22_X1 U23 ( .A1(NPC[31]), .A2(n73), .B1(BRANCH_ALU_OUT[31]), .B2(n71), 
        .ZN(n21) );
  NAND2_X1 U25 ( .A1(n23), .A2(n22), .ZN(PC_BUS[30]) );
  AOI22_X1 U26 ( .A1(NPC[30]), .A2(n73), .B1(BRANCH_ALU_OUT[30]), .B2(n71), 
        .ZN(n23) );
  AOI22_X1 U27 ( .A1(PC_next[30]), .A2(n6), .B1(OUT_PC_target_i[30]), .B2(n7), 
        .ZN(n22) );
  NAND2_X1 U28 ( .A1(n24), .A2(n25), .ZN(PC_BUS[2]) );
  AOI22_X1 U29 ( .A1(NPC[2]), .A2(n73), .B1(BRANCH_ALU_OUT[2]), .B2(n71), .ZN(
        n25) );
  AOI22_X1 U30 ( .A1(PC_next[2]), .A2(n6), .B1(OUT_PC_target_i[2]), .B2(n7), 
        .ZN(n24) );
  NAND2_X1 U31 ( .A1(n26), .A2(n27), .ZN(PC_BUS[29]) );
  AOI22_X1 U32 ( .A1(NPC[29]), .A2(n73), .B1(BRANCH_ALU_OUT[29]), .B2(n71), 
        .ZN(n27) );
  AOI22_X1 U33 ( .A1(PC_next[29]), .A2(n6), .B1(OUT_PC_target_i[29]), .B2(n7), 
        .ZN(n26) );
  NAND2_X1 U34 ( .A1(n28), .A2(n29), .ZN(PC_BUS[28]) );
  AOI22_X1 U35 ( .A1(NPC[28]), .A2(n73), .B1(BRANCH_ALU_OUT[28]), .B2(n71), 
        .ZN(n29) );
  AOI22_X1 U36 ( .A1(PC_next[28]), .A2(n6), .B1(OUT_PC_target_i[28]), .B2(n7), 
        .ZN(n28) );
  NAND2_X1 U37 ( .A1(n30), .A2(n31), .ZN(PC_BUS[27]) );
  AOI22_X1 U38 ( .A1(NPC[27]), .A2(n73), .B1(BRANCH_ALU_OUT[27]), .B2(n71), 
        .ZN(n31) );
  AOI22_X1 U39 ( .A1(PC_next[27]), .A2(n6), .B1(OUT_PC_target_i[27]), .B2(n7), 
        .ZN(n30) );
  NAND2_X1 U40 ( .A1(n32), .A2(n33), .ZN(PC_BUS[26]) );
  AOI22_X1 U41 ( .A1(NPC[26]), .A2(n73), .B1(BRANCH_ALU_OUT[26]), .B2(n71), 
        .ZN(n33) );
  AOI22_X1 U42 ( .A1(PC_next[26]), .A2(n6), .B1(OUT_PC_target_i[26]), .B2(n7), 
        .ZN(n32) );
  NAND2_X1 U43 ( .A1(n34), .A2(n35), .ZN(PC_BUS[25]) );
  AOI22_X1 U44 ( .A1(NPC[25]), .A2(n73), .B1(BRANCH_ALU_OUT[25]), .B2(n71), 
        .ZN(n35) );
  AOI22_X1 U45 ( .A1(PC_next[25]), .A2(n6), .B1(OUT_PC_target_i[25]), .B2(n7), 
        .ZN(n34) );
  NAND2_X1 U46 ( .A1(n36), .A2(n37), .ZN(PC_BUS[24]) );
  AOI22_X1 U47 ( .A1(NPC[24]), .A2(n73), .B1(BRANCH_ALU_OUT[24]), .B2(n71), 
        .ZN(n37) );
  AOI22_X1 U48 ( .A1(PC_next[24]), .A2(n6), .B1(OUT_PC_target_i[24]), .B2(n7), 
        .ZN(n36) );
  NAND2_X1 U49 ( .A1(n38), .A2(n39), .ZN(PC_BUS[23]) );
  AOI22_X1 U50 ( .A1(NPC[23]), .A2(n73), .B1(BRANCH_ALU_OUT[23]), .B2(n71), 
        .ZN(n39) );
  AOI22_X1 U51 ( .A1(PC_next[23]), .A2(n6), .B1(OUT_PC_target_i[23]), .B2(n7), 
        .ZN(n38) );
  NAND2_X1 U52 ( .A1(n40), .A2(n41), .ZN(PC_BUS[22]) );
  AOI22_X1 U53 ( .A1(NPC[22]), .A2(n73), .B1(BRANCH_ALU_OUT[22]), .B2(n71), 
        .ZN(n41) );
  AOI22_X1 U54 ( .A1(PC_next[22]), .A2(n6), .B1(OUT_PC_target_i[22]), .B2(n7), 
        .ZN(n40) );
  NAND2_X1 U55 ( .A1(n42), .A2(n43), .ZN(PC_BUS[21]) );
  AOI22_X1 U56 ( .A1(NPC[21]), .A2(n73), .B1(BRANCH_ALU_OUT[21]), .B2(n71), 
        .ZN(n43) );
  AOI22_X1 U57 ( .A1(PC_next[21]), .A2(n6), .B1(OUT_PC_target_i[21]), .B2(n7), 
        .ZN(n42) );
  NAND2_X1 U58 ( .A1(n44), .A2(n45), .ZN(PC_BUS[20]) );
  AOI22_X1 U59 ( .A1(NPC[20]), .A2(n73), .B1(BRANCH_ALU_OUT[20]), .B2(n71), 
        .ZN(n45) );
  AOI22_X1 U60 ( .A1(PC_next[20]), .A2(n6), .B1(OUT_PC_target_i[20]), .B2(n7), 
        .ZN(n44) );
  NAND2_X1 U61 ( .A1(n46), .A2(n47), .ZN(PC_BUS[1]) );
  AOI22_X1 U62 ( .A1(NPC[1]), .A2(n73), .B1(BRANCH_ALU_OUT[1]), .B2(n71), .ZN(
        n47) );
  AOI22_X1 U63 ( .A1(PC_next[1]), .A2(n6), .B1(OUT_PC_target_i[1]), .B2(n7), 
        .ZN(n46) );
  NAND2_X1 U64 ( .A1(n49), .A2(n48), .ZN(PC_BUS[19]) );
  AOI22_X1 U65 ( .A1(NPC[19]), .A2(n73), .B1(BRANCH_ALU_OUT[19]), .B2(n71), 
        .ZN(n49) );
  AOI22_X1 U66 ( .A1(PC_next[19]), .A2(n6), .B1(OUT_PC_target_i[19]), .B2(n7), 
        .ZN(n48) );
  NAND2_X1 U67 ( .A1(n50), .A2(n51), .ZN(PC_BUS[18]) );
  AOI22_X1 U68 ( .A1(NPC[18]), .A2(n73), .B1(BRANCH_ALU_OUT[18]), .B2(n71), 
        .ZN(n51) );
  AOI22_X1 U69 ( .A1(PC_next[18]), .A2(n6), .B1(OUT_PC_target_i[18]), .B2(n7), 
        .ZN(n50) );
  NAND2_X1 U70 ( .A1(n52), .A2(n53), .ZN(PC_BUS[17]) );
  AOI22_X1 U71 ( .A1(NPC[17]), .A2(n73), .B1(BRANCH_ALU_OUT[17]), .B2(n71), 
        .ZN(n53) );
  AOI22_X1 U72 ( .A1(PC_next[17]), .A2(n6), .B1(OUT_PC_target_i[17]), .B2(n7), 
        .ZN(n52) );
  NAND2_X1 U73 ( .A1(n54), .A2(n55), .ZN(PC_BUS[16]) );
  AOI22_X1 U74 ( .A1(NPC[16]), .A2(n73), .B1(BRANCH_ALU_OUT[16]), .B2(n71), 
        .ZN(n55) );
  AOI22_X1 U75 ( .A1(PC_next[16]), .A2(n6), .B1(OUT_PC_target_i[16]), .B2(n7), 
        .ZN(n54) );
  NAND2_X1 U76 ( .A1(n56), .A2(n57), .ZN(PC_BUS[15]) );
  AOI22_X1 U77 ( .A1(NPC[15]), .A2(n73), .B1(BRANCH_ALU_OUT[15]), .B2(n71), 
        .ZN(n57) );
  AOI22_X1 U78 ( .A1(PC_next[15]), .A2(n6), .B1(OUT_PC_target_i[15]), .B2(n7), 
        .ZN(n56) );
  NAND2_X1 U79 ( .A1(n58), .A2(n59), .ZN(PC_BUS[14]) );
  AOI22_X1 U80 ( .A1(NPC[14]), .A2(n73), .B1(BRANCH_ALU_OUT[14]), .B2(n71), 
        .ZN(n59) );
  AOI22_X1 U81 ( .A1(PC_next[14]), .A2(n6), .B1(OUT_PC_target_i[14]), .B2(n7), 
        .ZN(n58) );
  NAND2_X1 U82 ( .A1(n60), .A2(n61), .ZN(PC_BUS[13]) );
  AOI22_X1 U83 ( .A1(NPC[13]), .A2(n73), .B1(BRANCH_ALU_OUT[13]), .B2(n71), 
        .ZN(n61) );
  AOI22_X1 U84 ( .A1(PC_next[13]), .A2(n6), .B1(OUT_PC_target_i[13]), .B2(n7), 
        .ZN(n60) );
  NAND2_X1 U85 ( .A1(n62), .A2(n63), .ZN(PC_BUS[12]) );
  AOI22_X1 U86 ( .A1(NPC[12]), .A2(n73), .B1(BRANCH_ALU_OUT[12]), .B2(n71), 
        .ZN(n63) );
  AOI22_X1 U87 ( .A1(PC_next[12]), .A2(n6), .B1(OUT_PC_target_i[12]), .B2(n7), 
        .ZN(n62) );
  NAND2_X1 U88 ( .A1(n64), .A2(n65), .ZN(PC_BUS[11]) );
  AOI22_X1 U89 ( .A1(NPC[11]), .A2(n73), .B1(BRANCH_ALU_OUT[11]), .B2(n71), 
        .ZN(n65) );
  AOI22_X1 U90 ( .A1(PC_next[11]), .A2(n6), .B1(OUT_PC_target_i[11]), .B2(n7), 
        .ZN(n64) );
  NAND2_X1 U91 ( .A1(n66), .A2(n67), .ZN(PC_BUS[10]) );
  AOI22_X1 U92 ( .A1(NPC[10]), .A2(n73), .B1(BRANCH_ALU_OUT[10]), .B2(n71), 
        .ZN(n67) );
  AOI22_X1 U93 ( .A1(PC_next[10]), .A2(n6), .B1(OUT_PC_target_i[10]), .B2(n7), 
        .ZN(n66) );
  NAND2_X1 U94 ( .A1(n68), .A2(n69), .ZN(PC_BUS[0]) );
  AOI22_X1 U95 ( .A1(NPC[0]), .A2(n73), .B1(BRANCH_ALU_OUT[0]), .B2(n71), .ZN(
        n69) );
  AOI22_X1 U98 ( .A1(PC_next[0]), .A2(n6), .B1(OUT_PC_target_i[0]), .B2(n7), 
        .ZN(n68) );
  AND2_X1 U96 ( .A1(BRANCH_CTRL_SIG), .A2(Flush_BTB), .ZN(n5) );
  INV_X1 U100 ( .A(Flush_BTB), .ZN(n70) );
  NAND2_X1 U22 ( .A1(n20), .A2(n21), .ZN(PC_BUS[31]) );
  AOI22_X1 U24 ( .A1(PC_next[31]), .A2(n6), .B1(OUT_PC_target_i[31]), .B2(n7), 
        .ZN(n20) );
  INV_X1 U97 ( .A(n5), .ZN(n1) );
  INV_X2 U99 ( .A(n1), .ZN(n71) );
  NOR2_X4 U101 ( .A1(Flush_BTB), .A2(OUTT_NT_i), .ZN(n6) );
  AND2_X4 U102 ( .A1(OUTT_NT_i), .A2(n70), .ZN(n7) );
  INV_X1 U103 ( .A(n4), .ZN(n72) );
  INV_X2 U104 ( .A(n72), .ZN(n73) );
  NOR2_X1 U105 ( .A1(n70), .A2(BRANCH_CTRL_SIG), .ZN(n4) );
endmodule


module DLX_IR_SIZE32_PC_SIZE32 ( Clk, Rst, Iaddr, Idata, Denable, Drd, Dwd, 
        Daddr, Ddatain, Ddataout, DataOut );
  output [31:0] Iaddr;
  input [31:0] Idata;
  output [31:0] Daddr;
  output [31:0] Ddatain;
  input [31:0] Ddataout;
  output [31:0] DataOut;
  input Clk, Rst;
  output Denable, Drd, Dwd;
  wire   n314, I_R_TYPE_i, N2, prevT_NT_i, Flush_BTB_i, BRANCH_CTRL_SIG,
         Flush_BTB, IR_LATCH_EN_i, PC_LATCH_EN_i, NPC_LATCH_EN_i, OUTT_NT_i,
         STALL_i, RegRF_LATCH_EN_i, RegA_LATCH_EN_i, RegB_LATCH_EN_i,
         RegIMM_LATCH_EN_i, RegRD1_LATCH_EN_i, SIGN_UNSIGN_i, RFR1_EN_i,
         RFR2_EN_i, MUX_IMM_SEL_i, JUMP_i, JUMP_EN_i, EQ_COND_i, MUXA_SEL_i,
         MUXB_SEL_i, ALU_OUTREG_EN_i, REGME_LATCH_EN_i, RegRD2_LATCH_EN_i,
         LMD_LATCH_EN_i, RALUOUT2_LATCH_EN_i, RegRD3_LATCH_EN_i,
         RPCplus8_LATCH_EN_i, WB_MUX_SEL_i, RF_WE_i, JandL_i, REGWRITE_DX_i,
         REGWRITE_XM_i, REGWRITE_MW_i, MEMREAD_DX_i, N4, N5, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313;
  wire   [15:0] INP2;
  wire   [31:26] IR;
  wire   [25:16] IMM26;
  wire   [4:0] RD;
  wire   [31:0] PC_BUS;
  wire   [31:0] NPC;
  wire   [31:0] PC_next;
  wire   [31:0] BRANCH_ALU_OUT;
  wire   [31:0] OUT_PC_target_i;
  wire   [4:0] ALU_OPCODE_i;

  AND2_X2 C628 ( .A1(prevT_NT_i), .A2(N4), .ZN(N5) );
  XOR2_X1 C627 ( .A(N5), .B(BRANCH_CTRL_SIG), .Z(Flush_BTB) );
  INV_X2 I_1 ( .A(I_R_TYPE_i), .ZN(N2) );
  DFFR_X1 \NPC_reg[0]  ( .D(n289), .CK(Clk), .RN(n311), .Q(NPC[0]), .QN(n193)
         );
  DFFR_X1 Flush_BTB_i_reg ( .D(Flush_BTB), .CK(Clk), .RN(n313), .Q(Flush_BTB_i), .QN(N4) );
  DFFR_X1 \PC_reg[0]  ( .D(n287), .CK(Clk), .RN(n313), .Q(n314), .QN(n191) );
  DFFR_X1 \PC_reg[1]  ( .D(n286), .CK(Clk), .RN(n312), .Q(Iaddr[1]), .QN(n190)
         );
  DFFR_X1 \PC_reg[2]  ( .D(n285), .CK(Clk), .RN(n312), .Q(Iaddr[2]), .QN(n189)
         );
  DFFR_X1 \PC_reg[3]  ( .D(n284), .CK(Clk), .RN(n313), .Q(Iaddr[3]), .QN(n188)
         );
  DFFR_X1 \PC_reg[4]  ( .D(n283), .CK(Clk), .RN(n313), .Q(Iaddr[4]), .QN(n187)
         );
  DFFR_X1 \PC_reg[5]  ( .D(n282), .CK(Clk), .RN(n313), .Q(Iaddr[5]), .QN(n186)
         );
  DFFR_X1 \PC_reg[6]  ( .D(n281), .CK(Clk), .RN(n313), .Q(Iaddr[6]), .QN(n185)
         );
  DFFR_X1 \PC_reg[7]  ( .D(n280), .CK(Clk), .RN(n313), .Q(Iaddr[7]), .QN(n184)
         );
  DFFR_X1 \PC_reg[8]  ( .D(n279), .CK(Clk), .RN(n313), .Q(Iaddr[8]), .QN(n183)
         );
  DFFR_X1 \PC_reg[9]  ( .D(n278), .CK(Clk), .RN(n313), .Q(Iaddr[9]), .QN(n182)
         );
  DFFR_X1 \PC_reg[10]  ( .D(n277), .CK(Clk), .RN(n312), .Q(Iaddr[10]), .QN(
        n181) );
  DFFR_X1 \PC_reg[11]  ( .D(n276), .CK(Clk), .RN(n311), .Q(Iaddr[11]), .QN(
        n180) );
  DFFR_X1 \PC_reg[12]  ( .D(n275), .CK(Clk), .RN(n311), .Q(Iaddr[12]), .QN(
        n179) );
  DFFR_X1 \PC_reg[13]  ( .D(n274), .CK(Clk), .RN(n311), .Q(Iaddr[13]), .QN(
        n178) );
  DFFR_X1 \PC_reg[14]  ( .D(n273), .CK(Clk), .RN(n311), .Q(Iaddr[14]), .QN(
        n177) );
  DFFR_X1 \PC_reg[15]  ( .D(n272), .CK(Clk), .RN(n311), .Q(Iaddr[15]), .QN(
        n176) );
  DFFR_X1 \PC_reg[16]  ( .D(n271), .CK(Clk), .RN(n311), .Q(Iaddr[16]), .QN(
        n175) );
  DFFR_X1 \PC_reg[17]  ( .D(n270), .CK(Clk), .RN(n311), .Q(Iaddr[17]), .QN(
        n174) );
  DFFR_X1 \PC_reg[18]  ( .D(n269), .CK(Clk), .RN(n311), .Q(Iaddr[18]), .QN(
        n173) );
  DFFR_X1 \PC_reg[19]  ( .D(n268), .CK(Clk), .RN(n311), .Q(Iaddr[19]), .QN(
        n172) );
  DFFR_X1 \PC_reg[20]  ( .D(n267), .CK(Clk), .RN(n311), .Q(Iaddr[20]), .QN(
        n171) );
  DFFR_X1 \PC_reg[21]  ( .D(n266), .CK(Clk), .RN(n312), .Q(Iaddr[21]), .QN(
        n170) );
  DFFR_X1 \PC_reg[22]  ( .D(n265), .CK(Clk), .RN(n311), .Q(Iaddr[22]), .QN(
        n169) );
  DFFR_X1 \PC_reg[23]  ( .D(n264), .CK(Clk), .RN(n312), .Q(Iaddr[23]), .QN(
        n168) );
  DFFR_X1 \PC_reg[24]  ( .D(n263), .CK(Clk), .RN(n311), .Q(Iaddr[24]), .QN(
        n167) );
  DFFR_X1 \PC_reg[25]  ( .D(n262), .CK(Clk), .RN(n312), .Q(Iaddr[25]), .QN(
        n166) );
  DFFR_X1 \PC_reg[26]  ( .D(n261), .CK(Clk), .RN(n311), .Q(Iaddr[26]), .QN(
        n165) );
  DFFR_X1 \PC_reg[27]  ( .D(n260), .CK(Clk), .RN(n312), .Q(Iaddr[27]), .QN(
        n164) );
  DFFR_X1 \PC_reg[28]  ( .D(n259), .CK(Clk), .RN(n313), .Q(Iaddr[28]), .QN(
        n163) );
  DFFR_X1 \PC_reg[29]  ( .D(n258), .CK(Clk), .RN(n312), .Q(Iaddr[29]), .QN(
        n162) );
  DFFR_X1 \PC_reg[30]  ( .D(n257), .CK(Clk), .RN(n311), .Q(Iaddr[30]), .QN(
        n161) );
  DFFR_X1 \NPC_reg[1]  ( .D(n256), .CK(Clk), .RN(n312), .Q(NPC[1]), .QN(n160)
         );
  DFFR_X1 \NPC_reg[2]  ( .D(n255), .CK(Clk), .RN(n312), .Q(NPC[2]), .QN(n159)
         );
  DFFR_X1 \NPC_reg[3]  ( .D(n254), .CK(Clk), .RN(n312), .Q(NPC[3]), .QN(n158)
         );
  DFFR_X1 \NPC_reg[4]  ( .D(n253), .CK(Clk), .RN(n313), .Q(NPC[4]), .QN(n157)
         );
  DFFR_X1 \NPC_reg[5]  ( .D(n252), .CK(Clk), .RN(n313), .Q(NPC[5]), .QN(n156)
         );
  DFFR_X1 \NPC_reg[6]  ( .D(n251), .CK(Clk), .RN(n313), .Q(NPC[6]), .QN(n155)
         );
  DFFR_X1 \NPC_reg[7]  ( .D(n250), .CK(Clk), .RN(n313), .Q(NPC[7]), .QN(n154)
         );
  DFFR_X1 \NPC_reg[8]  ( .D(n249), .CK(Clk), .RN(n313), .Q(NPC[8]), .QN(n153)
         );
  DFFR_X1 \NPC_reg[9]  ( .D(n248), .CK(Clk), .RN(n313), .Q(NPC[9]), .QN(n152)
         );
  DFFR_X1 \NPC_reg[10]  ( .D(n247), .CK(Clk), .RN(n311), .Q(NPC[10]), .QN(n151) );
  DFFR_X1 \NPC_reg[11]  ( .D(n246), .CK(Clk), .RN(n311), .Q(NPC[11]), .QN(n150) );
  DFFR_X1 \NPC_reg[12]  ( .D(n245), .CK(Clk), .RN(n311), .Q(NPC[12]), .QN(n149) );
  DFFR_X1 \NPC_reg[13]  ( .D(n244), .CK(Clk), .RN(n311), .Q(NPC[13]), .QN(n148) );
  DFFR_X1 \NPC_reg[14]  ( .D(n243), .CK(Clk), .RN(n311), .Q(NPC[14]), .QN(n147) );
  DFFR_X1 \NPC_reg[15]  ( .D(n242), .CK(Clk), .RN(n311), .Q(NPC[15]), .QN(n146) );
  DFFR_X1 \NPC_reg[16]  ( .D(n241), .CK(Clk), .RN(n311), .Q(NPC[16]), .QN(n145) );
  DFFR_X1 \NPC_reg[17]  ( .D(n240), .CK(Clk), .RN(n311), .Q(NPC[17]), .QN(n144) );
  DFFR_X1 \NPC_reg[18]  ( .D(n239), .CK(Clk), .RN(n311), .Q(NPC[18]), .QN(n143) );
  DFFR_X1 \NPC_reg[19]  ( .D(n238), .CK(Clk), .RN(n311), .Q(NPC[19]), .QN(n142) );
  DFFR_X1 \NPC_reg[20]  ( .D(n237), .CK(Clk), .RN(n311), .Q(NPC[20]), .QN(n141) );
  DFFR_X1 \NPC_reg[21]  ( .D(n236), .CK(Clk), .RN(n312), .Q(NPC[21]), .QN(n140) );
  DFFR_X1 \NPC_reg[22]  ( .D(n235), .CK(Clk), .RN(n311), .Q(NPC[22]), .QN(n139) );
  DFFR_X1 \NPC_reg[23]  ( .D(n234), .CK(Clk), .RN(n312), .Q(NPC[23]), .QN(n138) );
  DFFR_X1 \NPC_reg[24]  ( .D(n233), .CK(Clk), .RN(n311), .Q(NPC[24]), .QN(n137) );
  DFFR_X1 \NPC_reg[25]  ( .D(n232), .CK(Clk), .RN(n312), .Q(NPC[25]), .QN(n136) );
  DFFR_X1 \NPC_reg[26]  ( .D(n231), .CK(Clk), .RN(n311), .Q(NPC[26]), .QN(n135) );
  DFFR_X1 \NPC_reg[27]  ( .D(n230), .CK(Clk), .RN(n312), .Q(NPC[27]), .QN(n134) );
  DFFR_X1 \NPC_reg[28]  ( .D(n229), .CK(Clk), .RN(n313), .Q(NPC[28]), .QN(n133) );
  DFFR_X1 \NPC_reg[29]  ( .D(n228), .CK(Clk), .RN(n312), .Q(NPC[29]), .QN(n132) );
  DFFR_X1 \NPC_reg[30]  ( .D(n227), .CK(Clk), .RN(n311), .Q(NPC[30]), .QN(n131) );
  DFFR_X1 \NPC_reg[31]  ( .D(n226), .CK(Clk), .RN(n313), .Q(NPC[31]), .QN(n130) );
  DFFR_X1 \IR_reg[0]  ( .D(n225), .CK(Clk), .RN(n312), .Q(INP2[0]), .QN(n129)
         );
  DFFR_X1 \IR_reg[1]  ( .D(n224), .CK(Clk), .RN(n312), .Q(INP2[1]), .QN(n128)
         );
  DFFR_X1 \IR_reg[2]  ( .D(n223), .CK(Clk), .RN(n312), .Q(INP2[2]), .QN(n127)
         );
  DFFR_X1 \IR_reg[3]  ( .D(n222), .CK(Clk), .RN(n312), .Q(INP2[3]), .QN(n126)
         );
  DFFR_X1 \IR_reg[4]  ( .D(n221), .CK(Clk), .RN(n312), .Q(INP2[4]), .QN(n125)
         );
  DFFR_X1 \IR_reg[5]  ( .D(n220), .CK(Clk), .RN(n312), .Q(INP2[5]), .QN(n124)
         );
  DFFR_X1 \IR_reg[6]  ( .D(n219), .CK(Clk), .RN(n312), .Q(INP2[6]), .QN(n123)
         );
  DFFR_X1 \IR_reg[7]  ( .D(n218), .CK(Clk), .RN(n312), .Q(INP2[7]), .QN(n122)
         );
  DFFR_X1 \IR_reg[8]  ( .D(n217), .CK(Clk), .RN(n312), .Q(INP2[8]), .QN(n121)
         );
  DFFR_X1 \IR_reg[9]  ( .D(n216), .CK(Clk), .RN(n312), .Q(INP2[9]), .QN(n120)
         );
  DFFR_X1 \IR_reg[10]  ( .D(n215), .CK(Clk), .RN(n312), .Q(INP2[10]), .QN(n119) );
  DFFR_X1 \IR_reg[11]  ( .D(n214), .CK(Clk), .RN(n312), .Q(INP2[11]), .QN(n118) );
  DFFR_X1 \IR_reg[12]  ( .D(n213), .CK(Clk), .RN(n312), .Q(INP2[12]), .QN(n117) );
  DFFR_X1 \IR_reg[13]  ( .D(n212), .CK(Clk), .RN(n312), .Q(INP2[13]), .QN(n116) );
  DFFR_X1 \IR_reg[14]  ( .D(n211), .CK(Clk), .RN(n312), .Q(INP2[14]), .QN(n115) );
  DFFR_X1 \IR_reg[15]  ( .D(n210), .CK(Clk), .RN(n312), .Q(INP2[15]), .QN(n114) );
  DFFR_X1 \IR_reg[16]  ( .D(n209), .CK(Clk), .RN(n312), .Q(IMM26[16]), .QN(
        n113) );
  DFFR_X1 \IR_reg[17]  ( .D(n208), .CK(Clk), .RN(n312), .Q(IMM26[17]), .QN(
        n112) );
  DFFR_X1 \IR_reg[18]  ( .D(n207), .CK(Clk), .RN(n312), .Q(IMM26[18]), .QN(
        n111) );
  DFFR_X1 \IR_reg[19]  ( .D(n206), .CK(Clk), .RN(n312), .Q(IMM26[19]), .QN(
        n110) );
  DFFR_X1 \IR_reg[20]  ( .D(n205), .CK(Clk), .RN(n312), .Q(IMM26[20]), .QN(
        n109) );
  DFFR_X1 \IR_reg[21]  ( .D(n204), .CK(Clk), .RN(n312), .Q(IMM26[21]), .QN(
        n108) );
  DFFR_X1 \IR_reg[22]  ( .D(n203), .CK(Clk), .RN(n312), .Q(IMM26[22]), .QN(
        n107) );
  DFFR_X1 \IR_reg[23]  ( .D(n202), .CK(Clk), .RN(n312), .Q(IMM26[23]), .QN(
        n106) );
  DFFR_X1 \IR_reg[24]  ( .D(n201), .CK(Clk), .RN(n312), .Q(IMM26[24]), .QN(
        n105) );
  DFFR_X1 \IR_reg[25]  ( .D(n200), .CK(Clk), .RN(n312), .Q(IMM26[25]), .QN(
        n104) );
  DFFR_X1 \IR_reg[26]  ( .D(n199), .CK(Clk), .RN(n312), .Q(IR[26]), .QN(n103)
         );
  DFFR_X1 \IR_reg[27]  ( .D(n198), .CK(Clk), .RN(n312), .Q(IR[27]), .QN(n102)
         );
  DFFR_X1 \IR_reg[28]  ( .D(n197), .CK(Clk), .RN(n312), .Q(IR[28]), .QN(n101)
         );
  DFFR_X1 \IR_reg[29]  ( .D(n196), .CK(Clk), .RN(n312), .Q(IR[29]), .QN(n100)
         );
  DFFR_X1 \IR_reg[30]  ( .D(n195), .CK(Clk), .RN(n313), .Q(IR[30]), .QN(n99)
         );
  DFFR_X1 \IR_reg[31]  ( .D(n194), .CK(Clk), .RN(n313), .Q(IR[31]), .QN(n98)
         );
  OAI21_X1 U3 ( .B1(n304), .B2(n98), .A(n2), .ZN(n194) );
  NAND2_X1 U4 ( .A1(Idata[31]), .A2(n301), .ZN(n2) );
  OAI21_X1 U5 ( .B1(n304), .B2(n99), .A(n3), .ZN(n195) );
  NAND2_X1 U6 ( .A1(Idata[30]), .A2(n301), .ZN(n3) );
  OAI21_X1 U7 ( .B1(n303), .B2(n100), .A(n4), .ZN(n196) );
  NAND2_X1 U8 ( .A1(Idata[29]), .A2(n301), .ZN(n4) );
  OAI21_X1 U9 ( .B1(n303), .B2(n101), .A(n5), .ZN(n197) );
  NAND2_X1 U10 ( .A1(Idata[28]), .A2(n301), .ZN(n5) );
  OAI21_X1 U11 ( .B1(n303), .B2(n102), .A(n6), .ZN(n198) );
  NAND2_X1 U12 ( .A1(Idata[27]), .A2(n301), .ZN(n6) );
  OAI21_X1 U13 ( .B1(n302), .B2(n103), .A(n7), .ZN(n199) );
  NAND2_X1 U14 ( .A1(Idata[26]), .A2(n301), .ZN(n7) );
  OAI21_X1 U15 ( .B1(n303), .B2(n104), .A(n8), .ZN(n200) );
  NAND2_X1 U16 ( .A1(Idata[25]), .A2(n301), .ZN(n8) );
  OAI21_X1 U17 ( .B1(n302), .B2(n105), .A(n9), .ZN(n201) );
  NAND2_X1 U18 ( .A1(Idata[24]), .A2(n300), .ZN(n9) );
  OAI21_X1 U19 ( .B1(n302), .B2(n106), .A(n10), .ZN(n202) );
  NAND2_X1 U20 ( .A1(Idata[23]), .A2(n301), .ZN(n10) );
  OAI21_X1 U21 ( .B1(n302), .B2(n107), .A(n11), .ZN(n203) );
  NAND2_X1 U22 ( .A1(Idata[22]), .A2(n300), .ZN(n11) );
  OAI21_X1 U23 ( .B1(n301), .B2(n108), .A(n12), .ZN(n204) );
  NAND2_X1 U24 ( .A1(Idata[21]), .A2(n300), .ZN(n12) );
  OAI21_X1 U25 ( .B1(n301), .B2(n109), .A(n13), .ZN(n205) );
  NAND2_X1 U26 ( .A1(Idata[20]), .A2(n300), .ZN(n13) );
  OAI21_X1 U27 ( .B1(n302), .B2(n110), .A(n14), .ZN(n206) );
  NAND2_X1 U28 ( .A1(Idata[19]), .A2(n300), .ZN(n14) );
  OAI21_X1 U29 ( .B1(n301), .B2(n111), .A(n15), .ZN(n207) );
  NAND2_X1 U30 ( .A1(Idata[18]), .A2(n300), .ZN(n15) );
  OAI21_X1 U31 ( .B1(n301), .B2(n112), .A(n16), .ZN(n208) );
  NAND2_X1 U32 ( .A1(Idata[17]), .A2(n300), .ZN(n16) );
  OAI21_X1 U33 ( .B1(n302), .B2(n113), .A(n17), .ZN(n209) );
  NAND2_X1 U34 ( .A1(Idata[16]), .A2(n300), .ZN(n17) );
  OAI21_X1 U35 ( .B1(n302), .B2(n114), .A(n18), .ZN(n210) );
  NAND2_X1 U36 ( .A1(Idata[15]), .A2(n300), .ZN(n18) );
  OAI21_X1 U37 ( .B1(n302), .B2(n115), .A(n19), .ZN(n211) );
  NAND2_X1 U38 ( .A1(Idata[14]), .A2(n300), .ZN(n19) );
  OAI21_X1 U39 ( .B1(n302), .B2(n116), .A(n20), .ZN(n212) );
  NAND2_X1 U40 ( .A1(Idata[13]), .A2(n300), .ZN(n20) );
  OAI21_X1 U41 ( .B1(n302), .B2(n117), .A(n21), .ZN(n213) );
  NAND2_X1 U42 ( .A1(Idata[12]), .A2(n299), .ZN(n21) );
  OAI21_X1 U43 ( .B1(n302), .B2(n118), .A(n22), .ZN(n214) );
  NAND2_X1 U44 ( .A1(Idata[11]), .A2(n299), .ZN(n22) );
  OAI21_X1 U45 ( .B1(n303), .B2(n119), .A(n23), .ZN(n215) );
  NAND2_X1 U46 ( .A1(Idata[10]), .A2(n299), .ZN(n23) );
  OAI21_X1 U47 ( .B1(n302), .B2(n120), .A(n24), .ZN(n216) );
  NAND2_X1 U48 ( .A1(Idata[9]), .A2(n299), .ZN(n24) );
  OAI21_X1 U49 ( .B1(n303), .B2(n121), .A(n25), .ZN(n217) );
  NAND2_X1 U50 ( .A1(Idata[8]), .A2(n299), .ZN(n25) );
  OAI21_X1 U51 ( .B1(n303), .B2(n122), .A(n26), .ZN(n218) );
  NAND2_X1 U52 ( .A1(Idata[7]), .A2(n299), .ZN(n26) );
  OAI21_X1 U53 ( .B1(n303), .B2(n123), .A(n27), .ZN(n219) );
  NAND2_X1 U54 ( .A1(Idata[6]), .A2(n299), .ZN(n27) );
  OAI21_X1 U55 ( .B1(n303), .B2(n124), .A(n28), .ZN(n220) );
  NAND2_X1 U56 ( .A1(Idata[5]), .A2(n299), .ZN(n28) );
  OAI21_X1 U57 ( .B1(n303), .B2(n125), .A(n29), .ZN(n221) );
  NAND2_X1 U58 ( .A1(Idata[4]), .A2(n299), .ZN(n29) );
  OAI21_X1 U59 ( .B1(n303), .B2(n126), .A(n30), .ZN(n222) );
  NAND2_X1 U60 ( .A1(Idata[3]), .A2(n299), .ZN(n30) );
  OAI21_X1 U61 ( .B1(n303), .B2(n127), .A(n31), .ZN(n223) );
  NAND2_X1 U62 ( .A1(Idata[2]), .A2(n299), .ZN(n31) );
  OAI21_X1 U63 ( .B1(n304), .B2(n128), .A(n32), .ZN(n224) );
  NAND2_X1 U64 ( .A1(Idata[1]), .A2(n299), .ZN(n32) );
  OAI21_X1 U65 ( .B1(n304), .B2(n129), .A(n33), .ZN(n225) );
  NAND2_X1 U66 ( .A1(Idata[0]), .A2(n300), .ZN(n33) );
  OAI21_X1 U67 ( .B1(n310), .B2(n130), .A(n34), .ZN(n226) );
  NAND2_X1 U68 ( .A1(n296), .A2(n307), .ZN(n34) );
  OAI21_X1 U69 ( .B1(n310), .B2(n131), .A(n35), .ZN(n227) );
  NAND2_X1 U70 ( .A1(PC_next[30]), .A2(n307), .ZN(n35) );
  OAI21_X1 U71 ( .B1(n309), .B2(n132), .A(n36), .ZN(n228) );
  NAND2_X1 U72 ( .A1(PC_next[29]), .A2(n307), .ZN(n36) );
  OAI21_X1 U73 ( .B1(n309), .B2(n133), .A(n37), .ZN(n229) );
  NAND2_X1 U74 ( .A1(PC_next[28]), .A2(n307), .ZN(n37) );
  OAI21_X1 U75 ( .B1(n309), .B2(n134), .A(n38), .ZN(n230) );
  NAND2_X1 U76 ( .A1(PC_next[27]), .A2(n307), .ZN(n38) );
  OAI21_X1 U77 ( .B1(n308), .B2(n135), .A(n39), .ZN(n231) );
  NAND2_X1 U78 ( .A1(PC_next[26]), .A2(n307), .ZN(n39) );
  OAI21_X1 U79 ( .B1(n309), .B2(n136), .A(n40), .ZN(n232) );
  NAND2_X1 U80 ( .A1(PC_next[25]), .A2(n307), .ZN(n40) );
  OAI21_X1 U81 ( .B1(n308), .B2(n137), .A(n41), .ZN(n233) );
  NAND2_X1 U82 ( .A1(PC_next[24]), .A2(n306), .ZN(n41) );
  OAI21_X1 U83 ( .B1(n308), .B2(n138), .A(n42), .ZN(n234) );
  NAND2_X1 U84 ( .A1(PC_next[23]), .A2(n307), .ZN(n42) );
  OAI21_X1 U85 ( .B1(n308), .B2(n139), .A(n43), .ZN(n235) );
  NAND2_X1 U86 ( .A1(PC_next[22]), .A2(n306), .ZN(n43) );
  OAI21_X1 U87 ( .B1(n307), .B2(n140), .A(n44), .ZN(n236) );
  NAND2_X1 U88 ( .A1(PC_next[21]), .A2(n306), .ZN(n44) );
  OAI21_X1 U89 ( .B1(n307), .B2(n141), .A(n45), .ZN(n237) );
  NAND2_X1 U90 ( .A1(PC_next[20]), .A2(n306), .ZN(n45) );
  OAI21_X1 U91 ( .B1(n308), .B2(n142), .A(n46), .ZN(n238) );
  NAND2_X1 U92 ( .A1(PC_next[19]), .A2(n306), .ZN(n46) );
  OAI21_X1 U93 ( .B1(n307), .B2(n143), .A(n47), .ZN(n239) );
  NAND2_X1 U94 ( .A1(PC_next[18]), .A2(n306), .ZN(n47) );
  OAI21_X1 U95 ( .B1(n307), .B2(n144), .A(n48), .ZN(n240) );
  NAND2_X1 U96 ( .A1(PC_next[17]), .A2(n306), .ZN(n48) );
  OAI21_X1 U97 ( .B1(n308), .B2(n145), .A(n49), .ZN(n241) );
  NAND2_X1 U98 ( .A1(PC_next[16]), .A2(n306), .ZN(n49) );
  OAI21_X1 U99 ( .B1(n308), .B2(n146), .A(n50), .ZN(n242) );
  NAND2_X1 U100 ( .A1(PC_next[15]), .A2(n306), .ZN(n50) );
  OAI21_X1 U101 ( .B1(n308), .B2(n147), .A(n51), .ZN(n243) );
  NAND2_X1 U102 ( .A1(PC_next[14]), .A2(n306), .ZN(n51) );
  OAI21_X1 U103 ( .B1(n308), .B2(n148), .A(n52), .ZN(n244) );
  NAND2_X1 U104 ( .A1(PC_next[13]), .A2(n306), .ZN(n52) );
  OAI21_X1 U105 ( .B1(n308), .B2(n149), .A(n53), .ZN(n245) );
  NAND2_X1 U106 ( .A1(PC_next[12]), .A2(n305), .ZN(n53) );
  OAI21_X1 U107 ( .B1(n308), .B2(n150), .A(n54), .ZN(n246) );
  NAND2_X1 U108 ( .A1(PC_next[11]), .A2(n305), .ZN(n54) );
  OAI21_X1 U109 ( .B1(n309), .B2(n151), .A(n55), .ZN(n247) );
  NAND2_X1 U110 ( .A1(PC_next[10]), .A2(n305), .ZN(n55) );
  OAI21_X1 U111 ( .B1(n308), .B2(n152), .A(n56), .ZN(n248) );
  NAND2_X1 U112 ( .A1(PC_next[9]), .A2(n305), .ZN(n56) );
  OAI21_X1 U113 ( .B1(n309), .B2(n153), .A(n57), .ZN(n249) );
  NAND2_X1 U114 ( .A1(PC_next[8]), .A2(n305), .ZN(n57) );
  OAI21_X1 U115 ( .B1(n309), .B2(n154), .A(n58), .ZN(n250) );
  NAND2_X1 U116 ( .A1(PC_next[7]), .A2(n305), .ZN(n58) );
  OAI21_X1 U117 ( .B1(n309), .B2(n155), .A(n59), .ZN(n251) );
  NAND2_X1 U118 ( .A1(PC_next[6]), .A2(n305), .ZN(n59) );
  OAI21_X1 U119 ( .B1(n309), .B2(n156), .A(n60), .ZN(n252) );
  NAND2_X1 U120 ( .A1(PC_next[5]), .A2(n305), .ZN(n60) );
  OAI21_X1 U121 ( .B1(n309), .B2(n157), .A(n61), .ZN(n253) );
  NAND2_X1 U122 ( .A1(PC_next[4]), .A2(n305), .ZN(n61) );
  OAI21_X1 U123 ( .B1(n309), .B2(n158), .A(n62), .ZN(n254) );
  NAND2_X1 U124 ( .A1(PC_next[3]), .A2(n305), .ZN(n62) );
  OAI21_X1 U125 ( .B1(n309), .B2(n159), .A(n63), .ZN(n255) );
  NAND2_X1 U126 ( .A1(PC_next[2]), .A2(n305), .ZN(n63) );
  OAI21_X1 U127 ( .B1(n310), .B2(n160), .A(n64), .ZN(n256) );
  NAND2_X1 U128 ( .A1(PC_next[1]), .A2(n305), .ZN(n64) );
  OAI21_X1 U129 ( .B1(PC_LATCH_EN_i), .B2(n161), .A(n65), .ZN(n257) );
  NAND2_X1 U130 ( .A1(PC_LATCH_EN_i), .A2(PC_BUS[30]), .ZN(n65) );
  OAI21_X1 U131 ( .B1(PC_LATCH_EN_i), .B2(n162), .A(n66), .ZN(n258) );
  NAND2_X1 U132 ( .A1(PC_BUS[29]), .A2(PC_LATCH_EN_i), .ZN(n66) );
  OAI21_X1 U133 ( .B1(PC_LATCH_EN_i), .B2(n163), .A(n67), .ZN(n259) );
  NAND2_X1 U134 ( .A1(PC_BUS[28]), .A2(PC_LATCH_EN_i), .ZN(n67) );
  OAI21_X1 U135 ( .B1(PC_LATCH_EN_i), .B2(n164), .A(n68), .ZN(n260) );
  NAND2_X1 U136 ( .A1(PC_BUS[27]), .A2(PC_LATCH_EN_i), .ZN(n68) );
  OAI21_X1 U137 ( .B1(PC_LATCH_EN_i), .B2(n165), .A(n69), .ZN(n261) );
  NAND2_X1 U138 ( .A1(PC_BUS[26]), .A2(PC_LATCH_EN_i), .ZN(n69) );
  OAI21_X1 U139 ( .B1(PC_LATCH_EN_i), .B2(n166), .A(n70), .ZN(n262) );
  NAND2_X1 U140 ( .A1(PC_BUS[25]), .A2(PC_LATCH_EN_i), .ZN(n70) );
  OAI21_X1 U141 ( .B1(PC_LATCH_EN_i), .B2(n167), .A(n71), .ZN(n263) );
  NAND2_X1 U142 ( .A1(PC_BUS[24]), .A2(PC_LATCH_EN_i), .ZN(n71) );
  OAI21_X1 U143 ( .B1(PC_LATCH_EN_i), .B2(n168), .A(n72), .ZN(n264) );
  NAND2_X1 U144 ( .A1(PC_BUS[23]), .A2(PC_LATCH_EN_i), .ZN(n72) );
  OAI21_X1 U145 ( .B1(PC_LATCH_EN_i), .B2(n169), .A(n73), .ZN(n265) );
  NAND2_X1 U146 ( .A1(PC_BUS[22]), .A2(PC_LATCH_EN_i), .ZN(n73) );
  OAI21_X1 U147 ( .B1(PC_LATCH_EN_i), .B2(n170), .A(n74), .ZN(n266) );
  NAND2_X1 U148 ( .A1(PC_BUS[21]), .A2(PC_LATCH_EN_i), .ZN(n74) );
  OAI21_X1 U149 ( .B1(PC_LATCH_EN_i), .B2(n171), .A(n75), .ZN(n267) );
  NAND2_X1 U150 ( .A1(PC_BUS[20]), .A2(PC_LATCH_EN_i), .ZN(n75) );
  OAI21_X1 U151 ( .B1(PC_LATCH_EN_i), .B2(n172), .A(n76), .ZN(n268) );
  NAND2_X1 U152 ( .A1(PC_BUS[19]), .A2(PC_LATCH_EN_i), .ZN(n76) );
  OAI21_X1 U153 ( .B1(PC_LATCH_EN_i), .B2(n173), .A(n77), .ZN(n269) );
  NAND2_X1 U154 ( .A1(PC_BUS[18]), .A2(PC_LATCH_EN_i), .ZN(n77) );
  OAI21_X1 U155 ( .B1(PC_LATCH_EN_i), .B2(n174), .A(n78), .ZN(n270) );
  NAND2_X1 U156 ( .A1(PC_BUS[17]), .A2(PC_LATCH_EN_i), .ZN(n78) );
  OAI21_X1 U157 ( .B1(PC_LATCH_EN_i), .B2(n175), .A(n79), .ZN(n271) );
  NAND2_X1 U158 ( .A1(PC_BUS[16]), .A2(PC_LATCH_EN_i), .ZN(n79) );
  OAI21_X1 U159 ( .B1(PC_LATCH_EN_i), .B2(n176), .A(n80), .ZN(n272) );
  NAND2_X1 U160 ( .A1(PC_BUS[15]), .A2(PC_LATCH_EN_i), .ZN(n80) );
  OAI21_X1 U161 ( .B1(PC_LATCH_EN_i), .B2(n177), .A(n81), .ZN(n273) );
  NAND2_X1 U162 ( .A1(PC_BUS[14]), .A2(PC_LATCH_EN_i), .ZN(n81) );
  OAI21_X1 U163 ( .B1(PC_LATCH_EN_i), .B2(n178), .A(n82), .ZN(n274) );
  NAND2_X1 U164 ( .A1(PC_BUS[13]), .A2(PC_LATCH_EN_i), .ZN(n82) );
  OAI21_X1 U165 ( .B1(PC_LATCH_EN_i), .B2(n179), .A(n83), .ZN(n275) );
  NAND2_X1 U166 ( .A1(PC_BUS[12]), .A2(PC_LATCH_EN_i), .ZN(n83) );
  OAI21_X1 U167 ( .B1(PC_LATCH_EN_i), .B2(n180), .A(n84), .ZN(n276) );
  NAND2_X1 U168 ( .A1(PC_BUS[11]), .A2(PC_LATCH_EN_i), .ZN(n84) );
  OAI21_X1 U169 ( .B1(PC_LATCH_EN_i), .B2(n181), .A(n85), .ZN(n277) );
  NAND2_X1 U170 ( .A1(PC_BUS[10]), .A2(PC_LATCH_EN_i), .ZN(n85) );
  OAI21_X1 U171 ( .B1(PC_LATCH_EN_i), .B2(n182), .A(n86), .ZN(n278) );
  NAND2_X1 U172 ( .A1(PC_BUS[9]), .A2(PC_LATCH_EN_i), .ZN(n86) );
  OAI21_X1 U173 ( .B1(PC_LATCH_EN_i), .B2(n183), .A(n87), .ZN(n279) );
  NAND2_X1 U174 ( .A1(PC_BUS[8]), .A2(PC_LATCH_EN_i), .ZN(n87) );
  OAI21_X1 U175 ( .B1(PC_LATCH_EN_i), .B2(n184), .A(n88), .ZN(n280) );
  NAND2_X1 U176 ( .A1(PC_BUS[7]), .A2(PC_LATCH_EN_i), .ZN(n88) );
  OAI21_X1 U177 ( .B1(PC_LATCH_EN_i), .B2(n185), .A(n89), .ZN(n281) );
  NAND2_X1 U178 ( .A1(PC_BUS[6]), .A2(PC_LATCH_EN_i), .ZN(n89) );
  OAI21_X1 U179 ( .B1(PC_LATCH_EN_i), .B2(n186), .A(n90), .ZN(n282) );
  NAND2_X1 U180 ( .A1(PC_BUS[5]), .A2(PC_LATCH_EN_i), .ZN(n90) );
  OAI21_X1 U181 ( .B1(PC_LATCH_EN_i), .B2(n187), .A(n91), .ZN(n283) );
  NAND2_X1 U182 ( .A1(PC_BUS[4]), .A2(PC_LATCH_EN_i), .ZN(n91) );
  OAI21_X1 U183 ( .B1(PC_LATCH_EN_i), .B2(n188), .A(n92), .ZN(n284) );
  NAND2_X1 U184 ( .A1(PC_BUS[3]), .A2(PC_LATCH_EN_i), .ZN(n92) );
  OAI21_X1 U185 ( .B1(PC_LATCH_EN_i), .B2(n189), .A(n93), .ZN(n285) );
  NAND2_X1 U186 ( .A1(PC_BUS[2]), .A2(PC_LATCH_EN_i), .ZN(n93) );
  OAI21_X1 U187 ( .B1(PC_LATCH_EN_i), .B2(n190), .A(n94), .ZN(n286) );
  NAND2_X1 U188 ( .A1(PC_BUS[1]), .A2(PC_LATCH_EN_i), .ZN(n94) );
  OAI21_X1 U189 ( .B1(PC_LATCH_EN_i), .B2(n191), .A(n95), .ZN(n287) );
  NAND2_X1 U190 ( .A1(PC_BUS[0]), .A2(PC_LATCH_EN_i), .ZN(n95) );
  NAND2_X1 U192 ( .A1(PC_BUS[31]), .A2(PC_LATCH_EN_i), .ZN(n96) );
  OAI21_X1 U193 ( .B1(n310), .B2(n193), .A(n97), .ZN(n289) );
  NAND2_X1 U194 ( .A1(PC_next[0]), .A2(n306), .ZN(n97) );
  INV_X1 U195 ( .A(n290), .ZN(RD[4]) );
  AOI22_X1 U196 ( .A1(IMM26[20]), .A2(n291), .B1(N2), .B2(INP2[15]), .ZN(n290)
         );
  INV_X1 U197 ( .A(n292), .ZN(RD[3]) );
  AOI22_X1 U198 ( .A1(IMM26[19]), .A2(n291), .B1(INP2[14]), .B2(N2), .ZN(n292)
         );
  INV_X1 U199 ( .A(n293), .ZN(RD[2]) );
  AOI22_X1 U200 ( .A1(IMM26[18]), .A2(n291), .B1(INP2[13]), .B2(N2), .ZN(n293)
         );
  INV_X1 U201 ( .A(n294), .ZN(RD[1]) );
  AOI22_X1 U202 ( .A1(IMM26[17]), .A2(n291), .B1(INP2[12]), .B2(N2), .ZN(n294)
         );
  INV_X1 U203 ( .A(n295), .ZN(RD[0]) );
  AOI22_X1 U204 ( .A1(IMM26[16]), .A2(n291), .B1(INP2[11]), .B2(N2), .ZN(n295)
         );
  INV_X1 U205 ( .A(N2), .ZN(n291) );
  NPC_logic_PC_SIZE32 NPC_logic_0 ( .Flush_BTB(Flush_BTB), .BRANCH_CTRL_SIG(
        BRANCH_CTRL_SIG), .OUTT_NT_i(OUTT_NT_i), .PC_next(PC_next), 
        .BRANCH_ALU_OUT(BRANCH_ALU_OUT), .OUT_PC_target_i(OUT_PC_target_i), 
        .NPC(NPC), .PC_BUS(PC_BUS) );
  dlx_cu_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE29 CU_I ( .Clk(Clk), .Rst(
        n311), .Flush_BTB(Flush_BTB_i), .STALL(STALL_i), .IR_IN({IR, IMM26, 
        INP2}), .IR_LATCH_EN(IR_LATCH_EN_i), .NPC_LATCH_EN(NPC_LATCH_EN_i), 
        .I_R_type(I_R_TYPE_i), .REGF_LATCH_EN(RegRF_LATCH_EN_i), 
        .RegA_LATCH_EN(RegA_LATCH_EN_i), .RegB_LATCH_EN(RegB_LATCH_EN_i), 
        .RegIMM_LATCH_EN(RegIMM_LATCH_EN_i), .RegRD1_LATCH_EN(
        RegRD1_LATCH_EN_i), .SIGN_UNSIGN(SIGN_UNSIGN_i), .RFR1_EN(RFR1_EN_i), 
        .RFR2_EN(RFR2_EN_i), .MUX_IMM_SEL(MUX_IMM_SEL_i), .JUMP(JUMP_i), 
        .JUMP_EN(JUMP_EN_i), .EQ_COND(EQ_COND_i), .MUXA_SEL(MUXA_SEL_i), 
        .MUXB_SEL(MUXB_SEL_i), .ALU_OUTREG_EN(ALU_OUTREG_EN_i), 
        .REGME_LATCH_EN(REGME_LATCH_EN_i), .RegRD2_LATCH_EN(RegRD2_LATCH_EN_i), 
        .ALU_OPCODE(ALU_OPCODE_i), .DRAM_EN(Denable), .DRAM_RE(Drd), .DRAM_WE(
        Dwd), .LMD_LATCH_EN(LMD_LATCH_EN_i), .RALUOUT2_LATCH_EN(
        RALUOUT2_LATCH_EN_i), .RegRD3_LATCH_EN(RegRD3_LATCH_EN_i), 
        .PC_LATCH_EN(PC_LATCH_EN_i), .RPCplus8_LATCH_EN(RPCplus8_LATCH_EN_i), 
        .WB_MUX_SEL(WB_MUX_SEL_i), .RF_WE(RF_WE_i), .JandL(JandL_i), 
        .REGWRITE_DX(REGWRITE_DX_i), .REGWRITE_XM(REGWRITE_XM_i), 
        .REGWRITE_MW(REGWRITE_MW_i), .MEMREAD_DX(MEMREAD_DX_i) );
  datapath_NUMBIT32_ADDRESS_WIDTH_RF5_ADDRESS_WIDTH_DM32 DP_I ( .CLK(Clk), 
        .RST(n311), .INP1(NPC), .INP2(INP2), .IMM26({IMM26, INP2}), .RS1(
        IMM26[25:21]), .RS2(IMM26[20:16]), .RD(RD), .REGF_LATCH_EN(
        RegRF_LATCH_EN_i), .RegA_LATCH_EN(RegA_LATCH_EN_i), .RegB_LATCH_EN(
        RegB_LATCH_EN_i), .RegIMM_LATCH_EN(RegIMM_LATCH_EN_i), 
        .RegRD1_LATCH_EN(RegRD1_LATCH_EN_i), .SIGN_UNSIGN(SIGN_UNSIGN_i), 
        .RFR1_EN(RFR1_EN_i), .RFR2_EN(RFR2_EN_i), .MUX_IMM_SEL(MUX_IMM_SEL_i), 
        .JUMP(JUMP_i), .JUMP_EN(JUMP_EN_i), .EQ_COND(EQ_COND_i), .MUXA_SEL(
        MUXA_SEL_i), .MUXB_SEL(MUXB_SEL_i), .RALUOUT_LATCH_EN(ALU_OUTREG_EN_i), 
        .REGME_LATCH_EN(REGME_LATCH_EN_i), .RegRD2_LATCH_EN(RegRD2_LATCH_EN_i), 
        .ALU_OPCODE(ALU_OPCODE_i), .ADDR_DRAM(Daddr), .DATAIN_DRAM(Ddatain), 
        .DATAOUT_DRAM(Ddataout), .LMD_LATCH_EN(LMD_LATCH_EN_i), 
        .RALUOUT2_LATCH_EN(RALUOUT2_LATCH_EN_i), .RegRD3_LATCH_EN(
        RegRD3_LATCH_EN_i), .RPCplus8_LATCH_EN(RPCplus8_LATCH_EN_i), 
        .WB_MUX_SEL(WB_MUX_SEL_i), .RF_WE(RF_WE_i), .ROUT_LATCH_EN(1'b0), 
        .JandL(JandL_i), .BRANCH_CTRL_SIG(BRANCH_CTRL_SIG), .BRANCH_ALU_OUT(
        BRANCH_ALU_OUT), .Data_out(DataOut), .REGWRITE_XM(REGWRITE_XM_i), 
        .REGWRITE_MW(REGWRITE_MW_i) );
  BTB_PC_SIZE32_BTBSIZE5 BTB_0 ( .Reset(n311), .Clk(Clk), .Enable(1'b1), 
        .PC_read({n296, PC_next[30:0]}), .WR(JUMP_EN_i), .PC_write(NPC), 
        .SetT_NT(BRANCH_CTRL_SIG), .Set_target(BRANCH_ALU_OUT), 
        .OUT_PC_target(OUT_PC_target_i), .OUTT_NT(OUTT_NT_i), .prevT_NT(
        prevT_NT_i) );
  HazardUnit_NUMBIT32_ADDRESS_WIDTH_RF5_OP_CODE_SIZE6 HU_0 ( .CLK(Clk), .RST(
        n311), .RS1(IMM26[25:21]), .RS2(IMM26[20:16]), .REGWRITE_DX(
        REGWRITE_DX_i), .MEMREAD_DX(MEMREAD_DX_i), .RD(IMM26[20:16]), .OPCODE(
        IR), .STALL(STALL_i) );
  DLX_IR_SIZE32_PC_SIZE32_DW01_inc_1 add_365 ( .A({Iaddr[31:1], n314}), .SUM(
        PC_next) );
  DFFR_X1 \PC_reg[31]  ( .D(n288), .CK(Clk), .RN(n311), .Q(Iaddr[31]), .QN(
        n192) );
  BUF_X8 U206 ( .A(Rst), .Z(n311) );
  CLKBUF_X1 U207 ( .A(PC_next[31]), .Z(n296) );
  INV_X1 U208 ( .A(n191), .ZN(Iaddr[0]) );
  OR2_X1 U209 ( .A1(PC_LATCH_EN_i), .A2(n192), .ZN(n298) );
  NAND2_X1 U210 ( .A1(n298), .A2(n96), .ZN(n288) );
  CLKBUF_X1 U211 ( .A(IR_LATCH_EN_i), .Z(n299) );
  CLKBUF_X1 U212 ( .A(IR_LATCH_EN_i), .Z(n300) );
  CLKBUF_X1 U213 ( .A(IR_LATCH_EN_i), .Z(n301) );
  CLKBUF_X1 U214 ( .A(IR_LATCH_EN_i), .Z(n302) );
  CLKBUF_X1 U215 ( .A(IR_LATCH_EN_i), .Z(n303) );
  CLKBUF_X1 U216 ( .A(IR_LATCH_EN_i), .Z(n304) );
  CLKBUF_X1 U217 ( .A(NPC_LATCH_EN_i), .Z(n305) );
  CLKBUF_X1 U218 ( .A(NPC_LATCH_EN_i), .Z(n306) );
  CLKBUF_X1 U219 ( .A(NPC_LATCH_EN_i), .Z(n307) );
  CLKBUF_X1 U220 ( .A(NPC_LATCH_EN_i), .Z(n308) );
  CLKBUF_X1 U221 ( .A(NPC_LATCH_EN_i), .Z(n309) );
  CLKBUF_X1 U222 ( .A(NPC_LATCH_EN_i), .Z(n310) );
  CLKBUF_X3 U223 ( .A(Rst), .Z(n312) );
  CLKBUF_X3 U224 ( .A(Rst), .Z(n313) );
endmodule

