library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

entity FP_ALU is
  port (
  clock
  );
end entity;

architecture arch of FP_ALU is

begin

end architecture;
