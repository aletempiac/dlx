
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX_IR_SIZE32_PC_SIZE32 is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type VHDLOUT_TYPE is range 0 to 2;
type VHDLOUT_TYPE_2 is range 0 to 5;
type aluOp is (ADDS, SUBS, ANDS, ORS, XORS, SLLS, SRLS, SRAS, SEQS, SNES, SLTS,
   SGTS, SLES, SGES, SLTUS, SGTUS, SLEUS, SGEUS, NOP);
attribute ENUM_ENCODING of aluOp : type is 
   "00000 00001 00010 00011 00100 00101 00110 00111 01000 01001 01010 01011 01100 01101 01110 01111 10000 10001 10010";
   
   -- Declarations for conversion functions.
   function integer_to_unsigned(arg, size : in INTEGER) return std_logic_vector
               ;
   function std_logic_vector_to_aluOp(arg : in std_logic_vector( 1 to 5 )) 
               return aluOp;
   function aluOp_to_std_logic_vector(arg : in aluOp) return std_logic_vector;

end CONV_PACK_DLX_IR_SIZE32_PC_SIZE32;

package body CONV_PACK_DLX_IR_SIZE32_PC_SIZE32 is
   
   -- integer type to std_logic_vector function
   function integer_to_unsigned(arg, size : in INTEGER) return std_logic_vector
   is 
      variable result: std_logic_vector(size-1 downto 0);
      variable temp: INTEGER;
      -- synopsys built_in SYN_INTEGER_TO_UNSIGNED
   begin
      temp := arg;
      for i in 0 to size-1 loop
         if (temp mod 2) = 1 then
            result(i) := '1';
         else
            result(i) := '0';
         end if;
         temp := temp / 2;
      end loop;
      return result;
   end;
   
   -- std_logic_vector to enum type function
   function std_logic_vector_to_aluOp(arg : in std_logic_vector( 1 to 5 )) 
   return aluOp is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when "00000" => return ADDS;
         when "00001" => return SUBS;
         when "00010" => return ANDS;
         when "00011" => return ORS;
         when "00100" => return XORS;
         when "00101" => return SLLS;
         when "00110" => return SRLS;
         when "00111" => return SRAS;
         when "01000" => return SEQS;
         when "01001" => return SNES;
         when "01010" => return SLTS;
         when "01011" => return SGTS;
         when "01100" => return SLES;
         when "01101" => return SGES;
         when "01110" => return SLTUS;
         when "01111" => return SGTUS;
         when "10000" => return SLEUS;
         when "10001" => return SGEUS;
         when "10010" => return NOP;
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return ADDS;
      end case;
   end;
   
   -- enum type to std_logic_vector function
   function aluOp_to_std_logic_vector(arg : in aluOp) return std_logic_vector 
   is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when ADDS => return "00000";
         when SUBS => return "00001";
         when ANDS => return "00010";
         when ORS => return "00011";
         when XORS => return "00100";
         when SLLS => return "00101";
         when SRLS => return "00110";
         when SRAS => return "00111";
         when SEQS => return "01000";
         when SNES => return "01001";
         when SLTS => return "01010";
         when SGTS => return "01011";
         when SLES => return "01100";
         when SGES => return "01101";
         when SLTUS => return "01110";
         when SGTUS => return "01111";
         when SLEUS => return "10000";
         when SGEUS => return "10001";
         when NOP => return "10010";
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return "00000";
      end case;
   end;

end CONV_PACK_DLX_IR_SIZE32_PC_SIZE32;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity DLX_IR_SIZE32_PC_SIZE32_DW01_inc_1 is

   port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector (31
         downto 0));

end DLX_IR_SIZE32_PC_SIZE32_DW01_inc_1;

architecture SYN_cla of DLX_IR_SIZE32_PC_SIZE32_DW01_inc_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X2
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106 : std_logic;

begin
   
   U2 : XNOR2_X2 port map( A => A(4), B => n54, ZN => SUM(4));
   U3 : INV_X1 port map( A => n32, ZN => n54);
   U4 : NOR2_X1 port map( A1 => n72, A2 => n24, ZN => n1);
   U5 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => n66);
   U6 : AND2_X1 port map( A1 => n3, A2 => A(26), ZN => n2);
   U7 : INV_X1 port map( A => n25, ZN => n3);
   U8 : OR2_X1 port map( A1 => n24, A2 => n72, ZN => n4);
   U9 : OR2_X1 port map( A1 => n20, A2 => n21, ZN => n5);
   U10 : OR2_X2 port map( A1 => n5, A2 => n6, ZN => n85);
   U11 : OR2_X1 port map( A1 => n7, A2 => n39, ZN => n6);
   U12 : INV_X1 port map( A => A(18), ZN => n7);
   U13 : INV_X1 port map( A => A(25), ZN => n24);
   U14 : NOR2_X1 port map( A1 => n24, A2 => n72, ZN => n23);
   U15 : NOR2_X1 port map( A1 => n59, A2 => n60, ZN => n57);
   U16 : XNOR2_X1 port map( A => n57, B => n58, ZN => SUM(31));
   U17 : OR2_X2 port map( A1 => n20, A2 => n21, ZN => n89);
   U18 : NOR2_X2 port map( A1 => n43, A2 => n101, ZN => n42);
   U19 : OR2_X2 port map( A1 => n8, A2 => n9, ZN => n101);
   U20 : NOR2_X2 port map( A1 => n41, A2 => n85, ZN => n40);
   U21 : NAND2_X1 port map( A1 => n30, A2 => A(8), ZN => n8);
   U22 : OR2_X1 port map( A1 => n10, A2 => n36, ZN => n9);
   U23 : INV_X1 port map( A => A(10), ZN => n10);
   U24 : NAND2_X1 port map( A1 => n40, A2 => A(20), ZN => n11);
   U25 : OR2_X1 port map( A1 => n11, A2 => n12, ZN => n76);
   U26 : OR2_X1 port map( A1 => n13, A2 => n34, ZN => n12);
   U27 : INV_X1 port map( A => A(22), ZN => n13);
   U28 : OR2_X1 port map( A1 => n11, A2 => n12, ZN => n14);
   U29 : OR2_X2 port map( A1 => n14, A2 => n15, ZN => n72);
   U30 : OR2_X1 port map( A1 => n16, A2 => n29, ZN => n15);
   U31 : INV_X1 port map( A => A(24), ZN => n16);
   U32 : NAND2_X1 port map( A1 => n42, A2 => A(12), ZN => n17);
   U33 : OR2_X1 port map( A1 => n17, A2 => n18, ZN => n93);
   U34 : OR2_X1 port map( A1 => n19, A2 => n27, ZN => n18);
   U35 : INV_X1 port map( A => A(14), ZN => n19);
   U36 : OR2_X1 port map( A1 => n17, A2 => n18, ZN => n20);
   U37 : OR2_X1 port map( A1 => n22, A2 => n45, ZN => n21);
   U38 : INV_X1 port map( A => A(16), ZN => n22);
   U39 : NOR2_X1 port map( A1 => n103, A2 => n36, ZN => n35);
   U40 : INV_X32 port map( A => A(27), ZN => n25);
   U41 : INV_X1 port map( A => n26, ZN => n94);
   U42 : NOR2_X1 port map( A1 => n27, A2 => n97, ZN => n26);
   U43 : INV_X32 port map( A => A(13), ZN => n27);
   U44 : INV_X1 port map( A => n28, ZN => n73);
   U45 : NOR2_X1 port map( A1 => n29, A2 => n76, ZN => n28);
   U46 : INV_X1 port map( A => n35, ZN => n102);
   U47 : INV_X1 port map( A => A(11), ZN => n43);
   U48 : INV_X32 port map( A => A(23), ZN => n29);
   U49 : AND2_X1 port map( A1 => A(1), A2 => A(0), ZN => n37);
   U50 : INV_X1 port map( A => n37, ZN => n62);
   U51 : INV_X2 port map( A => n30, ZN => n48);
   U52 : INV_X2 port map( A => n31, ZN => n51);
   U53 : NAND2_X1 port map( A1 => A(6), A2 => n31, ZN => n104);
   U54 : NAND2_X1 port map( A1 => A(4), A2 => n32, ZN => n105);
   U55 : AND2_X2 port map( A1 => A(7), A2 => n49, ZN => n30);
   U56 : AND2_X2 port map( A1 => A(5), A2 => n52, ZN => n31);
   U57 : NOR2_X1 port map( A1 => n34, A2 => n80, ZN => n33);
   U58 : INV_X1 port map( A => A(9), ZN => n36);
   U59 : INV_X1 port map( A => n33, ZN => n77);
   U60 : AND2_X2 port map( A1 => A(3), A2 => n55, ZN => n32);
   U61 : INV_X32 port map( A => A(21), ZN => n34);
   U62 : NOR2_X1 port map( A1 => n39, A2 => n89, ZN => n38);
   U63 : INV_X1 port map( A => n38, ZN => n86);
   U64 : INV_X32 port map( A => A(17), ZN => n39);
   U65 : INV_X1 port map( A => n42, ZN => n98);
   U66 : INV_X1 port map( A => n40, ZN => n81);
   U67 : INV_X32 port map( A => A(19), ZN => n41);
   U68 : NOR2_X1 port map( A1 => n45, A2 => n93, ZN => n44);
   U69 : INV_X1 port map( A => n44, ZN => n90);
   U70 : INV_X32 port map( A => A(15), ZN => n45);
   U71 : NAND2_X1 port map( A1 => A(8), A2 => n30, ZN => n103);
   U72 : NAND2_X1 port map( A1 => A(28), A2 => n65, ZN => n64);
   U73 : XNOR2_X1 port map( A => A(6), B => n51, ZN => SUM(6));
   U74 : XNOR2_X1 port map( A => A(2), B => n62, ZN => SUM(2));
   U75 : XNOR2_X1 port map( A => A(26), B => n4, ZN => SUM(26));
   U76 : XNOR2_X1 port map( A => A(16), B => n90, ZN => SUM(16));
   U77 : XNOR2_X1 port map( A => A(22), B => n77, ZN => SUM(22));
   U78 : XNOR2_X1 port map( A => A(12), B => n98, ZN => SUM(12));
   U79 : INV_X1 port map( A => A(0), ZN => SUM(0));
   U80 : XNOR2_X1 port map( A => A(10), B => n102, ZN => SUM(10));
   U81 : XNOR2_X1 port map( A => A(8), B => n48, ZN => SUM(8));
   U82 : XNOR2_X1 port map( A => A(20), B => n81, ZN => SUM(20));
   U83 : XNOR2_X1 port map( A => A(18), B => n86, ZN => SUM(18));
   U84 : XNOR2_X1 port map( A => A(28), B => n66, ZN => SUM(28));
   U85 : XNOR2_X1 port map( A => A(0), B => n83, ZN => SUM(1));
   U86 : XNOR2_X1 port map( A => A(24), B => n73, ZN => SUM(24));
   U87 : XNOR2_X1 port map( A => A(14), B => n94, ZN => SUM(14));
   U88 : NAND2_X1 port map( A1 => A(29), A2 => n61, ZN => n59);
   U89 : NAND2_X1 port map( A1 => A(26), A2 => n23, ZN => n69);
   U90 : NAND2_X1 port map( A1 => A(20), A2 => n40, ZN => n80);
   U91 : NAND2_X1 port map( A1 => A(12), A2 => n42, ZN => n97);
   U92 : NAND2_X1 port map( A1 => A(2), A2 => n37, ZN => n106);
   U93 : XNOR2_X1 port map( A => n46, B => n47, ZN => SUM(9));
   U94 : INV_X2 port map( A => A(9), ZN => n47);
   U95 : XNOR2_X1 port map( A => n49, B => n50, ZN => SUM(7));
   U96 : INV_X2 port map( A => A(7), ZN => n50);
   U97 : XNOR2_X1 port map( A => n52, B => n53, ZN => SUM(5));
   U98 : INV_X2 port map( A => A(5), ZN => n53);
   U99 : XNOR2_X1 port map( A => n55, B => n56, ZN => SUM(3));
   U100 : INV_X2 port map( A => A(3), ZN => n56);
   U101 : INV_X2 port map( A => A(31), ZN => n58);
   U102 : INV_X2 port map( A => A(30), ZN => n60);
   U103 : XNOR2_X2 port map( A => A(30), B => n59, ZN => SUM(30));
   U104 : XNOR2_X1 port map( A => n61, B => n63, ZN => SUM(29));
   U105 : INV_X2 port map( A => A(29), ZN => n63);
   U106 : INV_X1 port map( A => n64, ZN => n61);
   U107 : INV_X1 port map( A => n66, ZN => n65);
   U108 : XNOR2_X1 port map( A => n67, B => n68, ZN => SUM(27));
   U109 : INV_X2 port map( A => A(27), ZN => n68);
   U110 : INV_X1 port map( A => n69, ZN => n67);
   U111 : XNOR2_X1 port map( A => n70, B => n71, ZN => SUM(25));
   U112 : INV_X2 port map( A => A(25), ZN => n71);
   U113 : INV_X1 port map( A => n72, ZN => n70);
   U114 : XNOR2_X1 port map( A => n74, B => n75, ZN => SUM(23));
   U115 : INV_X2 port map( A => A(23), ZN => n75);
   U116 : INV_X1 port map( A => n76, ZN => n74);
   U117 : XNOR2_X1 port map( A => n78, B => n79, ZN => SUM(21));
   U118 : INV_X2 port map( A => A(21), ZN => n79);
   U119 : INV_X1 port map( A => n80, ZN => n78);
   U120 : INV_X2 port map( A => A(1), ZN => n83);
   U121 : XNOR2_X1 port map( A => n82, B => n84, ZN => SUM(19));
   U122 : INV_X2 port map( A => A(19), ZN => n84);
   U123 : INV_X1 port map( A => n85, ZN => n82);
   U124 : XNOR2_X1 port map( A => n87, B => n88, ZN => SUM(17));
   U125 : INV_X2 port map( A => A(17), ZN => n88);
   U126 : INV_X1 port map( A => n89, ZN => n87);
   U127 : XNOR2_X1 port map( A => n91, B => n92, ZN => SUM(15));
   U128 : INV_X2 port map( A => A(15), ZN => n92);
   U129 : INV_X1 port map( A => n93, ZN => n91);
   U130 : XNOR2_X1 port map( A => n95, B => n96, ZN => SUM(13));
   U131 : INV_X2 port map( A => A(13), ZN => n96);
   U132 : INV_X1 port map( A => n97, ZN => n95);
   U133 : XNOR2_X1 port map( A => n99, B => n100, ZN => SUM(11));
   U134 : INV_X2 port map( A => A(11), ZN => n100);
   U135 : INV_X1 port map( A => n101, ZN => n99);
   U136 : INV_X1 port map( A => n103, ZN => n46);
   U137 : INV_X1 port map( A => n104, ZN => n49);
   U138 : INV_X1 port map( A => n105, ZN => n52);
   U139 : INV_X1 port map( A => n106, ZN => n55);

end SYN_cla;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_1 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1;

architecture SYN_BEHAVIORAL of FA_1 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U2 : INV_X1 port map( A => n11, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n10, B2 => Ci, ZN => n11);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_2 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2;

architecture SYN_BEHAVIORAL of FA_2 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U2 : INV_X1 port map( A => n12, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_3 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_3;

architecture SYN_BEHAVIORAL of FA_3 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_4 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_4;

architecture SYN_BEHAVIORAL of FA_4 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8, n9, n10 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => n8, B => Ci, Z => S);
   U2 : INV_X1 port map( A => n9, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => n10, B1 => n8, B2 => Ci, ZN => n9);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n8);
   U5 : CLKBUF_X1 port map( A => A, Z => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_5 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_5;

architecture SYN_BEHAVIORAL of FA_5 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_6 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_6;

architecture SYN_BEHAVIORAL of FA_6 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U2 : INV_X1 port map( A => n12, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_7 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_7;

architecture SYN_BEHAVIORAL of FA_7 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_8 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_8;

architecture SYN_BEHAVIORAL of FA_8 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => n8, B => Ci, Z => S);
   U2 : INV_X1 port map( A => n9, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n8, B2 => Ci, ZN => n9);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_9 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_9;

architecture SYN_BEHAVIORAL of FA_9 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U2 : INV_X1 port map( A => n13, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n13);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_10 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_10;

architecture SYN_BEHAVIORAL of FA_10 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U2 : INV_X1 port map( A => n13, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n13);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_11 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_11;

architecture SYN_BEHAVIORAL of FA_11 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_12 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_12;

architecture SYN_BEHAVIORAL of FA_12 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n10, n11 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U2 : INV_X1 port map( A => n11, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n10, B2 => Ci, ZN => n11);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_13 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_13;

architecture SYN_BEHAVIORAL of FA_13 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U2 : INV_X1 port map( A => n13, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n13);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_14 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_14;

architecture SYN_BEHAVIORAL of FA_14 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U2 : INV_X1 port map( A => n13, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n13);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_15 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_15;

architecture SYN_BEHAVIORAL of FA_15 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_16 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_16;

architecture SYN_BEHAVIORAL of FA_16 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U2 : INV_X1 port map( A => n10, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n10);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_17 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_17;

architecture SYN_BEHAVIORAL of FA_17 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U2 : INV_X1 port map( A => n13, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n13);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_18 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_18;

architecture SYN_BEHAVIORAL of FA_18 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_19 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_19;

architecture SYN_BEHAVIORAL of FA_19 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_20 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_20;

architecture SYN_BEHAVIORAL of FA_20 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U2 : INV_X1 port map( A => n10, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n10);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_21 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_21;

architecture SYN_BEHAVIORAL of FA_21 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U2 : INV_X1 port map( A => n13, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n13);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_22 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_22;

architecture SYN_BEHAVIORAL of FA_22 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_23 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_23;

architecture SYN_BEHAVIORAL of FA_23 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_24 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_24;

architecture SYN_BEHAVIORAL of FA_24 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U2 : INV_X1 port map( A => n10, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n10);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_25 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_25;

architecture SYN_BEHAVIORAL of FA_25 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U2 : INV_X1 port map( A => n13, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n13);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_26 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_26;

architecture SYN_BEHAVIORAL of FA_26 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_27 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_27;

architecture SYN_BEHAVIORAL of FA_27 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_28 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_28;

architecture SYN_BEHAVIORAL of FA_28 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U2 : INV_X1 port map( A => n10, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n10);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U5 : CLKBUF_X1 port map( A => n9, Z => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_29 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_29;

architecture SYN_BEHAVIORAL of FA_29 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U2 : INV_X1 port map( A => n9, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n8, B2 => Ci, ZN => n9);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_30 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_30;

architecture SYN_BEHAVIORAL of FA_30 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_31 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_31;

architecture SYN_BEHAVIORAL of FA_31 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_32 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_32;

architecture SYN_BEHAVIORAL of FA_32 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8, n9, n10 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U2 : INV_X1 port map( A => n9, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n8, B2 => Ci, ZN => n9);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n8);
   U5 : CLKBUF_X1 port map( A => n8, Z => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_33 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_33;

architecture SYN_BEHAVIORAL of FA_33 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U2 : INV_X1 port map( A => n9, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n8, B2 => Ci, ZN => n9);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_34 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_34;

architecture SYN_BEHAVIORAL of FA_34 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_35 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_35;

architecture SYN_BEHAVIORAL of FA_35 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_36 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_36;

architecture SYN_BEHAVIORAL of FA_36 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U2 : INV_X1 port map( A => n10, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n10);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U5 : CLKBUF_X1 port map( A => n9, Z => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_37 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_37;

architecture SYN_BEHAVIORAL of FA_37 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U2 : INV_X1 port map( A => n9, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n8, B2 => Ci, ZN => n9);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_38 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_38;

architecture SYN_BEHAVIORAL of FA_38 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_39 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_39;

architecture SYN_BEHAVIORAL of FA_39 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_40 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_40;

architecture SYN_BEHAVIORAL of FA_40 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8, n9, n10 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n10, Z => S);
   U2 : INV_X1 port map( A => n9, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n8, B2 => Ci, ZN => n9);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n8);
   U5 : CLKBUF_X1 port map( A => n8, Z => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_41 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_41;

architecture SYN_BEHAVIORAL of FA_41 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U2 : INV_X1 port map( A => n9, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n8, B2 => Ci, ZN => n9);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_42 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_42;

architecture SYN_BEHAVIORAL of FA_42 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_43 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_43;

architecture SYN_BEHAVIORAL of FA_43 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7, n8, n9, n10 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n9);
   U5 : NAND2_X1 port map( A1 => n7, A2 => Ci, ZN => n10);
   U6 : AND2_X1 port map( A1 => n9, A2 => n10, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_44 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_44;

architecture SYN_BEHAVIORAL of FA_44 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => n8, B => Ci, Z => S);
   U2 : INV_X1 port map( A => n9, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n8, B2 => Ci, ZN => n9);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_45 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_45;

architecture SYN_BEHAVIORAL of FA_45 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U2 : INV_X1 port map( A => n9, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n8, B2 => Ci, ZN => n9);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_46 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_46;

architecture SYN_BEHAVIORAL of FA_46 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_47 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_47;

architecture SYN_BEHAVIORAL of FA_47 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_48 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_48;

architecture SYN_BEHAVIORAL of FA_48 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_49 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_49;

architecture SYN_BEHAVIORAL of FA_49 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U2 : INV_X1 port map( A => n9, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n8, B2 => Ci, ZN => n9);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_50 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_50;

architecture SYN_BEHAVIORAL of FA_50 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_51 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_51;

architecture SYN_BEHAVIORAL of FA_51 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_52 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_52;

architecture SYN_BEHAVIORAL of FA_52 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U2 : INV_X1 port map( A => n9, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n8, B2 => Ci, ZN => n9);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_53 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_53;

architecture SYN_BEHAVIORAL of FA_53 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U2 : INV_X1 port map( A => n9, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n8, B2 => Ci, ZN => n9);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_54 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_54;

architecture SYN_BEHAVIORAL of FA_54 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_55 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_55;

architecture SYN_BEHAVIORAL of FA_55 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_56 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_56;

architecture SYN_BEHAVIORAL of FA_56 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U2 : INV_X1 port map( A => n9, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n8, B2 => Ci, ZN => n9);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_57 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_57;

architecture SYN_BEHAVIORAL of FA_57 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8, n9 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U2 : INV_X1 port map( A => n9, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n8, B2 => Ci, ZN => n9);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_58 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_58;

architecture SYN_BEHAVIORAL of FA_58 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n10, n11, n12 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => n10, B => n8, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n8);
   U2 : NAND2_X1 port map( A1 => n11, A2 => n12, ZN => Co);
   U3 : CLKBUF_X1 port map( A => Ci, Z => n10);
   U5 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n11);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => n8, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_59 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_59;

architecture SYN_BEHAVIORAL of FA_59 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_60 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_60;

architecture SYN_BEHAVIORAL of FA_60 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n12, n13 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => n12, B => Ci, Z => S);
   U2 : INV_X1 port map( A => n13, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n12, B2 => Ci, ZN => n13);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_61 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_61;

architecture SYN_BEHAVIORAL of FA_61 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U2 : INV_X1 port map( A => n10, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n10);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_62 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_62;

architecture SYN_BEHAVIORAL of FA_62 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_63 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_63;

architecture SYN_BEHAVIORAL of FA_63 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7, n8, n9 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => n9, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U5 : CLKBUF_X1 port map( A => Ci, Z => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_0 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_0;

architecture SYN_BEHAVIORAL of FA_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n10, n12, n13, n14, n15 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => n10, B => Ci, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);
   U2 : OAI22_X1 port map( A1 => n12, A2 => n13, B1 => n14, B2 => n15, ZN => Co
                           );
   U3 : INV_X1 port map( A => B, ZN => n12);
   U5 : INV_X1 port map( A => A, ZN => n13);
   U6 : INV_X1 port map( A => n10, ZN => n14);
   U7 : INV_X1 port map( A => Ci, ZN => n15);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_N4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end RCA_N4_1;

architecture SYN_STRUCTURAL of RCA_N4_1 is

   component FA_1
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_3
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_4
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port, net4521 : std_logic;

begin
   
   FAI_1 : FA_4 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_3 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_2 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_1 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net4521);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_N4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end RCA_N4_2;

architecture SYN_STRUCTURAL of RCA_N4_2 is

   component FA_5
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_6
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_7
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_8
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port, net4521 : std_logic;

begin
   
   FAI_1 : FA_8 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_7 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_6 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_5 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net4521);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_N4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end RCA_N4_3;

architecture SYN_STRUCTURAL of RCA_N4_3 is

   component FA_9
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_10
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_11
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_12
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port, net4521 : std_logic;

begin
   
   FAI_1 : FA_12 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_11 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_10 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_9 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net4521);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_N4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end RCA_N4_4;

architecture SYN_STRUCTURAL of RCA_N4_4 is

   component FA_13
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_14
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_15
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_16
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port, net4521 : std_logic;

begin
   
   FAI_1 : FA_16 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_15 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_14 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_13 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net4521);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_N4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end RCA_N4_5;

architecture SYN_STRUCTURAL of RCA_N4_5 is

   component FA_17
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_18
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_19
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_20
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port, net4521 : std_logic;

begin
   
   FAI_1 : FA_20 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_19 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_18 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_17 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net4521);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_N4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end RCA_N4_6;

architecture SYN_STRUCTURAL of RCA_N4_6 is

   component FA_21
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_22
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_23
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_24
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port, net4521 : std_logic;

begin
   
   FAI_1 : FA_24 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_23 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_22 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_21 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net4521);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_N4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end RCA_N4_7;

architecture SYN_STRUCTURAL of RCA_N4_7 is

   component FA_25
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_26
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_27
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_28
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port, net4521 : std_logic;

begin
   
   FAI_1 : FA_28 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_27 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_26 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_25 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net4521);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_N4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end RCA_N4_8;

architecture SYN_STRUCTURAL of RCA_N4_8 is

   component FA_29
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_30
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_31
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_32
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port, net4521 : std_logic;

begin
   
   FAI_1 : FA_32 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_31 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_30 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_29 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net4521);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_N4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end RCA_N4_9;

architecture SYN_STRUCTURAL of RCA_N4_9 is

   component FA_33
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_34
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_35
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_36
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port, net4521 : std_logic;

begin
   
   FAI_1 : FA_36 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_35 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_34 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_33 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net4521);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_N4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end RCA_N4_10;

architecture SYN_STRUCTURAL of RCA_N4_10 is

   component FA_37
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_38
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_39
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_40
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port, net4521 : std_logic;

begin
   
   FAI_1 : FA_40 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_39 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_38 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_37 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net4521);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_N4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end RCA_N4_11;

architecture SYN_STRUCTURAL of RCA_N4_11 is

   component FA_41
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_42
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_43
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_44
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port, net4521 : std_logic;

begin
   
   FAI_1 : FA_44 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_43 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_42 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_41 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net4521);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_N4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end RCA_N4_12;

architecture SYN_STRUCTURAL of RCA_N4_12 is

   component FA_45
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_46
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_47
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_48
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port, net4521 : std_logic;

begin
   
   FAI_1 : FA_48 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_47 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_46 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_45 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net4521);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_N4_13 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end RCA_N4_13;

architecture SYN_STRUCTURAL of RCA_N4_13 is

   component FA_49
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_50
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_51
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_52
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port, net4521 : std_logic;

begin
   
   FAI_1 : FA_52 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_51 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_50 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_49 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net4521);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_N4_14 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end RCA_N4_14;

architecture SYN_STRUCTURAL of RCA_N4_14 is

   component FA_53
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_54
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_55
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_56
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port, net4521 : std_logic;

begin
   
   FAI_1 : FA_56 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_55 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_54 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_53 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net4521);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_N4_15 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end RCA_N4_15;

architecture SYN_STRUCTURAL of RCA_N4_15 is

   component FA_57
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_58
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_59
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_60
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port, net4521 : std_logic;

begin
   
   FAI_1 : FA_60 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_59 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_58 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_57 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net4521);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_N4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end RCA_N4_0;

architecture SYN_STRUCTURAL of RCA_N4_0 is

   component FA_61
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_62
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_63
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_0
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port, net4521 : std_logic;

begin
   
   FAI_1 : FA_0 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_63 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_62 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_61 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net4521);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity CSB_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_1;

architecture SYN_structural of CSB_1 is

   component MUX2_X2
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component RCA_N4_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_2
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA_0 : RCA_N4_2 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => sum0_3_port, 
                           S(2) => sum0_2_port, S(1) => sum0_1_port, S(0) => 
                           sum0_0_port);
   RCA_1 : RCA_N4_1 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => sum1_3_port, 
                           S(2) => sum1_2_port, S(1) => sum1_1_port, S(0) => 
                           sum1_0_port);
   U3 : MUX2_X2 port map( A => sum0_3_port, B => sum1_3_port, S => Ci, Z => 
                           S(3));
   U4 : MUX2_X1 port map( A => sum0_2_port, B => sum1_2_port, S => Ci, Z => 
                           S(2));
   U5 : MUX2_X2 port map( A => sum0_0_port, B => sum1_0_port, S => Ci, Z => 
                           S(0));
   U6 : MUX2_X2 port map( A => sum0_1_port, B => sum1_1_port, S => Ci, Z => 
                           S(1));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity CSB_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_2;

architecture SYN_structural of CSB_2 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component RCA_N4_3
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   U4 : MUX2_X1 port map( A => sum0_2_port, B => sum1_2_port, S => Ci, Z => 
                           S(2));
   U5 : MUX2_X1 port map( A => sum0_1_port, B => sum1_1_port, S => Ci, Z => 
                           S(1));
   RCA_0 : RCA_N4_4 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => sum0_3_port, 
                           S(2) => sum0_2_port, S(1) => sum0_1_port, S(0) => 
                           sum0_0_port);
   RCA_1 : RCA_N4_3 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => sum1_3_port, 
                           S(2) => sum1_2_port, S(1) => sum1_1_port, S(0) => 
                           sum1_0_port);
   U3 : MUX2_X1 port map( A => sum0_0_port, B => sum1_0_port, S => Ci, Z => 
                           S(0));
   U6 : MUX2_X1 port map( A => sum0_3_port, B => sum1_3_port, S => Ci, Z => 
                           S(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity CSB_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_3;

architecture SYN_structural of CSB_3 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component RCA_N4_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_6
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   U3 : MUX2_X1 port map( A => sum0_3_port, B => sum1_3_port, S => Ci, Z => 
                           S(3));
   U4 : MUX2_X1 port map( A => sum0_2_port, B => sum1_2_port, S => Ci, Z => 
                           S(2));
   RCA_0 : RCA_N4_6 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => sum0_3_port, 
                           S(2) => sum0_2_port, S(1) => sum0_1_port, S(0) => 
                           sum0_0_port);
   RCA_1 : RCA_N4_5 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => sum1_3_port, 
                           S(2) => sum1_2_port, S(1) => sum1_1_port, S(0) => 
                           sum1_0_port);
   U5 : MUX2_X1 port map( A => sum0_0_port, B => sum1_0_port, S => Ci, Z => 
                           S(0));
   U6 : MUX2_X1 port map( A => sum0_1_port, B => sum1_1_port, S => Ci, Z => 
                           S(1));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity CSB_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_4;

architecture SYN_structural of CSB_4 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component RCA_N4_7
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_8
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA_0 : RCA_N4_8 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => sum0_3_port, 
                           S(2) => sum0_2_port, S(1) => sum0_1_port, S(0) => 
                           sum0_0_port);
   RCA_1 : RCA_N4_7 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => sum1_3_port, 
                           S(2) => sum1_2_port, S(1) => sum1_1_port, S(0) => 
                           sum1_0_port);
   U5 : MUX2_X1 port map( A => sum0_1_port, B => sum1_1_port, S => Ci, Z => 
                           S(1));
   U4 : MUX2_X1 port map( A => sum0_2_port, B => sum1_2_port, S => Ci, Z => 
                           S(2));
   U3 : MUX2_X1 port map( A => sum0_3_port, B => sum1_3_port, S => Ci, Z => 
                           S(3));
   U6 : MUX2_X1 port map( A => sum0_0_port, B => sum1_0_port, S => Ci, Z => 
                           S(0));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity CSB_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_5;

architecture SYN_structural of CSB_5 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component RCA_N4_9
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_10
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   U3 : MUX2_X1 port map( A => sum0_3_port, B => sum1_3_port, S => Ci, Z => 
                           S(3));
   U4 : MUX2_X1 port map( A => sum0_2_port, B => sum1_2_port, S => Ci, Z => 
                           S(2));
   U5 : MUX2_X1 port map( A => sum0_1_port, B => sum1_1_port, S => Ci, Z => 
                           S(1));
   RCA_0 : RCA_N4_10 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port);
   RCA_1 : RCA_N4_9 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => sum1_3_port, 
                           S(2) => sum1_2_port, S(1) => sum1_1_port, S(0) => 
                           sum1_0_port);
   U6 : MUX2_X1 port map( A => sum0_0_port, B => sum1_0_port, S => Ci, Z => 
                           S(0));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity CSB_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_6;

architecture SYN_structural of CSB_6 is

   component RCA_N4_11
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_12
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   U3 : MUX2_X1 port map( A => sum0_3_port, B => sum1_3_port, S => Ci, Z => 
                           S(3));
   U4 : MUX2_X1 port map( A => sum0_2_port, B => sum1_2_port, S => Ci, Z => 
                           S(2));
   U5 : MUX2_X1 port map( A => sum0_1_port, B => sum1_1_port, S => Ci, Z => 
                           S(1));
   U6 : MUX2_X1 port map( A => sum0_0_port, B => sum1_0_port, S => Ci, Z => 
                           S(0));
   RCA_0 : RCA_N4_12 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port);
   RCA_1 : RCA_N4_11 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity CSB_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_7;

architecture SYN_structural of CSB_7 is

   component MUX2_X2
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component RCA_N4_13
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_14
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   U4 : MUX2_X1 port map( A => sum0_2_port, B => sum1_2_port, S => Ci, Z => 
                           S(2));
   U5 : MUX2_X1 port map( A => sum0_1_port, B => sum1_1_port, S => Ci, Z => 
                           S(1));
   U6 : MUX2_X1 port map( A => sum0_0_port, B => sum1_0_port, S => Ci, Z => 
                           S(0));
   RCA_0 : RCA_N4_14 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port);
   RCA_1 : RCA_N4_13 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port);
   U3 : MUX2_X2 port map( A => sum0_3_port, B => sum1_3_port, S => Ci, Z => 
                           S(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity CSB_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_0;

architecture SYN_structural of CSB_0 is

   component MUX2_X2
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component RCA_N4_15
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   U4 : MUX2_X1 port map( A => sum0_2_port, B => sum1_2_port, S => Ci, Z => 
                           S(2));
   U5 : MUX2_X1 port map( A => sum0_1_port, B => sum1_1_port, S => Ci, Z => 
                           S(1));
   U6 : MUX2_X1 port map( A => sum0_0_port, B => sum1_0_port, S => Ci, Z => 
                           S(0));
   RCA_0 : RCA_N4_0 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => sum0_3_port, 
                           S(2) => sum0_2_port, S(1) => sum0_1_port, S(0) => 
                           sum0_0_port);
   RCA_1 : RCA_N4_15 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port);
   U3 : MUX2_X2 port map( A => sum0_3_port, B => sum1_3_port, S => Ci, Z => 
                           S(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_1 is

   port( pi, gi, gj : in std_logic;  gout : out std_logic);

end G_1;

architecture SYN_behav of G_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U1 : OAI21_X2 port map( B1 => n5, B2 => n6, A => n7, ZN => gout);
   U2 : INV_X1 port map( A => gj, ZN => n5);
   U3 : INV_X1 port map( A => pi, ZN => n6);
   U4 : INV_X1 port map( A => gi, ZN => n7);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_2 is

   port( pi, gi, gj : in std_logic;  gout : out std_logic);

end G_2;

architecture SYN_behav of G_2 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gj, B2 => pi, A => gi, ZN => n4);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_3 is

   port( pi, gi, gj : in std_logic;  gout : out std_logic);

end G_3;

architecture SYN_behav of G_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n6, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gj, B2 => pi, A => gi, ZN => n6);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_4 is

   port( pi, gi, gj : in std_logic;  gout : out std_logic);

end G_4;

architecture SYN_behav of G_4 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => gout);
   U2 : AOI21_X1 port map( B1 => pi, B2 => gj, A => gi, ZN => n4);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_1 is

   port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);

end PG_1;

architecture SYN_behav of PG_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => pj, A2 => pi, ZN => pout);
   U2 : INV_X1 port map( A => n4, ZN => gout);
   U3 : AOI21_X1 port map( B1 => gj, B2 => pi, A => gi, ZN => n4);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_2 is

   port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);

end PG_2;

architecture SYN_behav of PG_2 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => pj, A2 => pi, ZN => pout);
   U2 : INV_X1 port map( A => n4, ZN => gout);
   U3 : AOI21_X1 port map( B1 => gj, B2 => pi, A => gi, ZN => n4);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_5 is

   port( pi, gi, gj : in std_logic;  gout : out std_logic);

end G_5;

architecture SYN_behav of G_5 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => gout);
   U2 : AOI21_X1 port map( B1 => pi, B2 => gj, A => gi, ZN => n4);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_6 is

   port( pi, gi, gj : in std_logic;  gout : out std_logic);

end G_6;

architecture SYN_behav of G_6 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n6, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gj, B2 => pi, A => gi, ZN => n6);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_3 is

   port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);

end PG_3;

architecture SYN_behav of PG_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => pj, A2 => pi, ZN => pout);
   U2 : INV_X1 port map( A => n4, ZN => gout);
   U3 : AOI21_X1 port map( B1 => gj, B2 => pi, A => gi, ZN => n4);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_4 is

   port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);

end PG_4;

architecture SYN_behav of PG_4 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => pj, A2 => pi, ZN => pout);
   U2 : INV_X1 port map( A => n7, ZN => gout);
   U3 : AOI21_X1 port map( B1 => gj, B2 => pi, A => gi, ZN => n7);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_5 is

   port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);

end PG_5;

architecture SYN_behav of PG_5 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => pj, A2 => pi, ZN => pout);
   U2 : INV_X1 port map( A => n6, ZN => gout);
   U3 : AOI21_X1 port map( B1 => gj, B2 => pi, A => gi, ZN => n6);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_7 is

   port( pi, gi, gj : in std_logic;  gout : out std_logic);

end G_7;

architecture SYN_behav of G_7 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gj, B2 => pi, A => gi, ZN => n4);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_6 is

   port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);

end PG_6;

architecture SYN_behav of PG_6 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => pj, A2 => pi, ZN => pout);
   U2 : INV_X1 port map( A => n4, ZN => gout);
   U3 : AOI21_X1 port map( B1 => gj, B2 => pi, A => gi, ZN => n4);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_7 is

   port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);

end PG_7;

architecture SYN_behav of PG_7 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => pj, A2 => pi, ZN => pout);
   U2 : INV_X1 port map( A => n4, ZN => gout);
   U3 : AOI21_X1 port map( B1 => gj, B2 => pi, A => gi, ZN => n4);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_8 is

   port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);

end PG_8;

architecture SYN_behav of PG_8 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => pj, A2 => pi, ZN => pout);
   U2 : INV_X1 port map( A => n4, ZN => gout);
   U3 : AOI21_X1 port map( B1 => gj, B2 => pi, A => gi, ZN => n4);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_9 is

   port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);

end PG_9;

architecture SYN_behav of PG_9 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => pj, A2 => pi, ZN => pout);
   U2 : INV_X1 port map( A => n4, ZN => gout);
   U3 : AOI21_X1 port map( B1 => gj, B2 => pi, A => gi, ZN => n4);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_10 is

   port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);

end PG_10;

architecture SYN_behav of PG_10 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => pj, A2 => pi, ZN => pout);
   U2 : INV_X1 port map( A => n4, ZN => gout);
   U3 : AOI21_X1 port map( B1 => gj, B2 => pi, A => gi, ZN => n4);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_11 is

   port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);

end PG_11;

architecture SYN_behav of PG_11 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => pj, A2 => pi, ZN => pout);
   U2 : INV_X1 port map( A => n4, ZN => gout);
   U3 : AOI21_X1 port map( B1 => gj, B2 => pi, A => gi, ZN => n4);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_12 is

   port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);

end PG_12;

architecture SYN_behav of PG_12 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => pj, A2 => pi, ZN => pout);
   U2 : INV_X1 port map( A => n4, ZN => gout);
   U3 : AOI21_X1 port map( B1 => gj, B2 => pi, A => gi, ZN => n4);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_8 is

   port( pi, gi, gj : in std_logic;  gout : out std_logic);

end G_8;

architecture SYN_behav of G_8 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gj, B2 => pi, A => gi, ZN => n4);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_13 is

   port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);

end PG_13;

architecture SYN_behav of PG_13 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => pj, A2 => pi, ZN => pout);
   U2 : INV_X1 port map( A => n4, ZN => gout);
   U3 : AOI21_X1 port map( B1 => gj, B2 => pi, A => gi, ZN => n4);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_14 is

   port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);

end PG_14;

architecture SYN_behav of PG_14 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => pj, A2 => pi, ZN => pout);
   U2 : INV_X1 port map( A => n4, ZN => gout);
   U3 : AOI21_X1 port map( B1 => gj, B2 => pi, A => gi, ZN => n4);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_15 is

   port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);

end PG_15;

architecture SYN_behav of PG_15 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => pj, A2 => pi, ZN => pout);
   U2 : INV_X1 port map( A => n4, ZN => gout);
   U3 : AOI21_X1 port map( B1 => gj, B2 => pi, A => gi, ZN => n4);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_16 is

   port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);

end PG_16;

architecture SYN_behav of PG_16 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => pj, A2 => pi, ZN => pout);
   U2 : INV_X1 port map( A => n4, ZN => gout);
   U3 : AOI21_X1 port map( B1 => gj, B2 => pi, A => gi, ZN => n4);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_17 is

   port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);

end PG_17;

architecture SYN_behav of PG_17 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => pi, A2 => pj, ZN => pout);
   U2 : INV_X1 port map( A => n4, ZN => gout);
   U3 : AOI21_X1 port map( B1 => pi, B2 => gj, A => gi, ZN => n4);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_18 is

   port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);

end PG_18;

architecture SYN_behav of PG_18 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => pj, A2 => pi, ZN => pout);
   U2 : INV_X1 port map( A => n4, ZN => gout);
   U3 : AOI21_X1 port map( B1 => gj, B2 => pi, A => gi, ZN => n4);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_19 is

   port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);

end PG_19;

architecture SYN_behav of PG_19 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => pj, A2 => pi, ZN => pout);
   U2 : INV_X1 port map( A => n4, ZN => gout);
   U3 : AOI21_X1 port map( B1 => pi, B2 => gj, A => gi, ZN => n4);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_20 is

   port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);

end PG_20;

architecture SYN_behav of PG_20 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => pj, A2 => pi, ZN => pout);
   U2 : INV_X1 port map( A => n4, ZN => gout);
   U3 : AOI21_X1 port map( B1 => gj, B2 => pi, A => gi, ZN => n4);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_21 is

   port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);

end PG_21;

architecture SYN_behav of PG_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7, n8 : std_logic;

begin
   
   U1 : OAI21_X1 port map( B1 => n6, B2 => n7, A => n8, ZN => gout);
   U2 : INV_X1 port map( A => pi, ZN => n6);
   U3 : INV_X1 port map( A => gj, ZN => n7);
   U4 : INV_X1 port map( A => gi, ZN => n8);
   U5 : AND2_X1 port map( A1 => pi, A2 => pj, ZN => pout);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_22 is

   port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);

end PG_22;

architecture SYN_behav of PG_22 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => pi, A2 => pj, ZN => pout);
   U2 : INV_X1 port map( A => n5, ZN => gout);
   U3 : AOI21_X1 port map( B1 => pi, B2 => gj, A => gi, ZN => n5);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_23 is

   port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);

end PG_23;

architecture SYN_behav of PG_23 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => pi, A2 => pj, ZN => pout);
   U2 : INV_X1 port map( A => n5, ZN => gout);
   U3 : AOI21_X1 port map( B1 => pi, B2 => gj, A => gi, ZN => n5);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_24 is

   port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);

end PG_24;

architecture SYN_behav of PG_24 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => pj, A2 => pi, ZN => pout);
   U2 : INV_X1 port map( A => n5, ZN => gout);
   U3 : AOI21_X1 port map( B1 => gj, B2 => pi, A => gi, ZN => n5);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_25 is

   port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);

end PG_25;

architecture SYN_behav of PG_25 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => pi, A2 => pj, ZN => pout);
   U2 : INV_X1 port map( A => n7, ZN => gout);
   U3 : AOI21_X1 port map( B1 => pi, B2 => gj, A => gi, ZN => n7);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_26 is

   port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);

end PG_26;

architecture SYN_behav of PG_26 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => pi, A2 => pj, ZN => pout);
   U2 : INV_X1 port map( A => n7, ZN => gout);
   U3 : AOI21_X1 port map( B1 => gj, B2 => pi, A => gi, ZN => n7);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_0 is

   port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);

end PG_0;

architecture SYN_behav of PG_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => pi, A2 => pj, ZN => pout);
   U2 : INV_X1 port map( A => n7, ZN => gout);
   U3 : AOI21_X1 port map( B1 => pi, B2 => gj, A => gi, ZN => n7);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_0 is

   port( pi, gi, gj : in std_logic;  gout : out std_logic);

end G_0;

architecture SYN_behav of G_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => gout);
   U2 : AOI21_X1 port map( B1 => gj, B2 => pi, A => gi, ZN => n4);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity prop_gen_1 is

   port( a, b : in std_logic;  prop, gen : out std_logic);

end prop_gen_1;

architecture SYN_behav of prop_gen_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => prop);
   U2 : AND2_X1 port map( A1 => b, A2 => a, ZN => gen);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity prop_gen_2 is

   port( a, b : in std_logic;  prop, gen : out std_logic);

end prop_gen_2;

architecture SYN_behav of prop_gen_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => prop);
   U2 : AND2_X1 port map( A1 => b, A2 => a, ZN => gen);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity prop_gen_3 is

   port( a, b : in std_logic;  prop, gen : out std_logic);

end prop_gen_3;

architecture SYN_behav of prop_gen_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => prop);
   U2 : AND2_X1 port map( A1 => b, A2 => a, ZN => gen);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity prop_gen_4 is

   port( a, b : in std_logic;  prop, gen : out std_logic);

end prop_gen_4;

architecture SYN_behav of prop_gen_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => prop);
   U2 : AND2_X1 port map( A1 => b, A2 => a, ZN => gen);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity prop_gen_5 is

   port( a, b : in std_logic;  prop, gen : out std_logic);

end prop_gen_5;

architecture SYN_behav of prop_gen_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => prop);
   U2 : AND2_X1 port map( A1 => b, A2 => a, ZN => gen);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity prop_gen_6 is

   port( a, b : in std_logic;  prop, gen : out std_logic);

end prop_gen_6;

architecture SYN_behav of prop_gen_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => prop);
   U2 : AND2_X1 port map( A1 => b, A2 => a, ZN => gen);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity prop_gen_7 is

   port( a, b : in std_logic;  prop, gen : out std_logic);

end prop_gen_7;

architecture SYN_behav of prop_gen_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => prop);
   U2 : AND2_X1 port map( A1 => b, A2 => a, ZN => gen);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity prop_gen_8 is

   port( a, b : in std_logic;  prop, gen : out std_logic);

end prop_gen_8;

architecture SYN_behav of prop_gen_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => prop);
   U2 : AND2_X1 port map( A1 => b, A2 => a, ZN => gen);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity prop_gen_9 is

   port( a, b : in std_logic;  prop, gen : out std_logic);

end prop_gen_9;

architecture SYN_behav of prop_gen_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => a, B => b, Z => prop);
   U2 : AND2_X1 port map( A1 => b, A2 => a, ZN => gen);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity prop_gen_10 is

   port( a, b : in std_logic;  prop, gen : out std_logic);

end prop_gen_10;

architecture SYN_behav of prop_gen_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => prop);
   U2 : AND2_X1 port map( A1 => b, A2 => a, ZN => gen);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity prop_gen_11 is

   port( a, b : in std_logic;  prop, gen : out std_logic);

end prop_gen_11;

architecture SYN_behav of prop_gen_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => prop);
   U2 : AND2_X1 port map( A1 => b, A2 => a, ZN => gen);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity prop_gen_12 is

   port( a, b : in std_logic;  prop, gen : out std_logic);

end prop_gen_12;

architecture SYN_behav of prop_gen_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => prop);
   U2 : AND2_X1 port map( A1 => b, A2 => a, ZN => gen);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity prop_gen_13 is

   port( a, b : in std_logic;  prop, gen : out std_logic);

end prop_gen_13;

architecture SYN_behav of prop_gen_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => prop);
   U2 : AND2_X1 port map( A1 => b, A2 => a, ZN => gen);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity prop_gen_14 is

   port( a, b : in std_logic;  prop, gen : out std_logic);

end prop_gen_14;

architecture SYN_behav of prop_gen_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => prop);
   U2 : AND2_X1 port map( A1 => b, A2 => a, ZN => gen);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity prop_gen_15 is

   port( a, b : in std_logic;  prop, gen : out std_logic);

end prop_gen_15;

architecture SYN_behav of prop_gen_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => prop);
   U2 : AND2_X1 port map( A1 => b, A2 => a, ZN => gen);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity prop_gen_16 is

   port( a, b : in std_logic;  prop, gen : out std_logic);

end prop_gen_16;

architecture SYN_behav of prop_gen_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => prop);
   U2 : AND2_X1 port map( A1 => b, A2 => a, ZN => gen);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity prop_gen_17 is

   port( a, b : in std_logic;  prop, gen : out std_logic);

end prop_gen_17;

architecture SYN_behav of prop_gen_17 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U2 : AND2_X1 port map( A1 => a, A2 => b, ZN => gen);
   U1 : XOR2_X1 port map( A => a, B => b, Z => prop);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity prop_gen_18 is

   port( a, b : in std_logic;  prop, gen : out std_logic);

end prop_gen_18;

architecture SYN_behav of prop_gen_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => prop);
   U2 : AND2_X1 port map( A1 => b, A2 => a, ZN => gen);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity prop_gen_19 is

   port( a, b : in std_logic;  prop, gen : out std_logic);

end prop_gen_19;

architecture SYN_behav of prop_gen_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => prop);
   U2 : AND2_X1 port map( A1 => b, A2 => a, ZN => gen);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity prop_gen_20 is

   port( a, b : in std_logic;  prop, gen : out std_logic);

end prop_gen_20;

architecture SYN_behav of prop_gen_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => prop);
   U2 : AND2_X1 port map( A1 => b, A2 => a, ZN => gen);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity prop_gen_21 is

   port( a, b : in std_logic;  prop, gen : out std_logic);

end prop_gen_21;

architecture SYN_behav of prop_gen_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => a, B => b, Z => prop);
   U2 : AND2_X1 port map( A1 => b, A2 => a, ZN => gen);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity prop_gen_22 is

   port( a, b : in std_logic;  prop, gen : out std_logic);

end prop_gen_22;

architecture SYN_behav of prop_gen_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => prop);
   U2 : AND2_X1 port map( A1 => b, A2 => a, ZN => gen);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity prop_gen_23 is

   port( a, b : in std_logic;  prop, gen : out std_logic);

end prop_gen_23;

architecture SYN_behav of prop_gen_23 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => prop);
   U2 : AND2_X1 port map( A1 => b, A2 => n1, ZN => gen);
   U3 : CLKBUF_X1 port map( A => a, Z => n1);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity prop_gen_24 is

   port( a, b : in std_logic;  prop, gen : out std_logic);

end prop_gen_24;

architecture SYN_behav of prop_gen_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => prop);
   U2 : AND2_X1 port map( A1 => b, A2 => a, ZN => gen);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity prop_gen_25 is

   port( a, b : in std_logic;  prop, gen : out std_logic);

end prop_gen_25;

architecture SYN_behav of prop_gen_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => a, B => b, Z => prop);
   U2 : AND2_X1 port map( A1 => b, A2 => a, ZN => gen);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity prop_gen_26 is

   port( a, b : in std_logic;  prop, gen : out std_logic);

end prop_gen_26;

architecture SYN_behav of prop_gen_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => prop);
   U2 : AND2_X1 port map( A1 => b, A2 => a, ZN => gen);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity prop_gen_27 is

   port( a, b : in std_logic;  prop, gen : out std_logic);

end prop_gen_27;

architecture SYN_behav of prop_gen_27 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => prop);
   U2 : AND2_X1 port map( A1 => b, A2 => a, ZN => gen);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity prop_gen_28 is

   port( a, b : in std_logic;  prop, gen : out std_logic);

end prop_gen_28;

architecture SYN_behav of prop_gen_28 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => prop);
   U2 : AND2_X1 port map( A1 => b, A2 => a, ZN => gen);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity prop_gen_29 is

   port( a, b : in std_logic;  prop, gen : out std_logic);

end prop_gen_29;

architecture SYN_behav of prop_gen_29 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U2 : AND2_X1 port map( A1 => b, A2 => n1, ZN => gen);
   U1 : XOR2_X1 port map( A => b, B => a, Z => prop);
   U3 : CLKBUF_X1 port map( A => a, Z => n1);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity prop_gen_30 is

   port( a, b : in std_logic;  prop, gen : out std_logic);

end prop_gen_30;

architecture SYN_behav of prop_gen_30 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => prop);
   U2 : AND2_X1 port map( A1 => b, A2 => a, ZN => gen);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity prop_gen_0 is

   port( a, b : in std_logic;  prop, gen : out std_logic);

end prop_gen_0;

architecture SYN_behav of prop_gen_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => prop);
   U2 : AND2_X1 port map( A1 => b, A2 => a, ZN => gen);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity prop_gen_Cin is

   port( a, b, cin : in std_logic;  prop, gen : out std_logic);

end prop_gen_Cin;

architecture SYN_Behavioral of prop_gen_Cin is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n20, n21, n22 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n22, Z => prop);
   U5 : OAI21_X1 port map( B1 => a, B2 => b, A => cin, ZN => n20);
   U2 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => gen);
   U3 : NAND2_X1 port map( A1 => a, A2 => b, ZN => n21);
   U4 : CLKBUF_X1 port map( A => a, Z => n22);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity shifter is

   port( R : in std_logic_vector (31 downto 0);  Offset : in std_logic_vector 
         (4 downto 0);  Conf : in std_logic_vector (0 to 1);  Shift_OUT : out 
         std_logic_vector (31 downto 0));

end shifter;

architecture SYN_Struct of shifter is

   component AOI221_X4
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, 
      n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, 
      n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, 
      n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, 
      n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, 
      n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, 
      n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, 
      n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, 
      n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, 
      n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, 
      n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, 
      n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, 
      n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, 
      n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, 
      n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, 
      n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, 
      n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, 
      n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n461, n462, 
      n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, 
      n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, 
      n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497 : 
      std_logic;

begin
   
   U2 : AOI221_X1 port map( B1 => n324, B2 => R(21), C1 => n325, C2 => R(5), A 
                           => n479, ZN => n281);
   U3 : AOI221_X1 port map( B1 => n324, B2 => R(25), C1 => n325, C2 => R(9), A 
                           => n326, ZN => n256);
   U4 : AOI222_X1 port map( A1 => n423, A2 => R(31), B1 => R(7), B2 => n298, C1
                           => R(15), C2 => n299, ZN => n430);
   U5 : NOR3_X2 port map( A1 => n470, A2 => Offset(3), A3 => n372, ZN => n324);
   U6 : NOR2_X2 port map( A1 => n486, A2 => n487, ZN => n257);
   U7 : NOR2_X2 port map( A1 => n483, A2 => n486, ZN => n259);
   U8 : NOR3_X2 port map( A1 => Offset(3), A2 => Offset(4), A3 => n470, ZN => 
                           n325);
   U9 : NOR3_X2 port map( A1 => n371, A2 => Offset(3), A3 => n372, ZN => n338);
   U10 : NOR3_X4 port map( A1 => n470, A2 => Offset(4), A3 => n370, ZN => n423)
                           ;
   U11 : NOR2_X2 port map( A1 => n484, A2 => n487, ZN => n270);
   U12 : NOR3_X4 port map( A1 => n371, A2 => Offset(4), A3 => n370, ZN => n298)
                           ;
   U13 : NOR2_X4 port map( A1 => n483, A2 => n484, ZN => n268);
   U14 : NOR3_X4 port map( A1 => Offset(3), A2 => Offset(4), A3 => n371, ZN => 
                           n299);
   U15 : MUX2_X1 port map( A => n247, B => n248, S => Offset(0), Z => 
                           Shift_OUT(9));
   U16 : MUX2_X1 port map( A => n249, B => n247, S => Offset(0), Z => 
                           Shift_OUT(8));
   U17 : INV_X1 port map( A => n250, ZN => n247);
   U18 : OAI221_X1 port map( B1 => n251, B2 => n252, C1 => n253, C2 => n254, A 
                           => n255, ZN => n250);
   U19 : AOI22_X1 port map( A1 => n256, A2 => n257, B1 => n258, B2 => n259, ZN 
                           => n255);
   U20 : MUX2_X1 port map( A => n260, B => n249, S => Offset(0), Z => 
                           Shift_OUT(7));
   U21 : INV_X1 port map( A => n261, ZN => n249);
   U22 : OAI221_X1 port map( B1 => n262, B2 => n263, C1 => n264, C2 => n265, A 
                           => n266, ZN => n261);
   U23 : AOI22_X1 port map( A1 => n267, A2 => n268, B1 => n269, B2 => n270, ZN 
                           => n266);
   U24 : MUX2_X1 port map( A => n271, B => n260, S => Offset(0), Z => 
                           Shift_OUT(6));
   U25 : INV_X1 port map( A => n272, ZN => n260);
   U26 : OAI221_X1 port map( B1 => n251, B2 => n254, C1 => n262, C2 => n273, A 
                           => n274, ZN => n272);
   U27 : AOI22_X1 port map( A1 => n256, A2 => n259, B1 => n258, B2 => n270, ZN 
                           => n274);
   U28 : INV_X1 port map( A => n275, ZN => n273);
   U29 : MUX2_X1 port map( A => n276, B => n271, S => Offset(0), Z => 
                           Shift_OUT(5));
   U30 : INV_X1 port map( A => n277, ZN => n271);
   U31 : OAI221_X1 port map( B1 => n265, B2 => n263, C1 => n264, C2 => n253, A 
                           => n278, ZN => n277);
   U32 : AOI22_X1 port map( A1 => n269, A2 => n268, B1 => n279, B2 => n257, ZN 
                           => n278);
   U33 : MUX2_X1 port map( A => n280, B => n276, S => Offset(0), Z => 
                           Shift_OUT(4));
   U34 : AOI221_X1 port map( B1 => n259, B2 => n275, C1 => n257, C2 => n281, A 
                           => n282, ZN => n276);
   U35 : INV_X1 port map( A => n283, ZN => n282);
   U36 : AOI22_X1 port map( A1 => n256, A2 => n270, B1 => n258, B2 => n268, ZN 
                           => n283);
   U37 : MUX2_X1 port map( A => n284, B => n280, S => Offset(0), Z => 
                           Shift_OUT(3));
   U38 : INV_X1 port map( A => n285, ZN => n280);
   U39 : OAI221_X1 port map( B1 => n253, B2 => n263, C1 => n264, C2 => n251, A 
                           => n286, ZN => n285);
   U40 : AOI22_X1 port map( A1 => n287, A2 => n257, B1 => n279, B2 => n259, ZN 
                           => n286);
   U41 : INV_X1 port map( A => n288, ZN => n279);
   U42 : INV_X1 port map( A => n289, ZN => n263);
   U43 : MUX2_X1 port map( A => n290, B => n291, S => Offset(0), Z => 
                           Shift_OUT(31));
   U44 : OAI221_X1 port map( B1 => n292, B2 => n251, C1 => n293, C2 => n253, A 
                           => n294, ZN => n291);
   U45 : AOI22_X1 port map( A1 => n259, A2 => n295, B1 => n257, B2 => n296, ZN 
                           => n294);
   U46 : INV_X1 port map( A => n297, ZN => n295);
   U47 : AOI221_X1 port map( B1 => R(22), B2 => n298, C1 => R(30), C2 => n299, 
                           A => n300, ZN => n292);
   U48 : OAI221_X1 port map( B1 => n301, B2 => n302, C1 => n303, C2 => n304, A 
                           => n305, ZN => n300);
   U49 : MUX2_X1 port map( A => n306, B => n290, S => Offset(0), Z => 
                           Shift_OUT(30));
   U50 : INV_X1 port map( A => n307, ZN => n290);
   U51 : OAI221_X1 port map( B1 => n308, B2 => n309, C1 => n253, C2 => n310, A 
                           => n311, ZN => n307);
   U52 : AOI22_X1 port map( A1 => n312, A2 => n259, B1 => n313, B2 => n257, ZN 
                           => n311);
   U53 : OAI221_X1 port map( B1 => n314, B2 => n315, C1 => n316, C2 => n317, A 
                           => n268, ZN => n309);
   U54 : OAI221_X1 port map( B1 => n318, B2 => n302, C1 => n319, C2 => n304, A 
                           => n305, ZN => n308);
   U55 : MUX2_X1 port map( A => n320, B => n284, S => Offset(0), Z => 
                           Shift_OUT(2));
   U56 : AOI221_X1 port map( B1 => n257, B2 => n321, C1 => n270, C2 => n275, A 
                           => n322, ZN => n284);
   U57 : INV_X1 port map( A => n323, ZN => n322);
   U58 : AOI22_X1 port map( A1 => n256, A2 => n268, B1 => n281, B2 => n259, ZN 
                           => n323);
   U59 : OAI221_X1 port map( B1 => n327, B2 => n328, C1 => n329, C2 => n316, A 
                           => n330, ZN => n326);
   U60 : MUX2_X1 port map( A => n331, B => n306, S => Offset(0), Z => 
                           Shift_OUT(29));
   U61 : AOI221_X1 port map( B1 => n268, B2 => n293, C1 => n270, C2 => n297, A 
                           => n332, ZN => n306);
   U62 : OAI22_X1 port map( A1 => n296, A2 => n265, B1 => n333, B2 => n262, ZN 
                           => n332);
   U63 : INV_X1 port map( A => n334, ZN => n293);
   U64 : OAI221_X1 port map( B1 => n316, B2 => n335, C1 => n314, C2 => n336, A 
                           => n337, ZN => n334);
   U66 : MUX2_X1 port map( A => n341, B => n331, S => Offset(0), Z => 
                           Shift_OUT(28));
   U67 : INV_X1 port map( A => n342, ZN => n331);
   U68 : OAI221_X1 port map( B1 => n251, B2 => n310, C1 => n253, C2 => n343, A 
                           => n344, ZN => n342);
   U69 : AOI22_X1 port map( A1 => n313, A2 => n259, B1 => n345, B2 => n257, ZN 
                           => n344);
   U70 : OAI221_X1 port map( B1 => n316, B2 => n346, C1 => n314, C2 => n347, A 
                           => n348, ZN => n310);
   U72 : MUX2_X1 port map( A => n349, B => n341, S => Offset(0), Z => 
                           Shift_OUT(27));
   U73 : AOI221_X1 port map( B1 => n268, B2 => n297, C1 => n270, C2 => n350, A 
                           => n351, ZN => n341);
   U74 : OAI22_X1 port map( A1 => n333, A2 => n265, B1 => n352, B2 => n262, ZN 
                           => n351);
   U75 : AOI221_X1 port map( B1 => R(18), B2 => n298, C1 => n299, C2 => R(26), 
                           A => n353, ZN => n297);
   U76 : OAI221_X1 port map( B1 => n304, B2 => n354, C1 => n302, C2 => n355, A 
                           => n305, ZN => n353);
   U77 : INV_X1 port map( A => n339, ZN => n302);
   U78 : INV_X1 port map( A => n338, ZN => n304);
   U79 : MUX2_X1 port map( A => n356, B => n349, S => Offset(0), Z => 
                           Shift_OUT(26));
   U80 : AOI221_X1 port map( B1 => n268, B2 => n312, C1 => n270, C2 => n313, A 
                           => n357, ZN => n349);
   U81 : OAI22_X1 port map( A1 => n358, A2 => n265, B1 => n359, B2 => n262, ZN 
                           => n357);
   U82 : INV_X1 port map( A => n360, ZN => n313);
   U83 : INV_X1 port map( A => n343, ZN => n312);
   U84 : OAI221_X1 port map( B1 => n314, B2 => n327, C1 => n316, C2 => n361, A 
                           => n362, ZN => n343);
   U86 : MUX2_X1 port map( A => n363, B => n356, S => Offset(0), Z => 
                           Shift_OUT(25));
   U87 : AOI221_X1 port map( B1 => n268, B2 => n350, C1 => n270, C2 => n364, A 
                           => n365, ZN => n356);
   U88 : OAI22_X1 port map( A1 => n352, A2 => n265, B1 => n366, B2 => n262, ZN 
                           => n365);
   U89 : INV_X1 port map( A => n296, ZN => n350);
   U90 : OAI221_X1 port map( B1 => n314, B2 => n367, C1 => n316, C2 => n368, A 
                           => n369, ZN => n296);
   U92 : NOR3_X1 port map( A1 => n370, A2 => n371, A3 => n372, ZN => n339);
   U93 : MUX2_X1 port map( A => n373, B => n363, S => Offset(0), Z => 
                           Shift_OUT(24));
   U94 : AOI221_X1 port map( B1 => n259, B2 => n374, C1 => n257, C2 => n375, A 
                           => n376, ZN => n363);
   U95 : OAI22_X1 port map( A1 => n360, A2 => n251, B1 => n358, B2 => n253, ZN 
                           => n376);
   U96 : OAI211_X1 port map( C1 => n377, C2 => n378, A => n379, B => n380, ZN 
                           => n360);
   U97 : AOI222_X1 port map( A1 => R(23), A2 => n299, B1 => n338, B2 => R(7), 
                           C1 => R(15), C2 => n298, ZN => n380);
   U98 : MUX2_X1 port map( A => n381, B => n373, S => Offset(0), Z => 
                           Shift_OUT(23));
   U99 : AOI221_X1 port map( B1 => n268, B2 => n364, C1 => n270, C2 => n382, A 
                           => n383, ZN => n373);
   U100 : OAI22_X1 port map( A1 => n366, A2 => n265, B1 => n384, B2 => n262, ZN
                           => n383);
   U101 : INV_X1 port map( A => n333, ZN => n364);
   U102 : OAI211_X1 port map( C1 => n378, C2 => n385, A => n379, B => n386, ZN 
                           => n333);
   U103 : AOI222_X1 port map( A1 => R(22), A2 => n299, B1 => n338, B2 => R(6), 
                           C1 => R(14), C2 => n298, ZN => n386);
   U104 : MUX2_X1 port map( A => n387, B => n381, S => Offset(0), Z => 
                           Shift_OUT(22));
   U105 : AOI221_X1 port map( B1 => n268, B2 => n345, C1 => n270, C2 => n374, A
                           => n388, ZN => n381);
   U106 : OAI22_X1 port map( A1 => n389, A2 => n265, B1 => n390, B2 => n262, ZN
                           => n388);
   U107 : INV_X1 port map( A => n358, ZN => n345);
   U108 : OAI211_X1 port map( C1 => n378, C2 => n317, A => n379, B => n391, ZN 
                           => n358);
   U109 : AOI222_X1 port map( A1 => R(21), A2 => n299, B1 => n338, B2 => R(5), 
                           C1 => R(13), C2 => n298, ZN => n391);
   U110 : MUX2_X1 port map( A => n392, B => n387, S => Offset(0), Z => 
                           Shift_OUT(21));
   U111 : AOI221_X1 port map( B1 => n268, B2 => n382, C1 => n270, C2 => n393, A
                           => n394, ZN => n387);
   U112 : OAI22_X1 port map( A1 => n384, A2 => n265, B1 => n395, B2 => n262, ZN
                           => n394);
   U113 : INV_X1 port map( A => n352, ZN => n382);
   U114 : OAI211_X1 port map( C1 => n378, C2 => n335, A => n379, B => n396, ZN 
                           => n352);
   U115 : AOI222_X1 port map( A1 => R(20), A2 => n299, B1 => n338, B2 => R(4), 
                           C1 => R(12), C2 => n298, ZN => n396);
   U116 : MUX2_X1 port map( A => n397, B => n392, S => Offset(0), Z => 
                           Shift_OUT(20));
   U117 : AOI221_X1 port map( B1 => n268, B2 => n374, C1 => n270, C2 => n375, A
                           => n398, ZN => n392);
   U118 : OAI22_X1 port map( A1 => n390, A2 => n265, B1 => n399, B2 => n262, ZN
                           => n398);
   U119 : INV_X1 port map( A => n389, ZN => n375);
   U120 : INV_X1 port map( A => n359, ZN => n374);
   U121 : OAI211_X1 port map( C1 => n378, C2 => n346, A => n379, B => n400, ZN 
                           => n359);
   U122 : AOI222_X1 port map( A1 => R(19), A2 => n299, B1 => n338, B2 => R(3), 
                           C1 => R(11), C2 => n298, ZN => n400);
   U123 : MUX2_X1 port map( A => n401, B => n320, S => Offset(0), Z => 
                           Shift_OUT(1));
   U124 : INV_X1 port map( A => n402, ZN => n320);
   U125 : OAI221_X1 port map( B1 => n262, B2 => n403, C1 => n253, C2 => n288, A
                           => n404, ZN => n402);
   U126 : AOI22_X1 port map( A1 => n289, A2 => n268, B1 => n287, B2 => n259, ZN
                           => n404);
   U127 : AOI221_X1 port map( B1 => n324, B2 => R(24), C1 => n325, C2 => R(8), 
                           A => n405, ZN => n289);
   U128 : OAI221_X1 port map( B1 => n367, B2 => n328, C1 => n406, C2 => n316, A
                           => n330, ZN => n405);
   U129 : MUX2_X1 port map( A => n407, B => n397, S => Offset(0), Z => 
                           Shift_OUT(19));
   U130 : AOI221_X1 port map( B1 => n268, B2 => n393, C1 => n270, C2 => n408, A
                           => n409, ZN => n397);
   U131 : OAI22_X1 port map( A1 => n395, A2 => n265, B1 => n410, B2 => n262, ZN
                           => n409);
   U132 : INV_X1 port map( A => n366, ZN => n393);
   U133 : OAI211_X1 port map( C1 => n411, C2 => n378, A => n379, B => n412, ZN 
                           => n366);
   U134 : AOI222_X1 port map( A1 => R(18), A2 => n299, B1 => n338, B2 => R(2), 
                           C1 => n298, C2 => R(10), ZN => n412);
   U135 : MUX2_X1 port map( A => n413, B => n407, S => Offset(0), Z => 
                           Shift_OUT(18));
   U136 : AOI221_X1 port map( B1 => n259, B2 => n414, C1 => n257, C2 => n415, A
                           => n416, ZN => n407);
   U137 : OAI22_X1 port map( A1 => n389, A2 => n251, B1 => n390, B2 => n253, ZN
                           => n416);
   U138 : OAI211_X1 port map( C1 => n378, C2 => n361, A => n379, B => n417, ZN 
                           => n389);
   U139 : AOI222_X1 port map( A1 => R(17), A2 => n299, B1 => n338, B2 => R(1), 
                           C1 => R(9), C2 => n298, ZN => n417);
   U140 : MUX2_X1 port map( A => n418, B => n413, S => Offset(0), Z => 
                           Shift_OUT(17));
   U141 : AOI221_X1 port map( B1 => n268, B2 => n408, C1 => n270, C2 => n419, A
                           => n420, ZN => n413);
   U142 : OAI22_X1 port map( A1 => n410, A2 => n265, B1 => n421, B2 => n262, ZN
                           => n420);
   U143 : INV_X1 port map( A => n384, ZN => n408);
   U144 : OAI211_X1 port map( C1 => n378, C2 => n368, A => n379, B => n422, ZN 
                           => n384);
   U145 : AOI222_X1 port map( A1 => R(16), A2 => n299, B1 => n338, B2 => R(0), 
                           C1 => R(8), C2 => n298, ZN => n422);
   U147 : MUX2_X1 port map( A => n425, B => n418, S => Offset(0), Z => 
                           Shift_OUT(16));
   U148 : AOI221_X1 port map( B1 => n259, B2 => n415, C1 => n257, C2 => n426, A
                           => n427, ZN => n418);
   U149 : OAI22_X1 port map( A1 => n390, A2 => n251, B1 => n399, B2 => n253, ZN
                           => n427);
   U150 : INV_X1 port map( A => n414, ZN => n399);
   U151 : OAI211_X1 port map( C1 => n378, C2 => n428, A => n497, B => n430, ZN 
                           => n390);
   U152 : MUX2_X1 port map( A => n431, B => n425, S => Offset(0), Z => 
                           Shift_OUT(15));
   U153 : AOI221_X1 port map( B1 => n268, B2 => n419, C1 => n270, C2 => n432, A
                           => n433, ZN => n425);
   U154 : OAI22_X1 port map( A1 => n421, A2 => n265, B1 => n434, B2 => n262, ZN
                           => n433);
   U155 : INV_X1 port map( A => n395, ZN => n419);
   U156 : OAI211_X1 port map( C1 => n328, C2 => n385, A => n497, B => n435, ZN 
                           => n395);
   U157 : AOI222_X1 port map( A1 => R(14), A2 => n299, B1 => R(6), B2 => n298, 
                           C1 => R(22), C2 => n325, ZN => n435);
   U158 : MUX2_X1 port map( A => n436, B => n431, S => Offset(0), Z => 
                           Shift_OUT(14));
   U159 : INV_X1 port map( A => n437, ZN => n431);
   U160 : OAI221_X1 port map( B1 => n265, B2 => n438, C1 => n262, C2 => n252, A
                           => n439, ZN => n437);
   U161 : AOI22_X1 port map( A1 => n414, A2 => n268, B1 => n415, B2 => n270, ZN
                           => n439);
   U162 : AOI211_X1 port map( C1 => n325, C2 => R(21), A => n424, B => n440, ZN
                           => n414);
   U163 : OAI222_X1 port map( A1 => n317, A2 => n328, B1 => n318, B2 => n314, 
                           C1 => n319, C2 => n316, ZN => n440);
   U164 : INV_X1 port map( A => R(5), ZN => n318);
   U165 : MUX2_X1 port map( A => n441, B => n436, S => Offset(0), Z => 
                           Shift_OUT(13));
   U166 : AOI221_X1 port map( B1 => n257, B2 => n267, C1 => n268, C2 => n432, A
                           => n442, ZN => n436);
   U167 : OAI22_X1 port map( A1 => n421, A2 => n253, B1 => n265, B2 => n434, ZN
                           => n442);
   U168 : INV_X1 port map( A => n410, ZN => n432);
   U169 : OAI211_X1 port map( C1 => n378, C2 => n336, A => n497, B => n443, ZN 
                           => n410);
   U170 : AOI222_X1 port map( A1 => R(28), A2 => n423, B1 => R(4), B2 => n298, 
                           C1 => R(12), C2 => n299, ZN => n443);
   U171 : MUX2_X1 port map( A => n444, B => n441, S => Offset(0), Z => 
                           Shift_OUT(12));
   U172 : INV_X1 port map( A => n445, ZN => n441);
   U173 : OAI221_X1 port map( B1 => n265, B2 => n252, C1 => n262, C2 => n254, A
                           => n446, ZN => n445);
   U174 : AOI22_X1 port map( A1 => n415, A2 => n268, B1 => n426, B2 => n270, ZN
                           => n446);
   U175 : INV_X1 port map( A => n447, ZN => n415);
   U176 : OAI211_X1 port map( C1 => n328, C2 => n346, A => n497, B => n448, ZN 
                           => n447);
   U177 : AOI222_X1 port map( A1 => R(11), A2 => n299, B1 => R(3), B2 => n298, 
                           C1 => R(19), C2 => n325, ZN => n448);
   U178 : MUX2_X1 port map( A => n449, B => n444, S => Offset(0), Z => 
                           Shift_OUT(11));
   U179 : AOI221_X1 port map( B1 => n267, B2 => n259, C1 => n257, C2 => n269, A
                           => n450, ZN => n444);
   U180 : OAI22_X1 port map( A1 => n421, A2 => n251, B1 => n253, B2 => n434, ZN
                           => n450);
   U181 : INV_X1 port map( A => n451, ZN => n421);
   U182 : AOI211_X1 port map( C1 => R(18), C2 => n325, A => n424, B => n452, ZN
                           => n451);
   U183 : OAI222_X1 port map( A1 => n411, A2 => n328, B1 => n314, B2 => n355, 
                           C1 => n354, C2 => n316, ZN => n452);
   U184 : INV_X1 port map( A => n298, ZN => n314);
   U185 : INV_X1 port map( A => n496, ZN => n424);
   U186 : MUX2_X1 port map( A => n248, B => n449, S => Offset(0), Z => 
                           Shift_OUT(10));
   U187 : INV_X1 port map( A => n453, ZN => n449);
   U188 : OAI221_X1 port map( B1 => n253, B2 => n252, C1 => n265, C2 => n254, A
                           => n454, ZN => n453);
   U189 : AOI22_X1 port map( A1 => n258, A2 => n257, B1 => n426, B2 => n268, ZN
                           => n454);
   U190 : INV_X1 port map( A => n438, ZN => n426);
   U191 : OAI211_X1 port map( C1 => n378, C2 => n327, A => n497, B => n455, ZN 
                           => n438);
   U192 : AOI222_X1 port map( A1 => R(25), A2 => n423, B1 => R(1), B2 => n298, 
                           C1 => R(9), C2 => n299, ZN => n455);
   U193 : AOI221_X1 port map( B1 => n423, B2 => R(19), C1 => n325, C2 => R(11),
                           A => n456, ZN => n258);
   U194 : OAI221_X1 port map( B1 => n346, B2 => n457, C1 => n458, C2 => n316, A
                           => n330, ZN => n456);
   U195 : INV_X1 port map( A => R(3), ZN => n458);
   U196 : OAI221_X1 port map( B1 => n328, B2 => n315, C1 => n378, C2 => n319, A
                           => n459, ZN => n254);
   U197 : AOI221_X1 port map( B1 => R(29), B2 => n324, C1 => R(5), C2 => n299, 
                           A => n494, ZN => n459);
   U198 : INV_X1 port map( A => R(21), ZN => n315);
   U199 : INV_X1 port map( A => n259, ZN => n265);
   U200 : OAI221_X1 port map( B1 => n377, B2 => n457, C1 => n378, C2 => n461, A
                           => n462, ZN => n252);
   U202 : INV_X1 port map( A => R(15), ZN => n461);
   U203 : AOI221_X1 port map( B1 => n270, B2 => n267, C1 => n259, C2 => n269, A
                           => n463, ZN => n248);
   U204 : OAI22_X1 port map( A1 => n262, A2 => n264, B1 => n251, B2 => n434, ZN
                           => n463);
   U205 : OAI211_X1 port map( C1 => n378, C2 => n367, A => n497, B => n464, ZN 
                           => n434);
   U206 : AOI222_X1 port map( A1 => R(24), A2 => n423, B1 => R(0), B2 => n298, 
                           C1 => R(8), C2 => n299, ZN => n464);
   U208 : INV_X1 port map( A => R(16), ZN => n367);
   U209 : INV_X1 port map( A => n268, ZN => n251);
   U210 : OAI221_X1 port map( B1 => n457, B2 => n411, C1 => n378, C2 => n354, A
                           => n465, ZN => n264);
   U211 : AOI221_X1 port map( B1 => R(18), B2 => n423, C1 => R(2), C2 => n299, 
                           A => n494, ZN => n465);
   U213 : INV_X1 port map( A => R(26), ZN => n411);
   U214 : AOI221_X1 port map( B1 => n423, B2 => R(20), C1 => n325, C2 => R(12),
                           A => n466, ZN => n269);
   U215 : OAI221_X1 port map( B1 => n335, B2 => n457, C1 => n467, C2 => n316, A
                           => n330, ZN => n466);
   U216 : INV_X1 port map( A => R(4), ZN => n467);
   U217 : AOI221_X1 port map( B1 => n423, B2 => R(22), C1 => n325, C2 => R(14),
                           A => n468, ZN => n267);
   U218 : OAI221_X1 port map( B1 => n385, B2 => n457, C1 => n301, C2 => n316, A
                           => n330, ZN => n468);
   U220 : INV_X1 port map( A => n305, ZN => n340);
   U221 : NAND2_X1 port map( A1 => R(31), A2 => Conf(0), ZN => n305);
   U222 : INV_X1 port map( A => n299, ZN => n316);
   U223 : INV_X1 port map( A => n470, ZN => n371);
   U224 : INV_X1 port map( A => R(30), ZN => n385);
   U225 : MUX2_X1 port map( A => n471, B => n401, S => Offset(0), Z => 
                           Shift_OUT(0));
   U226 : AOI221_X1 port map( B1 => n270, B2 => n281, C1 => n268, C2 => n275, A
                           => n472, ZN => n401);
   U227 : INV_X1 port map( A => n473, ZN => n472);
   U228 : AOI21_X1 port map( B1 => n321, B2 => n259, A => n474, ZN => n473);
   U229 : AOI211_X1 port map( C1 => R(9), C2 => n423, A => n475, B => n262, ZN 
                           => n474);
   U230 : OAI222_X1 port map( A1 => n378, A2 => n329, B1 => n457, B2 => n327, 
                           C1 => n476, C2 => n361, ZN => n475);
   U231 : INV_X1 port map( A => R(25), ZN => n361);
   U232 : INV_X1 port map( A => R(17), ZN => n327);
   U233 : INV_X1 port map( A => R(1), ZN => n329);
   U234 : AOI221_X1 port map( B1 => n325, B2 => R(3), C1 => n423, C2 => R(11), 
                           A => n477, ZN => n321);
   U235 : OAI22_X1 port map( A1 => n347, A2 => n457, B1 => n346, B2 => n476, ZN
                           => n477);
   U236 : INV_X1 port map( A => R(27), ZN => n346);
   U237 : INV_X1 port map( A => R(19), ZN => n347);
   U238 : AOI221_X1 port map( B1 => n325, B2 => R(7), C1 => n423, C2 => R(15), 
                           A => n478, ZN => n275);
   U239 : OAI22_X1 port map( A1 => n428, A2 => n457, B1 => n476, B2 => n377, ZN
                           => n478);
   U240 : INV_X1 port map( A => R(31), ZN => n377);
   U241 : INV_X1 port map( A => R(23), ZN => n428);
   U242 : OAI22_X1 port map( A1 => n319, A2 => n328, B1 => n317, B2 => n476, ZN
                           => n479);
   U243 : INV_X1 port map( A => R(29), ZN => n317);
   U244 : INV_X1 port map( A => R(13), ZN => n319);
   U245 : OAI221_X1 port map( B1 => n480, B2 => n262, C1 => n287, C2 => n253, A
                           => n481, ZN => n471);
   U246 : AOI22_X1 port map( A1 => n259, A2 => n403, B1 => n268, B2 => n288, ZN
                           => n481);
   U247 : OAI221_X1 port map( B1 => n328, B2 => n303, C1 => n378, C2 => n301, A
                           => n482, ZN => n288);
   U248 : AOI22_X1 port map( A1 => R(22), A2 => n324, B1 => R(30), B2 => n469, 
                           ZN => n482);
   U249 : INV_X1 port map( A => R(6), ZN => n301);
   U250 : INV_X1 port map( A => R(14), ZN => n303);
   U251 : OAI221_X1 port map( B1 => n355, B2 => n378, C1 => n328, C2 => n354, A
                           => n485, ZN => n403);
   U252 : AOI22_X1 port map( A1 => n324, A2 => R(18), B1 => R(26), B2 => n469, 
                           ZN => n485);
   U253 : INV_X1 port map( A => R(10), ZN => n354);
   U254 : INV_X1 port map( A => n423, ZN => n328);
   U255 : INV_X1 port map( A => R(2), ZN => n355);
   U256 : INV_X1 port map( A => n270, ZN => n253);
   U257 : INV_X1 port map( A => n486, ZN => n484);
   U258 : AOI221_X1 port map( B1 => n325, B2 => R(4), C1 => n423, C2 => R(12), 
                           A => n488, ZN => n287);
   U259 : OAI22_X1 port map( A1 => n336, A2 => n457, B1 => n335, B2 => n476, ZN
                           => n488);
   U260 : INV_X1 port map( A => R(28), ZN => n335);
   U261 : INV_X1 port map( A => n324, ZN => n457);
   U262 : INV_X1 port map( A => R(20), ZN => n336);
   U263 : INV_X1 port map( A => n257, ZN => n262);
   U264 : INV_X1 port map( A => n483, ZN => n487);
   U265 : NAND2_X1 port map( A1 => n489, A2 => n490, ZN => n483);
   U266 : MUX2_X1 port map( A => n470, B => n491, S => Offset(1), Z => n489);
   U267 : NAND2_X1 port map( A1 => Offset(0), A2 => n470, ZN => n491);
   U268 : XNOR2_X1 port map( A => n492, B => Offset(2), ZN => n486);
   U269 : NAND2_X1 port map( A1 => n470, A2 => n490, ZN => n492);
   U270 : OR2_X1 port map( A1 => Offset(0), A2 => Offset(1), ZN => n490);
   U271 : AOI221_X1 port map( B1 => R(8), B2 => n423, C1 => R(16), C2 => n324, 
                           A => n493, ZN => n480);
   U272 : OAI22_X1 port map( A1 => n476, A2 => n368, B1 => n378, B2 => n406, ZN
                           => n493);
   U273 : INV_X1 port map( A => R(0), ZN => n406);
   U274 : INV_X1 port map( A => n325, ZN => n378);
   U275 : INV_X1 port map( A => R(24), ZN => n368);
   U276 : INV_X1 port map( A => n469, ZN => n476);
   U277 : NOR3_X1 port map( A1 => n370, A2 => n470, A3 => n372, ZN => n469);
   U278 : INV_X1 port map( A => Offset(4), ZN => n372);
   U279 : INV_X1 port map( A => Offset(3), ZN => n370);
   U280 : NOR2_X1 port map( A1 => Conf(0), A2 => Conf(1), ZN => n470);
   U65 : OAI221_X1 port map( B1 => Offset(4), B2 => Offset(3), C1 => Conf(0), 
                           C2 => Conf(1), A => n340, ZN => n379);
   U71 : AND2_X2 port map( A1 => n469, A2 => n340, ZN => n494);
   U85 : INV_X4 port map( A => n494, ZN => n330);
   U91 : AOI221_X4 port map( B1 => n338, B2 => R(9), C1 => n339, C2 => R(1), A 
                           => n340, ZN => n362);
   U146 : AOI21_X1 port map( B1 => n340, B2 => n324, A => n494, ZN => n429);
   U201 : INV_X1 port map( A => n429, ZN => n495);
   U207 : INV_X1 port map( A => n495, ZN => n496);
   U212 : INV_X1 port map( A => n495, ZN => n497);
   U219 : AOI221_X4 port map( B1 => n338, B2 => R(12), C1 => n339, C2 => R(4), 
                           A => n340, ZN => n337);
   U281 : AOI221_X4 port map( B1 => n338, B2 => R(11), C1 => n339, C2 => R(3), 
                           A => n340, ZN => n348);
   U282 : AOI221_X4 port map( B1 => n338, B2 => R(8), C1 => n339, C2 => R(0), A
                           => n340, ZN => n369);
   U283 : AOI221_X4 port map( B1 => R(23), B2 => n423, C1 => R(7), C2 => n299, 
                           A => n494, ZN => n462);

end SYN_Struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ComparatorUnit is

   port( A_MSB, B_MSB : in std_logic;  SUBIN : in std_logic_vector (31 downto 
         0);  COUT, SIGN_UNSIGN : in std_logic;  OP : in std_logic_vector (0 to
         2);  CU_OUT : out std_logic_vector (31 downto 0));

end ComparatorUnit;

architecture SYN_Beh of ComparatorUnit is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X2
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, CU_OUT_0_port, net123593, n39, n50, n41, n40, 
      net124999, net124998, net124924, net124922, net125054, net125029, 
      net125028, net125025, net125024, net125023, net125022, net125021, 
      net124992, net124989, net124976, net124927, n34, n32, n30, net125020, 
      net124983, net124980, net124995, net125095, net125050, net124982, 
      net124967, net124965, net124964, net124963, net124925, net123651, 
      net123650, net123620, net123618, n36, n31, net125090, net125007, 
      net125006, net125005, net125004, net125002, net124994, net124993, n53, 
      n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68
      , n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81 : 
      std_logic;

begin
   CU_OUT <= ( X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      CU_OUT_0_port );
   
   X_Logic0_port <= '0';
   U67 : INV_X1 port map( A => A_MSB, ZN => n40);
   U76 : XOR2_X1 port map( A => B_MSB, B => A_MSB, Z => n50);
   U75 : AND2_X1 port map( A1 => SIGN_UNSIGN, A2 => n50, ZN => n41);
   syn379 : INV_X2 port map( A => n40, ZN => net124999);
   syn369 : NAND3_X1 port map( A1 => n80, A2 => net125028, A3 => net124989, ZN 
                           => n81);
   syn362 : NOR2_X2 port map( A1 => net125022, A2 => net125023, ZN => n79);
   U63 : OAI21_X1 port map( B1 => net123593, B2 => n39, A => n34, ZN => n30);
   syn489 : NAND2_X2 port map( A1 => OP(2), A2 => net125029, ZN => net124922);
   syn361 : NAND3_X1 port map( A1 => net125024, A2 => net125025, A3 => n71, ZN 
                           => net125023);
   U64 : INV_X1 port map( A => OP(1), ZN => n34);
   syn92 : INV_X2 port map( A => OP(2), ZN => net124925);
   U58 : AOI22_X1 port map( A1 => n30, A2 => OP(0), B1 => n31, B2 => n32, ZN =>
                           CU_OUT_0_port);
   syn309 : NAND3_X1 port map( A1 => net125004, A2 => net125005, A3 => 
                           net125007, ZN => net125006);
   syn294 : NOR2_X2 port map( A1 => n41, A2 => SUBIN(1), ZN => n60);
   syn411 : INV_X2 port map( A => SUBIN(15), ZN => n62);
   syn312 : NOR2_X2 port map( A1 => SUBIN(0), A2 => SUBIN(10), ZN => n63);
   syn316 : NOR2_X2 port map( A1 => SUBIN(4), A2 => SUBIN(9), ZN => n64);
   syn319 : NAND3_X1 port map( A1 => n63, A2 => n66, A3 => n64, ZN => n65);
   syn320 : NOR2_X2 port map( A1 => SUBIN(8), A2 => SUBIN(5), ZN => n67);
   syn324 : NOR2_X2 port map( A1 => SUBIN(6), A2 => SUBIN(2), ZN => n68);
   syn327 : NAND3_X1 port map( A1 => n67, A2 => n70, A3 => n68, ZN => n69);
   U59 : NAND2_X1 port map( A1 => net124983, A2 => net124964, ZN => n74);
   U60 : OR2_X1 port map( A1 => SUBIN(25), A2 => SUBIN(26), ZN => net124983);
   U61 : CLKBUF_X1 port map( A => n72, Z => n53);
   U62 : AND4_X1 port map( A1 => n58, A2 => n59, A3 => net125090, A4 => 
                           net124993, ZN => n54);
   U65 : NAND2_X1 port map( A1 => net125021, A2 => n53, ZN => net125022);
   U66 : OAI21_X1 port map( B1 => net125029, B2 => n34, A => OP(2), ZN => 
                           net124976);
   U68 : AND4_X1 port map( A1 => net124989, A2 => n72, A3 => n55, A4 => n56, ZN
                           => net125020);
   U69 : INV_X1 port map( A => SUBIN(25), ZN => n55);
   U70 : INV_X1 port map( A => SUBIN(26), ZN => n56);
   U71 : OAI211_X1 port map( C1 => net125095, C2 => net123650, A => n73, B => 
                           n74, ZN => net124965);
   U72 : NOR2_X1 port map( A1 => net124963, A2 => net124967, ZN => net123593);
   U73 : NOR2_X1 port map( A1 => n81, A2 => net124992, ZN => n78);
   U74 : OAI211_X1 port map( C1 => n54, C2 => net123650, A => n57, B => 
                           net123620, ZN => n31);
   U77 : INV_X1 port map( A => net124965, ZN => n57);
   U78 : NAND4_X1 port map( A1 => n58, A2 => n59, A3 => net124994, A4 => 
                           net124993, ZN => net124963);
   U79 : INV_X1 port map( A => net124995, ZN => n58);
   U80 : INV_X1 port map( A => OP(2), ZN => n59);
   U81 : NOR2_X1 port map( A1 => net125002, A2 => net125006, ZN => net124994);
   U82 : NOR2_X1 port map( A1 => n65, A2 => n69, ZN => net124993);
   U83 : NAND2_X1 port map( A1 => net125090, A2 => net124993, ZN => net124992);
   U84 : INV_X1 port map( A => SUBIN(7), ZN => n70);
   U85 : INV_X1 port map( A => SUBIN(11), ZN => n66);
   U86 : NAND3_X1 port map( A1 => n60, A2 => n62, A3 => n61, ZN => net125002);
   U87 : NOR2_X1 port map( A1 => net125002, A2 => net125006, ZN => net125090);
   U88 : NOR2_X1 port map( A1 => SUBIN(14), A2 => SUBIN(13), ZN => n61);
   U89 : INV_X1 port map( A => SUBIN(12), ZN => net125007);
   U90 : NOR2_X1 port map( A1 => SUBIN(17), A2 => SUBIN(16), ZN => net125005);
   U91 : NOR2_X1 port map( A1 => SUBIN(18), A2 => SUBIN(19), ZN => net125004);
   U92 : MUX2_X2 port map( A => net124998, B => net124999, S => n41, Z => 
                           net124924);
   U93 : NAND2_X1 port map( A1 => n36, A2 => OP(1), ZN => net123620);
   U94 : AND2_X1 port map( A1 => net125050, A2 => n75, ZN => n73);
   U95 : NAND2_X1 port map( A1 => net124964, A2 => SUBIN(27), ZN => n75);
   U96 : INV_X1 port map( A => net123650, ZN => net124964);
   U97 : OR2_X1 port map( A1 => n72, A2 => net123650, ZN => net125050);
   U98 : INV_X1 port map( A => SUBIN(24), ZN => n72);
   U99 : NAND2_X1 port map( A1 => net124924, A2 => net124925, ZN => n36);
   U100 : NAND2_X1 port map( A1 => n36, A2 => net124922, ZN => n39);
   U101 : INV_X1 port map( A => OP(1), ZN => net123618);
   U102 : OR2_X1 port map( A1 => OP(0), A2 => net123651, ZN => net123650);
   U103 : INV_X1 port map( A => net123618, ZN => net123651);
   U104 : AND3_X1 port map( A1 => net124980, A2 => net124982, A3 => n71, ZN => 
                           net125095);
   U105 : NAND2_X1 port map( A1 => net125020, A2 => net125095, ZN => net124967)
                           ;
   U106 : INV_X1 port map( A => SUBIN(23), ZN => n71);
   U107 : NOR2_X1 port map( A1 => SUBIN(29), A2 => SUBIN(28), ZN => net124982);
   U108 : NAND2_X1 port map( A1 => n76, A2 => n77, ZN => net124995);
   U109 : INV_X1 port map( A => net124995, ZN => net125028);
   U110 : NOR2_X1 port map( A1 => SUBIN(22), A2 => SUBIN(21), ZN => n77);
   U111 : NOR2_X2 port map( A1 => SUBIN(20), A2 => SUBIN(3), ZN => n76);
   U112 : NOR2_X1 port map( A1 => SUBIN(30), A2 => SUBIN(31), ZN => net124980);
   U113 : INV_X1 port map( A => SUBIN(27), ZN => net124989);
   U114 : INV_X1 port map( A => net124927, ZN => n32);
   U115 : AOI21_X1 port map( B1 => n78, B2 => n79, A => net124976, ZN => 
                           net124927);
   U116 : INV_X1 port map( A => net124924, ZN => net125029);
   U117 : INV_X1 port map( A => SUBIN(30), ZN => net125025);
   U118 : INV_X1 port map( A => SUBIN(31), ZN => net125024);
   U119 : NOR2_X1 port map( A1 => net125054, A2 => SUBIN(25), ZN => net125021);
   U120 : CLKBUF_X1 port map( A => SUBIN(26), Z => net125054);
   U121 : NOR2_X1 port map( A1 => SUBIN(29), A2 => SUBIN(28), ZN => n80);
   U122 : INV_X1 port map( A => COUT, ZN => net124998);

end SYN_Beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity logicunit is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic_vector 
         (2 downto 0);  LU_OUT : out std_logic_vector (31 downto 0));

end logicunit;

architecture SYN_Behavioral of logicunit is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
      n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, 
      n119, n120, n121, n122, n123, n124, n125, n126, n127, n128 : std_logic;

begin
   
   U1 : MUX2_X1 port map( A => n65, B => n66, S => B(9), Z => LU_OUT(9));
   U2 : MUX2_X1 port map( A => SEL(0), B => SEL(2), S => A(9), Z => n66);
   U3 : AND2_X1 port map( A1 => A(9), A2 => SEL(1), ZN => n65);
   U4 : MUX2_X1 port map( A => n67, B => n68, S => B(8), Z => LU_OUT(8));
   U5 : MUX2_X1 port map( A => SEL(0), B => SEL(2), S => A(8), Z => n68);
   U6 : AND2_X1 port map( A1 => SEL(1), A2 => A(8), ZN => n67);
   U7 : MUX2_X1 port map( A => n69, B => n70, S => B(7), Z => LU_OUT(7));
   U8 : MUX2_X1 port map( A => SEL(0), B => SEL(2), S => A(7), Z => n70);
   U9 : AND2_X1 port map( A1 => SEL(1), A2 => A(7), ZN => n69);
   U10 : MUX2_X1 port map( A => n71, B => n72, S => B(6), Z => LU_OUT(6));
   U11 : MUX2_X1 port map( A => SEL(0), B => SEL(2), S => A(6), Z => n72);
   U12 : AND2_X1 port map( A1 => SEL(1), A2 => A(6), ZN => n71);
   U13 : MUX2_X1 port map( A => n73, B => n74, S => B(5), Z => LU_OUT(5));
   U14 : MUX2_X1 port map( A => SEL(0), B => SEL(2), S => A(5), Z => n74);
   U15 : AND2_X1 port map( A1 => SEL(1), A2 => A(5), ZN => n73);
   U16 : MUX2_X1 port map( A => n75, B => n76, S => B(4), Z => LU_OUT(4));
   U17 : MUX2_X1 port map( A => SEL(0), B => SEL(2), S => A(4), Z => n76);
   U18 : AND2_X1 port map( A1 => SEL(1), A2 => A(4), ZN => n75);
   U19 : MUX2_X1 port map( A => n77, B => n78, S => B(3), Z => LU_OUT(3));
   U20 : MUX2_X1 port map( A => SEL(0), B => SEL(2), S => A(3), Z => n78);
   U21 : AND2_X1 port map( A1 => SEL(1), A2 => A(3), ZN => n77);
   U22 : MUX2_X1 port map( A => n79, B => n80, S => B(31), Z => LU_OUT(31));
   U23 : MUX2_X1 port map( A => SEL(0), B => SEL(2), S => A(31), Z => n80);
   U24 : AND2_X1 port map( A1 => SEL(1), A2 => A(31), ZN => n79);
   U25 : MUX2_X1 port map( A => n81, B => n82, S => B(30), Z => LU_OUT(30));
   U26 : MUX2_X1 port map( A => SEL(0), B => SEL(2), S => A(30), Z => n82);
   U27 : AND2_X1 port map( A1 => SEL(1), A2 => A(30), ZN => n81);
   U28 : MUX2_X1 port map( A => n83, B => n84, S => B(2), Z => LU_OUT(2));
   U29 : MUX2_X1 port map( A => SEL(0), B => SEL(2), S => A(2), Z => n84);
   U30 : AND2_X1 port map( A1 => SEL(1), A2 => A(2), ZN => n83);
   U31 : MUX2_X1 port map( A => n85, B => n86, S => B(29), Z => LU_OUT(29));
   U32 : MUX2_X1 port map( A => SEL(0), B => SEL(2), S => A(29), Z => n86);
   U33 : AND2_X1 port map( A1 => SEL(1), A2 => A(29), ZN => n85);
   U34 : MUX2_X1 port map( A => n87, B => n88, S => B(28), Z => LU_OUT(28));
   U35 : MUX2_X1 port map( A => SEL(0), B => SEL(2), S => A(28), Z => n88);
   U36 : AND2_X1 port map( A1 => SEL(1), A2 => A(28), ZN => n87);
   U37 : MUX2_X1 port map( A => n89, B => n90, S => B(27), Z => LU_OUT(27));
   U38 : MUX2_X1 port map( A => SEL(0), B => SEL(2), S => A(27), Z => n90);
   U39 : AND2_X1 port map( A1 => SEL(1), A2 => A(27), ZN => n89);
   U40 : MUX2_X1 port map( A => n91, B => n92, S => B(26), Z => LU_OUT(26));
   U41 : MUX2_X1 port map( A => SEL(0), B => SEL(2), S => A(26), Z => n92);
   U42 : AND2_X1 port map( A1 => SEL(1), A2 => A(26), ZN => n91);
   U43 : MUX2_X1 port map( A => n93, B => n94, S => B(25), Z => LU_OUT(25));
   U44 : MUX2_X1 port map( A => SEL(0), B => SEL(2), S => A(25), Z => n94);
   U45 : AND2_X1 port map( A1 => SEL(1), A2 => A(25), ZN => n93);
   U46 : MUX2_X1 port map( A => n95, B => n96, S => B(24), Z => LU_OUT(24));
   U47 : MUX2_X1 port map( A => SEL(0), B => SEL(2), S => A(24), Z => n96);
   U48 : AND2_X1 port map( A1 => SEL(1), A2 => A(24), ZN => n95);
   U49 : MUX2_X1 port map( A => n97, B => n98, S => B(23), Z => LU_OUT(23));
   U50 : MUX2_X1 port map( A => SEL(0), B => SEL(2), S => A(23), Z => n98);
   U51 : AND2_X1 port map( A1 => SEL(1), A2 => A(23), ZN => n97);
   U52 : MUX2_X1 port map( A => n99, B => n100, S => B(22), Z => LU_OUT(22));
   U53 : MUX2_X1 port map( A => SEL(0), B => SEL(2), S => A(22), Z => n100);
   U54 : AND2_X1 port map( A1 => SEL(1), A2 => A(22), ZN => n99);
   U55 : MUX2_X1 port map( A => n101, B => n102, S => B(21), Z => LU_OUT(21));
   U56 : MUX2_X1 port map( A => SEL(0), B => SEL(2), S => A(21), Z => n102);
   U57 : AND2_X1 port map( A1 => SEL(1), A2 => A(21), ZN => n101);
   U58 : MUX2_X1 port map( A => n103, B => n104, S => B(20), Z => LU_OUT(20));
   U59 : MUX2_X1 port map( A => SEL(0), B => SEL(2), S => A(20), Z => n104);
   U60 : AND2_X1 port map( A1 => SEL(1), A2 => A(20), ZN => n103);
   U61 : MUX2_X1 port map( A => n105, B => n106, S => B(1), Z => LU_OUT(1));
   U62 : MUX2_X1 port map( A => SEL(0), B => SEL(2), S => A(1), Z => n106);
   U63 : AND2_X1 port map( A1 => SEL(1), A2 => A(1), ZN => n105);
   U64 : MUX2_X1 port map( A => n107, B => n108, S => B(19), Z => LU_OUT(19));
   U65 : MUX2_X1 port map( A => SEL(0), B => SEL(2), S => A(19), Z => n108);
   U66 : AND2_X1 port map( A1 => SEL(1), A2 => A(19), ZN => n107);
   U67 : MUX2_X1 port map( A => n109, B => n110, S => B(18), Z => LU_OUT(18));
   U68 : MUX2_X1 port map( A => SEL(0), B => SEL(2), S => A(18), Z => n110);
   U69 : AND2_X1 port map( A1 => SEL(1), A2 => A(18), ZN => n109);
   U70 : MUX2_X1 port map( A => n111, B => n112, S => B(17), Z => LU_OUT(17));
   U71 : MUX2_X1 port map( A => SEL(0), B => SEL(2), S => A(17), Z => n112);
   U72 : AND2_X1 port map( A1 => SEL(1), A2 => A(17), ZN => n111);
   U73 : MUX2_X1 port map( A => n113, B => n114, S => B(16), Z => LU_OUT(16));
   U74 : MUX2_X1 port map( A => SEL(0), B => SEL(2), S => A(16), Z => n114);
   U75 : AND2_X1 port map( A1 => SEL(1), A2 => A(16), ZN => n113);
   U76 : MUX2_X1 port map( A => n115, B => n116, S => B(15), Z => LU_OUT(15));
   U77 : MUX2_X1 port map( A => SEL(0), B => SEL(2), S => A(15), Z => n116);
   U78 : AND2_X1 port map( A1 => SEL(1), A2 => A(15), ZN => n115);
   U79 : MUX2_X1 port map( A => n117, B => n118, S => B(14), Z => LU_OUT(14));
   U80 : MUX2_X1 port map( A => SEL(0), B => SEL(2), S => A(14), Z => n118);
   U81 : AND2_X1 port map( A1 => SEL(1), A2 => A(14), ZN => n117);
   U82 : MUX2_X1 port map( A => n119, B => n120, S => B(13), Z => LU_OUT(13));
   U83 : MUX2_X1 port map( A => SEL(0), B => SEL(2), S => A(13), Z => n120);
   U84 : AND2_X1 port map( A1 => SEL(1), A2 => A(13), ZN => n119);
   U85 : MUX2_X1 port map( A => n121, B => n122, S => B(12), Z => LU_OUT(12));
   U86 : MUX2_X1 port map( A => SEL(0), B => SEL(2), S => A(12), Z => n122);
   U87 : AND2_X1 port map( A1 => SEL(1), A2 => A(12), ZN => n121);
   U88 : MUX2_X1 port map( A => n123, B => n124, S => B(11), Z => LU_OUT(11));
   U89 : MUX2_X1 port map( A => SEL(0), B => SEL(2), S => A(11), Z => n124);
   U90 : AND2_X1 port map( A1 => SEL(1), A2 => A(11), ZN => n123);
   U91 : MUX2_X1 port map( A => n125, B => n126, S => B(10), Z => LU_OUT(10));
   U92 : MUX2_X1 port map( A => SEL(0), B => SEL(2), S => A(10), Z => n126);
   U93 : AND2_X1 port map( A1 => SEL(1), A2 => A(10), ZN => n125);
   U94 : MUX2_X1 port map( A => n127, B => n128, S => B(0), Z => LU_OUT(0));
   U95 : MUX2_X1 port map( A => SEL(0), B => SEL(2), S => A(0), Z => n128);
   U96 : AND2_X1 port map( A1 => SEL(1), A2 => A(0), ZN => n127);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity sumgen_N_blocks8 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector (7
         downto 0);  S : out std_logic_vector (31 downto 0));

end sumgen_N_blocks8;

architecture SYN_STRUCTURAL of sumgen_N_blocks8 is

   component CSB_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSB_2
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSB_3
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSB_4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSB_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSB_6
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSB_7
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSB_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   
   CSBI_0 : CSB_0 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => Ci(0), S(3) => S(3), S(2) => S(2), 
                           S(1) => S(1), S(0) => S(0));
   CSBI_1 : CSB_7 port map( A(3) => A(7), A(2) => A(6), A(1) => A(5), A(0) => 
                           A(4), B(3) => B(7), B(2) => B(6), B(1) => B(5), B(0)
                           => B(4), Ci => Ci(1), S(3) => S(7), S(2) => S(6), 
                           S(1) => S(5), S(0) => S(4));
   CSBI_2 : CSB_6 port map( A(3) => A(11), A(2) => A(10), A(1) => A(9), A(0) =>
                           A(8), B(3) => B(11), B(2) => B(10), B(1) => B(9), 
                           B(0) => B(8), Ci => Ci(2), S(3) => S(11), S(2) => 
                           S(10), S(1) => S(9), S(0) => S(8));
   CSBI_3 : CSB_5 port map( A(3) => A(15), A(2) => A(14), A(1) => A(13), A(0) 
                           => A(12), B(3) => B(15), B(2) => B(14), B(1) => 
                           B(13), B(0) => B(12), Ci => Ci(3), S(3) => S(15), 
                           S(2) => S(14), S(1) => S(13), S(0) => S(12));
   CSBI_4 : CSB_4 port map( A(3) => A(19), A(2) => A(18), A(1) => A(17), A(0) 
                           => A(16), B(3) => B(19), B(2) => B(18), B(1) => 
                           B(17), B(0) => B(16), Ci => Ci(4), S(3) => S(19), 
                           S(2) => S(18), S(1) => S(17), S(0) => S(16));
   CSBI_5 : CSB_3 port map( A(3) => A(23), A(2) => A(22), A(1) => A(21), A(0) 
                           => A(20), B(3) => B(23), B(2) => B(22), B(1) => 
                           B(21), B(0) => B(20), Ci => Ci(5), S(3) => S(23), 
                           S(2) => S(22), S(1) => S(21), S(0) => S(20));
   CSBI_6 : CSB_2 port map( A(3) => A(27), A(2) => A(26), A(1) => A(25), A(0) 
                           => A(24), B(3) => B(27), B(2) => B(26), B(1) => 
                           B(25), B(0) => B(24), Ci => Ci(6), S(3) => S(27), 
                           S(2) => S(26), S(1) => S(25), S(0) => S(24));
   CSBI_7 : CSB_1 port map( A(3) => A(31), A(2) => A(30), A(1) => A(29), A(0) 
                           => A(28), B(3) => B(31), B(2) => B(30), B(1) => 
                           B(29), B(0) => B(28), Ci => Ci(7), S(3) => S(31), 
                           S(2) => S(30), S(1) => S(29), S(0) => S(28));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity STCG_N32_L5 is

   port( A, B : in std_logic_vector (31 downto 0);  cin : in std_logic;  cout :
         out std_logic_vector (7 downto 0));

end STCG_N32_L5;

architecture SYN_struct of STCG_N32_L5 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component G_1
      port( pi, gi, gj : in std_logic;  gout : out std_logic);
   end component;
   
   component G_2
      port( pi, gi, gj : in std_logic;  gout : out std_logic);
   end component;
   
   component G_3
      port( pi, gi, gj : in std_logic;  gout : out std_logic);
   end component;
   
   component G_4
      port( pi, gi, gj : in std_logic;  gout : out std_logic);
   end component;
   
   component PG_1
      port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PG_2
      port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component G_5
      port( pi, gi, gj : in std_logic;  gout : out std_logic);
   end component;
   
   component G_6
      port( pi, gi, gj : in std_logic;  gout : out std_logic);
   end component;
   
   component PG_3
      port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PG_4
      port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PG_5
      port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component G_7
      port( pi, gi, gj : in std_logic;  gout : out std_logic);
   end component;
   
   component PG_6
      port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PG_7
      port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PG_8
      port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PG_9
      port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PG_10
      port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PG_11
      port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PG_12
      port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component G_8
      port( pi, gi, gj : in std_logic;  gout : out std_logic);
   end component;
   
   component PG_13
      port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PG_14
      port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PG_15
      port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PG_16
      port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PG_17
      port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PG_18
      port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PG_19
      port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PG_20
      port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PG_21
      port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PG_22
      port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PG_23
      port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PG_24
      port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PG_25
      port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PG_26
      port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component PG_0
      port( pi, gi, pj, gj : in std_logic;  pout, gout : out std_logic);
   end component;
   
   component G_0
      port( pi, gi, gj : in std_logic;  gout : out std_logic);
   end component;
   
   component prop_gen_1
      port( a, b : in std_logic;  prop, gen : out std_logic);
   end component;
   
   component prop_gen_2
      port( a, b : in std_logic;  prop, gen : out std_logic);
   end component;
   
   component prop_gen_3
      port( a, b : in std_logic;  prop, gen : out std_logic);
   end component;
   
   component prop_gen_4
      port( a, b : in std_logic;  prop, gen : out std_logic);
   end component;
   
   component prop_gen_5
      port( a, b : in std_logic;  prop, gen : out std_logic);
   end component;
   
   component prop_gen_6
      port( a, b : in std_logic;  prop, gen : out std_logic);
   end component;
   
   component prop_gen_7
      port( a, b : in std_logic;  prop, gen : out std_logic);
   end component;
   
   component prop_gen_8
      port( a, b : in std_logic;  prop, gen : out std_logic);
   end component;
   
   component prop_gen_9
      port( a, b : in std_logic;  prop, gen : out std_logic);
   end component;
   
   component prop_gen_10
      port( a, b : in std_logic;  prop, gen : out std_logic);
   end component;
   
   component prop_gen_11
      port( a, b : in std_logic;  prop, gen : out std_logic);
   end component;
   
   component prop_gen_12
      port( a, b : in std_logic;  prop, gen : out std_logic);
   end component;
   
   component prop_gen_13
      port( a, b : in std_logic;  prop, gen : out std_logic);
   end component;
   
   component prop_gen_14
      port( a, b : in std_logic;  prop, gen : out std_logic);
   end component;
   
   component prop_gen_15
      port( a, b : in std_logic;  prop, gen : out std_logic);
   end component;
   
   component prop_gen_16
      port( a, b : in std_logic;  prop, gen : out std_logic);
   end component;
   
   component prop_gen_17
      port( a, b : in std_logic;  prop, gen : out std_logic);
   end component;
   
   component prop_gen_18
      port( a, b : in std_logic;  prop, gen : out std_logic);
   end component;
   
   component prop_gen_19
      port( a, b : in std_logic;  prop, gen : out std_logic);
   end component;
   
   component prop_gen_20
      port( a, b : in std_logic;  prop, gen : out std_logic);
   end component;
   
   component prop_gen_21
      port( a, b : in std_logic;  prop, gen : out std_logic);
   end component;
   
   component prop_gen_22
      port( a, b : in std_logic;  prop, gen : out std_logic);
   end component;
   
   component prop_gen_23
      port( a, b : in std_logic;  prop, gen : out std_logic);
   end component;
   
   component prop_gen_24
      port( a, b : in std_logic;  prop, gen : out std_logic);
   end component;
   
   component prop_gen_25
      port( a, b : in std_logic;  prop, gen : out std_logic);
   end component;
   
   component prop_gen_26
      port( a, b : in std_logic;  prop, gen : out std_logic);
   end component;
   
   component prop_gen_27
      port( a, b : in std_logic;  prop, gen : out std_logic);
   end component;
   
   component prop_gen_28
      port( a, b : in std_logic;  prop, gen : out std_logic);
   end component;
   
   component prop_gen_29
      port( a, b : in std_logic;  prop, gen : out std_logic);
   end component;
   
   component prop_gen_30
      port( a, b : in std_logic;  prop, gen : out std_logic);
   end component;
   
   component prop_gen_0
      port( a, b : in std_logic;  prop, gen : out std_logic);
   end component;
   
   component prop_gen_Cin
      port( a, b, cin : in std_logic;  prop, gen : out std_logic);
   end component;
   
   signal cout_7_port, cout_6_port, cout_5_port, cout_4_port, cout_2_port, 
      gen_0_31_port, gen_0_30_port, gen_0_29_port, gen_0_28_port, gen_0_27_port
      , gen_0_26_port, gen_0_25_port, gen_0_24_port, gen_0_23_port, 
      gen_0_22_port, gen_0_21_port, gen_0_20_port, gen_0_19_port, gen_0_18_port
      , gen_0_17_port, gen_0_16_port, gen_0_15_port, gen_0_14_port, 
      gen_0_13_port, gen_0_12_port, gen_0_11_port, gen_0_10_port, gen_0_9_port,
      gen_0_8_port, gen_0_7_port, gen_0_6_port, gen_0_5_port, gen_0_4_port, 
      gen_0_3_port, gen_0_2_port, gen_0_1_port, gen_0_0_port, gen_1_31_port, 
      gen_1_29_port, gen_1_27_port, gen_1_25_port, gen_1_23_port, gen_1_21_port
      , gen_1_19_port, gen_1_17_port, gen_1_15_port, gen_1_13_port, 
      gen_1_11_port, gen_1_9_port, gen_1_7_port, gen_1_5_port, gen_1_3_port, 
      gen_1_1_port, gen_2_31_port, gen_2_23_port, gen_2_15_port, gen_2_7_port, 
      gen_3_31_port, gen_3_15_port, gen_4_31_port, gen_4_27_port, 
      prop_0_31_port, prop_0_30_port, prop_0_29_port, prop_0_28_port, 
      prop_0_27_port, prop_0_26_port, prop_0_25_port, prop_0_24_port, 
      prop_0_23_port, prop_0_22_port, prop_0_21_port, prop_0_20_port, 
      prop_0_19_port, prop_0_18_port, prop_0_17_port, prop_0_16_port, 
      prop_0_15_port, prop_0_14_port, prop_0_13_port, prop_0_12_port, 
      prop_0_11_port, prop_0_10_port, prop_0_9_port, prop_0_8_port, 
      prop_0_7_port, prop_0_6_port, prop_0_5_port, prop_0_4_port, prop_0_3_port
      , prop_0_2_port, prop_0_1_port, prop_1_31_port, prop_1_29_port, 
      prop_1_27_port, prop_1_25_port, prop_1_23_port, prop_1_21_port, 
      prop_1_19_port, prop_1_17_port, prop_1_15_port, prop_1_13_port, 
      prop_1_11_port, prop_1_9_port, prop_1_7_port, prop_1_5_port, 
      prop_1_3_port, prop_2_31_port, prop_2_27_port, prop_2_23_port, 
      prop_2_19_port, prop_2_15_port, prop_2_11_port, prop_2_7_port, 
      prop_3_31_port, prop_3_23_port, prop_3_15_port, prop_4_31_port, 
      prop_4_27_port, net4519, n1, n22, n23, n24, n37, n26, n36, n29, n30, 
      cout_1_port, n32, n33, cout_0_port, cout_3_port : std_logic;

begin
   cout <= ( cout_7_port, cout_6_port, cout_5_port, cout_4_port, cout_3_port, 
      cout_2_port, cout_1_port, cout_0_port );
   
   prop_gen_Cin0 : prop_gen_Cin port map( a => A(0), b => B(0), cin => cin, 
                           prop => net4519, gen => gen_0_0_port);
   prop_gen_i_1 : prop_gen_0 port map( a => A(1), b => B(1), prop => 
                           prop_0_1_port, gen => gen_0_1_port);
   prop_gen_i_2 : prop_gen_30 port map( a => A(2), b => B(2), prop => 
                           prop_0_2_port, gen => gen_0_2_port);
   prop_gen_i_3 : prop_gen_29 port map( a => A(3), b => B(3), prop => 
                           prop_0_3_port, gen => gen_0_3_port);
   prop_gen_i_4 : prop_gen_28 port map( a => A(4), b => B(4), prop => 
                           prop_0_4_port, gen => gen_0_4_port);
   prop_gen_i_5 : prop_gen_27 port map( a => A(5), b => B(5), prop => 
                           prop_0_5_port, gen => gen_0_5_port);
   prop_gen_i_6 : prop_gen_26 port map( a => A(6), b => B(6), prop => 
                           prop_0_6_port, gen => gen_0_6_port);
   prop_gen_i_7 : prop_gen_25 port map( a => A(7), b => B(7), prop => 
                           prop_0_7_port, gen => gen_0_7_port);
   prop_gen_i_8 : prop_gen_24 port map( a => A(8), b => B(8), prop => 
                           prop_0_8_port, gen => gen_0_8_port);
   prop_gen_i_9 : prop_gen_23 port map( a => A(9), b => B(9), prop => 
                           prop_0_9_port, gen => gen_0_9_port);
   prop_gen_i_10 : prop_gen_22 port map( a => A(10), b => B(10), prop => 
                           prop_0_10_port, gen => gen_0_10_port);
   prop_gen_i_11 : prop_gen_21 port map( a => A(11), b => B(11), prop => 
                           prop_0_11_port, gen => gen_0_11_port);
   prop_gen_i_12 : prop_gen_20 port map( a => A(12), b => B(12), prop => 
                           prop_0_12_port, gen => gen_0_12_port);
   prop_gen_i_13 : prop_gen_19 port map( a => A(13), b => B(13), prop => 
                           prop_0_13_port, gen => gen_0_13_port);
   prop_gen_i_14 : prop_gen_18 port map( a => A(14), b => B(14), prop => 
                           prop_0_14_port, gen => gen_0_14_port);
   prop_gen_i_15 : prop_gen_17 port map( a => A(15), b => B(15), prop => 
                           prop_0_15_port, gen => gen_0_15_port);
   prop_gen_i_16 : prop_gen_16 port map( a => A(16), b => B(16), prop => 
                           prop_0_16_port, gen => gen_0_16_port);
   prop_gen_i_17 : prop_gen_15 port map( a => A(17), b => B(17), prop => 
                           prop_0_17_port, gen => gen_0_17_port);
   prop_gen_i_18 : prop_gen_14 port map( a => A(18), b => B(18), prop => 
                           prop_0_18_port, gen => gen_0_18_port);
   prop_gen_i_19 : prop_gen_13 port map( a => A(19), b => B(19), prop => 
                           prop_0_19_port, gen => gen_0_19_port);
   prop_gen_i_20 : prop_gen_12 port map( a => A(20), b => B(20), prop => 
                           prop_0_20_port, gen => gen_0_20_port);
   prop_gen_i_21 : prop_gen_11 port map( a => A(21), b => B(21), prop => 
                           prop_0_21_port, gen => gen_0_21_port);
   prop_gen_i_22 : prop_gen_10 port map( a => A(22), b => B(22), prop => 
                           prop_0_22_port, gen => gen_0_22_port);
   prop_gen_i_23 : prop_gen_9 port map( a => A(23), b => B(23), prop => 
                           prop_0_23_port, gen => gen_0_23_port);
   prop_gen_i_24 : prop_gen_8 port map( a => A(24), b => B(24), prop => 
                           prop_0_24_port, gen => gen_0_24_port);
   prop_gen_i_25 : prop_gen_7 port map( a => A(25), b => B(25), prop => 
                           prop_0_25_port, gen => gen_0_25_port);
   prop_gen_i_26 : prop_gen_6 port map( a => A(26), b => B(26), prop => 
                           prop_0_26_port, gen => gen_0_26_port);
   prop_gen_i_27 : prop_gen_5 port map( a => A(27), b => B(27), prop => 
                           prop_0_27_port, gen => gen_0_27_port);
   prop_gen_i_28 : prop_gen_4 port map( a => A(28), b => B(28), prop => 
                           prop_0_28_port, gen => gen_0_28_port);
   prop_gen_i_29 : prop_gen_3 port map( a => A(29), b => B(29), prop => 
                           prop_0_29_port, gen => gen_0_29_port);
   prop_gen_i_30 : prop_gen_2 port map( a => A(30), b => B(30), prop => 
                           prop_0_30_port, gen => gen_0_30_port);
   prop_gen_i_31 : prop_gen_1 port map( a => A(31), b => B(31), prop => 
                           prop_0_31_port, gen => gen_0_31_port);
   G_1_1_1 : G_0 port map( pi => prop_0_1_port, gi => gen_0_1_port, gj => 
                           gen_0_0_port, gout => gen_1_1_port);
   PG_0_i_1_3 : PG_0 port map( pi => prop_0_3_port, gi => gen_0_3_port, pj => 
                           prop_0_2_port, gj => gen_0_2_port, pout => 
                           prop_1_3_port, gout => gen_1_3_port);
   PG_0_i_1_5 : PG_26 port map( pi => prop_0_5_port, gi => gen_0_5_port, pj => 
                           prop_0_4_port, gj => gen_0_4_port, pout => 
                           prop_1_5_port, gout => gen_1_5_port);
   PG_0_i_1_7 : PG_25 port map( pi => prop_0_7_port, gi => gen_0_7_port, pj => 
                           prop_0_6_port, gj => gen_0_6_port, pout => 
                           prop_1_7_port, gout => gen_1_7_port);
   PG_0_i_1_9 : PG_24 port map( pi => prop_0_9_port, gi => gen_0_9_port, pj => 
                           prop_0_8_port, gj => gen_0_8_port, pout => 
                           prop_1_9_port, gout => gen_1_9_port);
   PG_0_i_1_11 : PG_23 port map( pi => prop_0_11_port, gi => gen_0_11_port, pj 
                           => prop_0_10_port, gj => gen_0_10_port, pout => 
                           prop_1_11_port, gout => gen_1_11_port);
   PG_0_i_1_13 : PG_22 port map( pi => prop_0_13_port, gi => gen_0_13_port, pj 
                           => prop_0_12_port, gj => gen_0_12_port, pout => 
                           prop_1_13_port, gout => gen_1_13_port);
   PG_0_i_1_15 : PG_21 port map( pi => prop_0_15_port, gi => gen_0_15_port, pj 
                           => prop_0_14_port, gj => gen_0_14_port, pout => 
                           prop_1_15_port, gout => gen_1_15_port);
   PG_0_i_1_17 : PG_20 port map( pi => prop_0_17_port, gi => gen_0_17_port, pj 
                           => prop_0_16_port, gj => gen_0_16_port, pout => 
                           prop_1_17_port, gout => gen_1_17_port);
   PG_0_i_1_19 : PG_19 port map( pi => prop_0_19_port, gi => gen_0_19_port, pj 
                           => prop_0_18_port, gj => gen_0_18_port, pout => 
                           prop_1_19_port, gout => gen_1_19_port);
   PG_0_i_1_21 : PG_18 port map( pi => prop_0_21_port, gi => gen_0_21_port, pj 
                           => prop_0_20_port, gj => gen_0_20_port, pout => 
                           prop_1_21_port, gout => gen_1_21_port);
   PG_0_i_1_23 : PG_17 port map( pi => prop_0_23_port, gi => gen_0_23_port, pj 
                           => prop_0_22_port, gj => gen_0_22_port, pout => 
                           prop_1_23_port, gout => gen_1_23_port);
   PG_0_i_1_25 : PG_16 port map( pi => prop_0_25_port, gi => gen_0_25_port, pj 
                           => prop_0_24_port, gj => gen_0_24_port, pout => 
                           prop_1_25_port, gout => gen_1_25_port);
   PG_0_i_1_27 : PG_15 port map( pi => prop_0_27_port, gi => gen_0_27_port, pj 
                           => prop_0_26_port, gj => gen_0_26_port, pout => 
                           prop_1_27_port, gout => gen_1_27_port);
   PG_0_i_1_29 : PG_14 port map( pi => prop_0_29_port, gi => gen_0_29_port, pj 
                           => prop_0_28_port, gj => gen_0_28_port, pout => 
                           prop_1_29_port, gout => gen_1_29_port);
   PG_0_i_1_31 : PG_13 port map( pi => prop_0_31_port, gi => gen_0_31_port, pj 
                           => prop_0_30_port, gj => gen_0_30_port, pout => 
                           prop_1_31_port, gout => gen_1_31_port);
   G_23_2_3 : G_8 port map( pi => prop_1_3_port, gi => gen_1_3_port, gj => 
                           gen_1_1_port, gout => n37);
   PG_0_i_2_7 : PG_12 port map( pi => prop_1_7_port, gi => gen_1_7_port, pj => 
                           prop_1_5_port, gj => gen_1_5_port, pout => 
                           prop_2_7_port, gout => gen_2_7_port);
   PG_0_i_2_11 : PG_11 port map( pi => prop_1_11_port, gi => gen_1_11_port, pj 
                           => prop_1_9_port, gj => gen_1_9_port, pout => 
                           prop_2_11_port, gout => n24);
   PG_0_i_2_15 : PG_10 port map( pi => prop_1_15_port, gi => gen_1_15_port, pj 
                           => prop_1_13_port, gj => gen_1_13_port, pout => 
                           prop_2_15_port, gout => gen_2_15_port);
   PG_0_i_2_19 : PG_9 port map( pi => prop_1_19_port, gi => gen_1_19_port, pj 
                           => prop_1_17_port, gj => gen_1_17_port, pout => 
                           prop_2_19_port, gout => n22);
   PG_0_i_2_23 : PG_8 port map( pi => prop_1_23_port, gi => gen_1_23_port, pj 
                           => prop_1_21_port, gj => gen_1_21_port, pout => 
                           prop_2_23_port, gout => gen_2_23_port);
   PG_0_i_2_27 : PG_7 port map( pi => prop_1_27_port, gi => gen_1_27_port, pj 
                           => prop_1_25_port, gj => gen_1_25_port, pout => 
                           prop_2_27_port, gout => n1);
   PG_0_i_2_31 : PG_6 port map( pi => prop_1_31_port, gi => gen_1_31_port, pj 
                           => prop_1_29_port, gj => gen_1_29_port, pout => 
                           prop_2_31_port, gout => gen_2_31_port);
   G_23_3_7 : G_7 port map( pi => prop_2_7_port, gi => gen_2_7_port, gj => n37,
                           gout => n26);
   PG_0_i_3_15 : PG_5 port map( pi => prop_2_15_port, gi => gen_2_15_port, pj 
                           => prop_2_11_port, gj => n24, pout => prop_3_15_port
                           , gout => gen_3_15_port);
   PG_0_i_3_23 : PG_4 port map( pi => prop_2_23_port, gi => gen_2_23_port, pj 
                           => prop_2_19_port, gj => n22, pout => prop_3_23_port
                           , gout => n23);
   PG_0_i_3_31 : PG_3 port map( pi => prop_2_31_port, gi => gen_2_31_port, pj 
                           => prop_2_27_port, gj => n1, pout => prop_3_31_port,
                           gout => gen_3_31_port);
   G_jk_4_15_1_0 : G_6 port map( pi => prop_3_15_port, gi => gen_3_15_port, gj 
                           => n26, gout => n36);
   G_jk1_4_15_1_0 : G_5 port map( pi => prop_2_11_port, gi => n30, gj => n33, 
                           gout => cout_2_port);
   PG_jk_4_31_1_0 : PG_2 port map( pi => prop_3_31_port, gi => gen_3_31_port, 
                           pj => prop_3_23_port, gj => n29, pout => 
                           prop_4_31_port, gout => gen_4_31_port);
   PG_jk1_4_31_1_0 : PG_1 port map( pi => prop_2_27_port, gi => n1, pj => 
                           prop_3_23_port, gj => n23, pout => prop_4_27_port, 
                           gout => gen_4_27_port);
   G_jk_5_31_2_0 : G_4 port map( pi => prop_4_31_port, gi => gen_4_31_port, gj 
                           => n32, gout => cout_7_port);
   G_jk_5_31_2_1 : G_3 port map( pi => prop_4_27_port, gi => gen_4_27_port, gj 
                           => n36, gout => cout_6_port);
   G_jk_5_31_1_0 : G_2 port map( pi => prop_3_23_port, gi => n29, gj => n36, 
                           gout => cout_5_port);
   G_jk1_5_31_1_0 : G_1 port map( pi => prop_2_19_port, gi => n22, gj => n36, 
                           gout => cout_4_port);
   U1 : CLKBUF_X1 port map( A => n23, Z => n29);
   U2 : BUF_X2 port map( A => n36, Z => cout_3_port);
   U3 : CLKBUF_X1 port map( A => n24, Z => n30);
   U4 : BUF_X1 port map( A => n33, Z => cout_1_port);
   U5 : CLKBUF_X1 port map( A => n26, Z => n33);
   U6 : CLKBUF_X1 port map( A => cout_3_port, Z => n32);
   U7 : CLKBUF_X1 port map( A => n37, Z => cout_0_port);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity BTB_PC_SIZE32_BTBSIZE5_DW01_cmp6_0 is

   port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, GT,
         EQ, LE, GE, NE : out std_logic);

end BTB_PC_SIZE32_BTBSIZE5_DW01_cmp6_0;

architecture SYN_rpl of BTB_PC_SIZE32_BTBSIZE5_DW01_cmp6_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47 : std_logic;

begin
   
   U1 : NOR4_X1 port map( A1 => n1, A2 => n2, A3 => n3, A4 => n4, ZN => EQ);
   U2 : NAND4_X1 port map( A1 => n5, A2 => n6, A3 => n7, A4 => n8, ZN => n4);
   U3 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n8);
   U4 : XNOR2_X1 port map( A => B(4), B => A(4), ZN => n7);
   U5 : XNOR2_X1 port map( A => B(5), B => A(5), ZN => n6);
   U6 : XNOR2_X1 port map( A => B(6), B => A(6), ZN => n5);
   U7 : NAND4_X1 port map( A1 => n9, A2 => n10, A3 => n11, A4 => n12, ZN => n3)
                           ;
   U8 : OAI22_X1 port map( A1 => n13, A2 => n14, B1 => B(1), B2 => n13, ZN => 
                           n12);
   U9 : INV_X1 port map( A => A(1), ZN => n14);
   U10 : AND2_X1 port map( A1 => B(0), A2 => n15, ZN => n13);
   U11 : OAI22_X1 port map( A1 => A(1), A2 => n16, B1 => n16, B2 => n17, ZN => 
                           n11);
   U12 : INV_X1 port map( A => B(1), ZN => n17);
   U13 : NOR2_X1 port map( A1 => n15, A2 => B(0), ZN => n16);
   U14 : INV_X1 port map( A => A(0), ZN => n15);
   U15 : XNOR2_X1 port map( A => B(31), B => A(31), ZN => n10);
   U16 : XNOR2_X1 port map( A => B(2), B => A(2), ZN => n9);
   U17 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => n2);
   U18 : NOR4_X1 port map( A1 => n20, A2 => n21, A3 => n22, A4 => n23, ZN => 
                           n19);
   U19 : XOR2_X1 port map( A => B(10), B => A(10), Z => n23);
   U20 : XOR2_X1 port map( A => B(9), B => A(9), Z => n22);
   U21 : XOR2_X1 port map( A => B(8), B => A(8), Z => n21);
   U22 : XOR2_X1 port map( A => B(7), B => A(7), Z => n20);
   U23 : NOR4_X1 port map( A1 => n24, A2 => n25, A3 => n26, A4 => n27, ZN => 
                           n18);
   U24 : XOR2_X1 port map( A => B(14), B => A(14), Z => n27);
   U25 : XOR2_X1 port map( A => B(13), B => A(13), Z => n26);
   U26 : XOR2_X1 port map( A => B(12), B => A(12), Z => n25);
   U27 : XOR2_X1 port map( A => B(11), B => A(11), Z => n24);
   U28 : NAND4_X1 port map( A1 => n28, A2 => n29, A3 => n30, A4 => n31, ZN => 
                           n1);
   U29 : NOR4_X1 port map( A1 => n32, A2 => n33, A3 => n34, A4 => n35, ZN => 
                           n31);
   U30 : XOR2_X1 port map( A => B(18), B => A(18), Z => n35);
   U31 : XOR2_X1 port map( A => B(17), B => A(17), Z => n34);
   U32 : XOR2_X1 port map( A => B(16), B => A(16), Z => n33);
   U33 : XOR2_X1 port map( A => B(15), B => A(15), Z => n32);
   U34 : NOR4_X1 port map( A1 => n36, A2 => n37, A3 => n38, A4 => n39, ZN => 
                           n30);
   U35 : XOR2_X1 port map( A => B(22), B => A(22), Z => n39);
   U36 : XOR2_X1 port map( A => B(21), B => A(21), Z => n38);
   U37 : XOR2_X1 port map( A => B(20), B => A(20), Z => n37);
   U38 : XOR2_X1 port map( A => B(19), B => A(19), Z => n36);
   U39 : NOR4_X1 port map( A1 => n40, A2 => n41, A3 => n42, A4 => n43, ZN => 
                           n29);
   U40 : XOR2_X1 port map( A => B(26), B => A(26), Z => n43);
   U41 : XOR2_X1 port map( A => B(25), B => A(25), Z => n42);
   U42 : XOR2_X1 port map( A => B(24), B => A(24), Z => n41);
   U43 : XOR2_X1 port map( A => B(23), B => A(23), Z => n40);
   U44 : NOR4_X1 port map( A1 => n44, A2 => n45, A3 => n46, A4 => n47, ZN => 
                           n28);
   U45 : XOR2_X1 port map( A => B(30), B => A(30), Z => n47);
   U46 : XOR2_X1 port map( A => B(29), B => A(29), Z => n46);
   U47 : XOR2_X1 port map( A => B(28), B => A(28), Z => n45);
   U48 : XOR2_X1 port map( A => B(27), B => A(27), Z => n44);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ForwardingUnit_NUMBIT32_ADDRESS_WIDTH_RF5 is

   port( CLK, RST : in std_logic;  RS1, RS2, RD_XM, RD_MW : in std_logic_vector
         (4 downto 0);  REGWRITE_XM, REGWRITE_MW : in std_logic;  ForwardA, 
         forwardB : out std_logic_vector (1 downto 0);  ForwardC : out 
         std_logic;  ForwardD : out std_logic_vector (1 downto 0));

end ForwardingUnit_NUMBIT32_ADDRESS_WIDTH_RF5;

architecture SYN_beh of ForwardingUnit_NUMBIT32_ADDRESS_WIDTH_RF5 is

   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR4_X4
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal N13, N14, N15, N16, N17, N18, N19, N20, n19_port, n20_port, n21, n61,
      n62, n63, n64, n65, net78471, net78472, net78473, net78475, net78476, 
      net78477, net78478, net78479, net78481, net78482, net78630, net78629, 
      net78628, net78621, net78620, net78618, net78611, net78608, net78606, 
      net78605, net78601, net78593, net78592, net78566, net78565, net78564, 
      net78563, net78562, net78559, net78558, net95388, net95387, net95500, 
      net95502, net95508, net95512, net95523, net95526, net95528, net95530, 
      net95540, net95557, net95493, net98500, net98509, net95345, net95344, 
      net78582, net78580, net78572, net78571, net78569, net78570, net78568, 
      net78576, net78575, net78574, net78573, net78567, net78579, net78577, n1,
      n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n14_port, n15_port, n16_port, 
      n17_port, n18_port, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32
      , n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, 
      n47, n48, n49, n50, n51, net114862, net114863, net114864, net114865, 
      net114866, net114867, net114868, net114869, n52, n53, n54 : std_logic;

begin
   
   RS1_DX_reg_4_inst : DFF_X1 port map( D => N17, CK => CLK, Q => net114869, QN
                           => n19_port);
   RS1_DX_reg_3_inst : DFF_X1 port map( D => N16, CK => CLK, Q => net114868, QN
                           => n20_port);
   RS1_DX_reg_2_inst : DFF_X1 port map( D => N15, CK => CLK, Q => net114867, QN
                           => n21);
   RS1_DX_reg_1_inst : DFF_X1 port map( D => N14, CK => CLK, Q => net114866, QN
                           => net78482);
   RS1_DX_reg_0_inst : DFF_X1 port map( D => N13, CK => CLK, Q => net114865, QN
                           => net78481);
   RS2_DX_reg_2_inst : DFF_X1 port map( D => N20, CK => CLK, Q => net114864, QN
                           => net78478);
   RS2_DX_reg_1_inst : DFF_X1 port map( D => N19, CK => CLK, Q => net114863, QN
                           => net78477);
   RS2_DX_reg_0_inst : DFF_X1 port map( D => N18, CK => CLK, Q => net114862, QN
                           => net78476);
   RS2_DX_reg_4_inst : DFF_X1 port map( D => n9, CK => CLK, Q => net78559, QN 
                           => net95493);
   RS2_XM_reg_4_inst : DFF_X1 port map( D => n65, CK => CLK, Q => net78558, QN 
                           => net78475);
   RS2_XM_reg_3_inst : DFF_X1 port map( D => n64, CK => CLK, Q => n14_port, QN 
                           => n51);
   RS2_XM_reg_2_inst : DFF_X1 port map( D => n63, CK => CLK, Q => n5, QN => 
                           net78473);
   RS2_XM_reg_1_inst : DFF_X1 port map( D => n62, CK => CLK, Q => n4, QN => 
                           net78472);
   RS2_XM_reg_0_inst : DFF_X1 port map( D => n61, CK => CLK, Q => n3, QN => 
                           net78471);
   U3 : OR4_X1 port map( A1 => n35, A2 => net78592, A3 => net78608, A4 => n36, 
                           ZN => n1);
   U4 : INV_X2 port map( A => n1, ZN => ForwardC);
   U5 : NAND4_X2 port map( A1 => n37, A2 => net78611, A3 => n38, A4 => n39, ZN 
                           => n35);
   U6 : NOR2_X1 port map( A1 => n6, A2 => net78579, ZN => net78577);
   U7 : NAND4_X1 port map( A1 => net78577, A2 => net78575, A3 => net78576, A4 
                           => net78574, ZN => net78567);
   U8 : XNOR2_X1 port map( A => RD_XM(4), B => net95493, ZN => net78579);
   U9 : XOR2_X1 port map( A => RD_XM(3), B => net95526, Z => n6);
   U10 : BUF_X1 port map( A => RD_XM(4), Z => net95557);
   U11 : XNOR2_X1 port map( A => RD_XM(4), B => n19_port, ZN => net78628);
   U12 : XOR2_X1 port map( A => net95493, B => RD_MW(4), Z => net78580);
   U13 : BUF_X1 port map( A => RD_XM(3), Z => net95502);
   U14 : NOR2_X1 port map( A1 => net78559, A2 => net95526, ZN => net78573);
   U15 : OAI21_X1 port map( B1 => net78567, B2 => net78565, A => net78568, ZN 
                           => net78570);
   U16 : NOR2_X1 port map( A1 => net95388, A2 => net78567, ZN => forwardB(1));
   U17 : XOR2_X1 port map( A => net78476, B => RD_XM(0), Z => net78574);
   U18 : XOR2_X1 port map( A => net78477, B => RD_XM(1), Z => net78576);
   U19 : XOR2_X1 port map( A => net78478, B => RD_XM(2), Z => net78575);
   U20 : MUX2_X1 port map( A => net78471, B => net78476, S => n53, Z => 
                           net78564);
   U21 : XNOR2_X1 port map( A => RD_MW(0), B => net78476, ZN => net78571);
   U22 : NAND4_X1 port map( A1 => net78476, A2 => net78478, A3 => net78477, A4 
                           => net78573, ZN => net78568);
   U23 : CLKBUF_X1 port map( A => RD_XM(0), Z => net95512);
   U24 : MUX2_X1 port map( A => net78472, B => net78477, S => n53, Z => 
                           net78563);
   U25 : XNOR2_X1 port map( A => RD_MW(1), B => net78477, ZN => net78572);
   U26 : BUF_X1 port map( A => RD_XM(1), Z => net95528);
   U27 : MUX2_X1 port map( A => net78473, B => net78478, S => n53, Z => 
                           net78562);
   U28 : XOR2_X1 port map( A => net78478, B => RD_MW(2), Z => net78582);
   U29 : BUF_X1 port map( A => RD_XM(2), Z => net95540);
   U30 : NOR3_X2 port map( A1 => net78570, A2 => net78569, A3 => net95345, ZN 
                           => forwardB(0));
   U31 : INV_X2 port map( A => REGWRITE_XM, ZN => net78565);
   U32 : INV_X1 port map( A => net78568, ZN => net78566);
   U33 : MUX2_X1 port map( A => net78558, B => net78559, S => n53, Z => n65);
   U34 : INV_X1 port map( A => net95344, ZN => net95345);
   U35 : NOR2_X1 port map( A1 => net78572, A2 => net78571, ZN => net95344);
   U36 : NAND4_X1 port map( A1 => REGWRITE_MW, A2 => net78580, A3 => n7, A4 => 
                           net78582, ZN => net78569);
   U37 : XOR2_X1 port map( A => net78479, B => RD_MW(3), Z => n7);
   U38 : CLKBUF_X1 port map( A => RD_MW(0), Z => net98500);
   U39 : XOR2_X1 port map( A => RS1(0), B => RD_MW(0), Z => net78593);
   U40 : BUF_X2 port map( A => RD_MW(1), Z => net98509);
   U41 : NAND4_X1 port map( A1 => REGWRITE_MW, A2 => net78629, A3 => net78630, 
                           A4 => n8, ZN => net78618);
   U42 : INV_X1 port map( A => REGWRITE_MW, ZN => net78592);
   U43 : XOR2_X1 port map( A => n21, B => RD_MW(2), Z => n8);
   U44 : INV_X1 port map( A => RD_MW(2), ZN => net78606);
   U46 : BUF_X1 port map( A => RD_MW(3), Z => net95530);
   U47 : BUF_X2 port map( A => RD_MW(4), Z => net95508);
   U48 : AND2_X1 port map( A1 => RS2(4), A2 => n53, ZN => n9);
   U49 : XOR2_X1 port map( A => net78471, B => net98500, Z => net78611);
   U50 : XNOR2_X1 port map( A => net78481, B => net98500, ZN => net78620);
   U51 : XNOR2_X1 port map( A => net98509, B => RS1(1), ZN => net78605);
   U52 : XNOR2_X1 port map( A => net78472, B => net98509, ZN => net78608);
   U53 : XNOR2_X1 port map( A => net78482, B => net98509, ZN => net78621);
   U54 : CLKBUF_X1 port map( A => net95526, Z => net95523);
   U55 : CLKBUF_X1 port map( A => net95530, Z => net95500);
   U56 : NAND2_X1 port map( A1 => n11, A2 => n12, ZN => n10);
   U57 : AND4_X1 port map( A1 => n32, A2 => n33, A3 => n34, A4 => net78605, ZN 
                           => n11);
   U58 : NOR2_X1 port map( A1 => net78566, A2 => net78565, ZN => net95387);
   U59 : INV_X1 port map( A => net95387, ZN => net95388);
   U60 : NOR3_X1 port map( A1 => n18_port, A2 => n22, A3 => net78565, ZN => 
                           ForwardD(1));
   U61 : NOR2_X2 port map( A1 => n24, A2 => n10, ZN => ForwardD(0));
   U62 : NOR4_X4 port map( A1 => net78618, A2 => n44, A3 => net78620, A4 => 
                           net78621, ZN => ForwardA(0));
   U63 : NOR2_X1 port map( A1 => net78593, A2 => net78592, ZN => n12);
   U67 : MUX2_X1 port map( A => n14_port, B => net95523, S => n53, Z => n64);
   U68 : INV_X1 port map( A => net78562, ZN => n63);
   U69 : INV_X1 port map( A => net78563, ZN => n62);
   U70 : INV_X1 port map( A => net78564, ZN => n61);
   U71 : AND2_X1 port map( A1 => RS2(2), A2 => n53, ZN => N20);
   U72 : AND2_X1 port map( A1 => RS2(1), A2 => n53, ZN => N19);
   U73 : AND2_X1 port map( A1 => RS2(0), A2 => n53, ZN => N18);
   U74 : NOR2_X1 port map( A1 => n54, A2 => n15_port, ZN => N17);
   U75 : NOR2_X1 port map( A1 => n54, A2 => n16_port, ZN => N16);
   U76 : NOR2_X1 port map( A1 => n54, A2 => n17_port, ZN => N15);
   U77 : AND2_X1 port map( A1 => n53, A2 => RS1(1), ZN => N14);
   U78 : AND2_X1 port map( A1 => n53, A2 => RS1(0), ZN => N13);
   U79 : INV_X1 port map( A => n23, ZN => n22);
   U80 : OAI21_X1 port map( B1 => net78565, B2 => n18_port, A => n23, ZN => n24
                           );
   U81 : NAND4_X1 port map( A1 => n16_port, A2 => n15_port, A3 => n17_port, A4 
                           => n25, ZN => n23);
   U82 : NOR2_X1 port map( A1 => RS1(1), A2 => RS1(0), ZN => n25);
   U83 : INV_X1 port map( A => RS1(2), ZN => n17_port);
   U84 : NAND4_X1 port map( A1 => n29, A2 => n27, A3 => n28, A4 => n26, ZN => 
                           n18_port);
   U85 : NOR2_X1 port map( A1 => n30, A2 => n31, ZN => n29);
   U86 : XOR2_X1 port map( A => RS1(4), B => net95557, Z => n31);
   U87 : XOR2_X1 port map( A => RS1(3), B => net95502, Z => n30);
   U88 : XNOR2_X1 port map( A => net95528, B => RS1(1), ZN => n28);
   U89 : XOR2_X1 port map( A => net78601, B => RS1(2), Z => n27);
   U90 : INV_X1 port map( A => net95540, ZN => net78601);
   U91 : XNOR2_X1 port map( A => net95512, B => RS1(0), ZN => n26);
   U92 : XOR2_X1 port map( A => net78606, B => RS1(2), Z => n34);
   U93 : XOR2_X1 port map( A => net95530, B => n16_port, Z => n33);
   U94 : INV_X1 port map( A => RS1(3), ZN => n16_port);
   U95 : XOR2_X1 port map( A => net95508, B => n15_port, Z => n32);
   U96 : INV_X1 port map( A => RS1(4), ZN => n15_port);
   U97 : XOR2_X1 port map( A => net78473, B => net78606, Z => n36);
   U98 : NAND4_X1 port map( A1 => net78472, A2 => net78471, A3 => net78473, A4 
                           => n40, ZN => n39);
   U99 : NOR2_X1 port map( A1 => n14_port, A2 => net78558, ZN => n40);
   U100 : XOR2_X1 port map( A => n51, B => net95500, Z => n38);
   U101 : XOR2_X1 port map( A => net78475, B => net95508, Z => n37);
   U102 : NOR3_X1 port map( A1 => n41, A2 => n42, A3 => net78565, ZN => 
                           ForwardA(1));
   U103 : INV_X1 port map( A => n43, ZN => n42);
   U104 : OAI21_X1 port map( B1 => net78565, B2 => n41, A => n43, ZN => n44);
   U105 : NAND4_X1 port map( A1 => net78481, A2 => n21, A3 => net78482, A4 => 
                           n45, ZN => n43);
   U106 : AND2_X1 port map( A1 => n20_port, A2 => n19_port, ZN => n45);
   U107 : NAND4_X1 port map( A1 => n46, A2 => n47, A3 => n48, A4 => n49, ZN => 
                           n41);
   U108 : NOR2_X1 port map( A1 => n50, A2 => net78628, ZN => n49);
   U109 : XNOR2_X1 port map( A => net95502, B => n20_port, ZN => n50);
   U110 : XOR2_X1 port map( A => net78482, B => net95528, Z => n48);
   U111 : XOR2_X1 port map( A => n21, B => net95540, Z => n47);
   U112 : XOR2_X1 port map( A => net78481, B => net95512, Z => n46);
   U113 : XOR2_X1 port map( A => n20_port, B => net95530, Z => net78630);
   U114 : XOR2_X1 port map( A => n19_port, B => net95508, Z => net78629);
   RS2_DX_reg_3_inst : DFF_X1 port map( D => n52, CK => CLK, Q => net95526, QN 
                           => net78479);
   U45 : AND2_X1 port map( A1 => RS2(3), A2 => n53, ZN => n52);
   U64 : INV_X1 port map( A => n54, ZN => n53);
   U65 : INV_X2 port map( A => RST, ZN => n54);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_N5 is

   port( A, B : in std_logic_vector (4 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (4 downto 0));

end MUX21_GENERIC_N5;

architecture SYN_BEHAVIORAL_1 of MUX21_GENERIC_N5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Y(4));
   U2 : AOI22_X1 port map( A1 => SEL, A2 => A(4), B1 => B(4), B2 => n3, ZN => 
                           n2);
   U3 : INV_X1 port map( A => n4, ZN => Y(3));
   U4 : AOI22_X1 port map( A1 => A(3), A2 => SEL, B1 => B(3), B2 => n3, ZN => 
                           n4);
   U5 : INV_X1 port map( A => n5, ZN => Y(2));
   U6 : AOI22_X1 port map( A1 => A(2), A2 => SEL, B1 => B(2), B2 => n3, ZN => 
                           n5);
   U7 : INV_X1 port map( A => n6, ZN => Y(1));
   U8 : AOI22_X1 port map( A1 => A(1), A2 => SEL, B1 => B(1), B2 => n3, ZN => 
                           n6);
   U9 : INV_X1 port map( A => n7, ZN => Y(0));
   U10 : AOI22_X1 port map( A1 => A(0), A2 => SEL, B1 => B(0), B2 => n3, ZN => 
                           n7);
   U11 : INV_X1 port map( A => SEL, ZN => n3);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21 is

   port( A, B, SEL : in std_logic;  Y : out std_logic);

end MUX21;

architecture SYN_BEHAVIORAL_1 of MUX21 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n2, n3 : std_logic;

begin
   
   U3 : INV_X1 port map( A => SEL, ZN => n3);
   U1 : BUF_X2 port map( A => n4, Z => Y);
   U2 : INV_X1 port map( A => n2, ZN => n4);
   U4 : AOI22_X1 port map( A1 => SEL, A2 => A, B1 => B, B2 => n3, ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity BranchMgmt_NUMBIT32 is

   port( Rin : in std_logic_vector (31 downto 0);  Cond, Jump : in std_logic;  
         Branch : out std_logic);

end BranchMgmt_NUMBIT32;

architecture SYN_Behavioral of BranchMgmt_NUMBIT32 is

   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U2 : OR2_X1 port map( A1 => n2, A2 => Jump, ZN => Branch);
   U3 : XNOR2_X1 port map( A => n3, B => Cond, ZN => n2);
   U4 : NOR2_X1 port map( A1 => n4, A2 => n5, ZN => n3);
   U5 : NAND4_X1 port map( A1 => n6, A2 => n7, A3 => n8, A4 => n9, ZN => n5);
   U6 : NOR4_X1 port map( A1 => Rin(23), A2 => Rin(22), A3 => Rin(21), A4 => 
                           Rin(20), ZN => n9);
   U7 : NOR4_X1 port map( A1 => Rin(1), A2 => Rin(19), A3 => Rin(18), A4 => 
                           Rin(17), ZN => n8);
   U8 : NOR4_X1 port map( A1 => Rin(16), A2 => Rin(15), A3 => Rin(14), A4 => 
                           Rin(13), ZN => n7);
   U9 : NOR4_X1 port map( A1 => Rin(12), A2 => Rin(11), A3 => Rin(10), A4 => 
                           Rin(0), ZN => n6);
   U10 : NAND4_X1 port map( A1 => n12, A2 => n11, A3 => n10, A4 => n13, ZN => 
                           n4);
   U11 : NOR4_X1 port map( A1 => Rin(9), A2 => Rin(8), A3 => Rin(7), A4 => 
                           Rin(6), ZN => n13);
   U12 : NOR4_X1 port map( A1 => Rin(5), A2 => Rin(4), A3 => Rin(3), A4 => 
                           Rin(31), ZN => n12);
   U13 : NOR4_X1 port map( A1 => Rin(30), A2 => Rin(2), A3 => Rin(29), A4 => 
                           Rin(28), ZN => n11);
   U14 : NOR4_X1 port map( A1 => Rin(27), A2 => Rin(26), A3 => Rin(25), A4 => 
                           Rin(24), ZN => n10);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity signExtend_NUMBIT_in26_NUMBIT_out32 is

   port( in_s : in std_logic_vector (25 downto 0);  sign_unsign : in std_logic;
         out_s : out std_logic_vector (31 downto 0));

end signExtend_NUMBIT_in26_NUMBIT_out32;

architecture SYN_beh of signExtend_NUMBIT_in26_NUMBIT_out32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal out_s_31 : std_logic;

begin
   out_s <= ( out_s_31, out_s_31, out_s_31, out_s_31, out_s_31, out_s_31, 
      in_s(25), in_s(24), in_s(23), in_s(22), in_s(21), in_s(20), in_s(19), 
      in_s(18), in_s(17), in_s(16), in_s(15), in_s(14), in_s(13), in_s(12), 
      in_s(11), in_s(10), in_s(9), in_s(8), in_s(7), in_s(6), in_s(5), in_s(4),
      in_s(3), in_s(2), in_s(1), in_s(0) );
   
   U1 : AND2_X1 port map( A1 => sign_unsign, A2 => in_s(25), ZN => out_s_31);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity signExtend_NUMBIT_in16_NUMBIT_out32 is

   port( in_s : in std_logic_vector (15 downto 0);  sign_unsign : in std_logic;
         out_s : out std_logic_vector (31 downto 0));

end signExtend_NUMBIT_in16_NUMBIT_out32;

architecture SYN_beh of signExtend_NUMBIT_in16_NUMBIT_out32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal out_s_31 : std_logic;

begin
   out_s <= ( out_s_31, out_s_31, out_s_31, out_s_31, out_s_31, out_s_31, 
      out_s_31, out_s_31, out_s_31, out_s_31, out_s_31, out_s_31, out_s_31, 
      out_s_31, out_s_31, out_s_31, in_s(15), in_s(14), in_s(13), in_s(12), 
      in_s(11), in_s(10), in_s(9), in_s(8), in_s(7), in_s(6), in_s(5), in_s(4),
      in_s(3), in_s(2), in_s(1), in_s(0) );
   
   U1 : AND2_X1 port map( A1 => sign_unsign, A2 => in_s(15), ZN => out_s_31);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity register_file_NUMBIT32_BITADDR5 is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0));

end register_file_NUMBIT32_BITADDR5;

architecture SYN_A of register_file_NUMBIT32_BITADDR5 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal REGISTERS_1_31_port, REGISTERS_1_30_port, REGISTERS_1_29_port, 
      REGISTERS_1_28_port, REGISTERS_1_27_port, REGISTERS_1_26_port, 
      REGISTERS_1_25_port, REGISTERS_1_24_port, REGISTERS_1_23_port, 
      REGISTERS_1_22_port, REGISTERS_1_21_port, REGISTERS_1_20_port, 
      REGISTERS_1_19_port, REGISTERS_1_18_port, REGISTERS_1_17_port, 
      REGISTERS_1_16_port, REGISTERS_1_15_port, REGISTERS_1_14_port, 
      REGISTERS_1_13_port, REGISTERS_1_12_port, REGISTERS_1_11_port, 
      REGISTERS_1_10_port, REGISTERS_1_9_port, REGISTERS_1_8_port, 
      REGISTERS_1_7_port, REGISTERS_1_6_port, REGISTERS_1_5_port, 
      REGISTERS_1_4_port, REGISTERS_1_3_port, REGISTERS_1_2_port, 
      REGISTERS_1_1_port, REGISTERS_1_0_port, REGISTERS_2_31_port, 
      REGISTERS_2_30_port, REGISTERS_2_29_port, REGISTERS_2_28_port, 
      REGISTERS_2_27_port, REGISTERS_2_26_port, REGISTERS_2_25_port, 
      REGISTERS_2_24_port, REGISTERS_2_23_port, REGISTERS_2_22_port, 
      REGISTERS_2_21_port, REGISTERS_2_20_port, REGISTERS_2_19_port, 
      REGISTERS_2_18_port, REGISTERS_2_17_port, REGISTERS_2_16_port, 
      REGISTERS_2_15_port, REGISTERS_2_14_port, REGISTERS_2_13_port, 
      REGISTERS_2_12_port, REGISTERS_2_11_port, REGISTERS_2_10_port, 
      REGISTERS_2_9_port, REGISTERS_2_8_port, REGISTERS_2_7_port, 
      REGISTERS_2_6_port, REGISTERS_2_5_port, REGISTERS_2_4_port, 
      REGISTERS_2_3_port, REGISTERS_2_2_port, REGISTERS_2_1_port, 
      REGISTERS_2_0_port, REGISTERS_3_31_port, REGISTERS_3_30_port, 
      REGISTERS_3_29_port, REGISTERS_3_28_port, REGISTERS_3_27_port, 
      REGISTERS_3_26_port, REGISTERS_3_25_port, REGISTERS_3_24_port, 
      REGISTERS_3_23_port, REGISTERS_3_22_port, REGISTERS_3_21_port, 
      REGISTERS_3_20_port, REGISTERS_3_19_port, REGISTERS_3_18_port, 
      REGISTERS_3_17_port, REGISTERS_3_16_port, REGISTERS_3_15_port, 
      REGISTERS_3_14_port, REGISTERS_3_13_port, REGISTERS_3_12_port, 
      REGISTERS_3_11_port, REGISTERS_3_10_port, REGISTERS_3_9_port, 
      REGISTERS_3_8_port, REGISTERS_3_7_port, REGISTERS_3_6_port, 
      REGISTERS_3_5_port, REGISTERS_3_4_port, REGISTERS_3_3_port, 
      REGISTERS_3_2_port, REGISTERS_3_1_port, REGISTERS_3_0_port, 
      REGISTERS_4_31_port, REGISTERS_4_30_port, REGISTERS_4_29_port, 
      REGISTERS_4_28_port, REGISTERS_4_27_port, REGISTERS_4_26_port, 
      REGISTERS_4_25_port, REGISTERS_4_24_port, REGISTERS_4_23_port, 
      REGISTERS_4_22_port, REGISTERS_4_21_port, REGISTERS_4_20_port, 
      REGISTERS_4_19_port, REGISTERS_4_18_port, REGISTERS_4_17_port, 
      REGISTERS_4_16_port, REGISTERS_4_15_port, REGISTERS_4_14_port, 
      REGISTERS_4_13_port, REGISTERS_4_12_port, REGISTERS_4_11_port, 
      REGISTERS_4_10_port, REGISTERS_4_9_port, REGISTERS_4_8_port, 
      REGISTERS_4_7_port, REGISTERS_4_6_port, REGISTERS_4_5_port, 
      REGISTERS_4_4_port, REGISTERS_4_3_port, REGISTERS_4_2_port, 
      REGISTERS_4_1_port, REGISTERS_4_0_port, REGISTERS_5_31_port, 
      REGISTERS_5_30_port, REGISTERS_5_29_port, REGISTERS_5_28_port, 
      REGISTERS_5_27_port, REGISTERS_5_26_port, REGISTERS_5_25_port, 
      REGISTERS_5_24_port, REGISTERS_5_23_port, REGISTERS_5_22_port, 
      REGISTERS_5_21_port, REGISTERS_5_20_port, REGISTERS_5_19_port, 
      REGISTERS_5_18_port, REGISTERS_5_17_port, REGISTERS_5_16_port, 
      REGISTERS_5_15_port, REGISTERS_5_14_port, REGISTERS_5_13_port, 
      REGISTERS_5_12_port, REGISTERS_5_11_port, REGISTERS_5_10_port, 
      REGISTERS_5_9_port, REGISTERS_5_8_port, REGISTERS_5_7_port, 
      REGISTERS_5_6_port, REGISTERS_5_5_port, REGISTERS_5_4_port, 
      REGISTERS_5_3_port, REGISTERS_5_2_port, REGISTERS_5_1_port, 
      REGISTERS_5_0_port, REGISTERS_6_31_port, REGISTERS_6_30_port, 
      REGISTERS_6_29_port, REGISTERS_6_28_port, REGISTERS_6_27_port, 
      REGISTERS_6_26_port, REGISTERS_6_25_port, REGISTERS_6_24_port, 
      REGISTERS_6_23_port, REGISTERS_6_22_port, REGISTERS_6_21_port, 
      REGISTERS_6_20_port, REGISTERS_6_19_port, REGISTERS_6_18_port, 
      REGISTERS_6_17_port, REGISTERS_6_16_port, REGISTERS_6_15_port, 
      REGISTERS_6_14_port, REGISTERS_6_13_port, REGISTERS_6_12_port, 
      REGISTERS_6_11_port, REGISTERS_6_10_port, REGISTERS_6_9_port, 
      REGISTERS_6_8_port, REGISTERS_6_7_port, REGISTERS_6_6_port, 
      REGISTERS_6_5_port, REGISTERS_6_4_port, REGISTERS_6_3_port, 
      REGISTERS_6_2_port, REGISTERS_6_1_port, REGISTERS_6_0_port, 
      REGISTERS_7_31_port, REGISTERS_7_30_port, REGISTERS_7_29_port, 
      REGISTERS_7_28_port, REGISTERS_7_27_port, REGISTERS_7_26_port, 
      REGISTERS_7_25_port, REGISTERS_7_24_port, REGISTERS_7_23_port, 
      REGISTERS_7_22_port, REGISTERS_7_21_port, REGISTERS_7_20_port, 
      REGISTERS_7_19_port, REGISTERS_7_18_port, REGISTERS_7_17_port, 
      REGISTERS_7_16_port, REGISTERS_7_15_port, REGISTERS_7_14_port, 
      REGISTERS_7_13_port, REGISTERS_7_12_port, REGISTERS_7_11_port, 
      REGISTERS_7_10_port, REGISTERS_7_9_port, REGISTERS_7_8_port, 
      REGISTERS_7_7_port, REGISTERS_7_6_port, REGISTERS_7_5_port, 
      REGISTERS_7_4_port, REGISTERS_7_3_port, REGISTERS_7_2_port, 
      REGISTERS_7_1_port, REGISTERS_7_0_port, REGISTERS_8_31_port, 
      REGISTERS_8_30_port, REGISTERS_8_29_port, REGISTERS_8_28_port, 
      REGISTERS_8_27_port, REGISTERS_8_26_port, REGISTERS_8_25_port, 
      REGISTERS_8_24_port, REGISTERS_8_23_port, REGISTERS_8_22_port, 
      REGISTERS_8_21_port, REGISTERS_8_20_port, REGISTERS_8_19_port, 
      REGISTERS_8_18_port, REGISTERS_8_17_port, REGISTERS_8_16_port, 
      REGISTERS_8_15_port, REGISTERS_8_14_port, REGISTERS_8_13_port, 
      REGISTERS_8_12_port, REGISTERS_8_11_port, REGISTERS_8_10_port, 
      REGISTERS_8_9_port, REGISTERS_8_8_port, REGISTERS_8_7_port, 
      REGISTERS_8_6_port, REGISTERS_8_5_port, REGISTERS_8_4_port, 
      REGISTERS_8_3_port, REGISTERS_8_2_port, REGISTERS_8_1_port, 
      REGISTERS_8_0_port, REGISTERS_9_31_port, REGISTERS_9_30_port, 
      REGISTERS_9_29_port, REGISTERS_9_28_port, REGISTERS_9_27_port, 
      REGISTERS_9_26_port, REGISTERS_9_25_port, REGISTERS_9_24_port, 
      REGISTERS_9_23_port, REGISTERS_9_22_port, REGISTERS_9_21_port, 
      REGISTERS_9_20_port, REGISTERS_9_19_port, REGISTERS_9_18_port, 
      REGISTERS_9_17_port, REGISTERS_9_16_port, REGISTERS_9_15_port, 
      REGISTERS_9_14_port, REGISTERS_9_13_port, REGISTERS_9_12_port, 
      REGISTERS_9_11_port, REGISTERS_9_10_port, REGISTERS_9_9_port, 
      REGISTERS_9_8_port, REGISTERS_9_7_port, REGISTERS_9_6_port, 
      REGISTERS_9_5_port, REGISTERS_9_4_port, REGISTERS_9_3_port, 
      REGISTERS_9_2_port, REGISTERS_9_1_port, REGISTERS_9_0_port, 
      REGISTERS_10_31_port, REGISTERS_10_30_port, REGISTERS_10_29_port, 
      REGISTERS_10_28_port, REGISTERS_10_27_port, REGISTERS_10_26_port, 
      REGISTERS_10_25_port, REGISTERS_10_24_port, REGISTERS_10_23_port, 
      REGISTERS_10_22_port, REGISTERS_10_21_port, REGISTERS_10_20_port, 
      REGISTERS_10_19_port, REGISTERS_10_18_port, REGISTERS_10_17_port, 
      REGISTERS_10_16_port, REGISTERS_10_15_port, REGISTERS_10_14_port, 
      REGISTERS_10_13_port, REGISTERS_10_12_port, REGISTERS_10_11_port, 
      REGISTERS_10_10_port, REGISTERS_10_9_port, REGISTERS_10_8_port, 
      REGISTERS_10_7_port, REGISTERS_10_6_port, REGISTERS_10_5_port, 
      REGISTERS_10_4_port, REGISTERS_10_3_port, REGISTERS_10_2_port, 
      REGISTERS_10_1_port, REGISTERS_10_0_port, REGISTERS_11_31_port, 
      REGISTERS_11_30_port, REGISTERS_11_29_port, REGISTERS_11_28_port, 
      REGISTERS_11_27_port, REGISTERS_11_26_port, REGISTERS_11_25_port, 
      REGISTERS_11_24_port, REGISTERS_11_23_port, REGISTERS_11_22_port, 
      REGISTERS_11_21_port, REGISTERS_11_20_port, REGISTERS_11_19_port, 
      REGISTERS_11_18_port, REGISTERS_11_17_port, REGISTERS_11_16_port, 
      REGISTERS_11_15_port, REGISTERS_11_14_port, REGISTERS_11_13_port, 
      REGISTERS_11_12_port, REGISTERS_11_11_port, REGISTERS_11_10_port, 
      REGISTERS_11_9_port, REGISTERS_11_8_port, REGISTERS_11_7_port, 
      REGISTERS_11_6_port, REGISTERS_11_5_port, REGISTERS_11_4_port, 
      REGISTERS_11_3_port, REGISTERS_11_2_port, REGISTERS_11_1_port, 
      REGISTERS_11_0_port, REGISTERS_12_31_port, REGISTERS_12_30_port, 
      REGISTERS_12_29_port, REGISTERS_12_28_port, REGISTERS_12_27_port, 
      REGISTERS_12_26_port, REGISTERS_12_25_port, REGISTERS_12_24_port, 
      REGISTERS_12_23_port, REGISTERS_12_22_port, REGISTERS_12_21_port, 
      REGISTERS_12_20_port, REGISTERS_12_19_port, REGISTERS_12_18_port, 
      REGISTERS_12_17_port, REGISTERS_12_16_port, REGISTERS_12_15_port, 
      REGISTERS_12_14_port, REGISTERS_12_13_port, REGISTERS_12_12_port, 
      REGISTERS_12_11_port, REGISTERS_12_10_port, REGISTERS_12_9_port, 
      REGISTERS_12_8_port, REGISTERS_12_7_port, REGISTERS_12_6_port, 
      REGISTERS_12_5_port, REGISTERS_12_4_port, REGISTERS_12_3_port, 
      REGISTERS_12_2_port, REGISTERS_12_1_port, REGISTERS_12_0_port, 
      REGISTERS_13_31_port, REGISTERS_13_30_port, REGISTERS_13_29_port, 
      REGISTERS_13_28_port, REGISTERS_13_27_port, REGISTERS_13_26_port, 
      REGISTERS_13_25_port, REGISTERS_13_24_port, REGISTERS_13_23_port, 
      REGISTERS_13_22_port, REGISTERS_13_21_port, REGISTERS_13_20_port, 
      REGISTERS_13_19_port, REGISTERS_13_18_port, REGISTERS_13_17_port, 
      REGISTERS_13_16_port, REGISTERS_13_15_port, REGISTERS_13_14_port, 
      REGISTERS_13_13_port, REGISTERS_13_12_port, REGISTERS_13_11_port, 
      REGISTERS_13_10_port, REGISTERS_13_9_port, REGISTERS_13_8_port, 
      REGISTERS_13_7_port, REGISTERS_13_6_port, REGISTERS_13_5_port, 
      REGISTERS_13_4_port, REGISTERS_13_3_port, REGISTERS_13_2_port, 
      REGISTERS_13_1_port, REGISTERS_13_0_port, REGISTERS_14_31_port, 
      REGISTERS_14_30_port, REGISTERS_14_29_port, REGISTERS_14_28_port, 
      REGISTERS_14_27_port, REGISTERS_14_26_port, REGISTERS_14_25_port, 
      REGISTERS_14_24_port, REGISTERS_14_23_port, REGISTERS_14_22_port, 
      REGISTERS_14_21_port, REGISTERS_14_20_port, REGISTERS_14_19_port, 
      REGISTERS_14_18_port, REGISTERS_14_17_port, REGISTERS_14_16_port, 
      REGISTERS_14_15_port, REGISTERS_14_14_port, REGISTERS_14_13_port, 
      REGISTERS_14_12_port, REGISTERS_14_11_port, REGISTERS_14_10_port, 
      REGISTERS_14_9_port, REGISTERS_14_8_port, REGISTERS_14_7_port, 
      REGISTERS_14_6_port, REGISTERS_14_5_port, REGISTERS_14_4_port, 
      REGISTERS_14_3_port, REGISTERS_14_2_port, REGISTERS_14_1_port, 
      REGISTERS_14_0_port, REGISTERS_15_31_port, REGISTERS_15_30_port, 
      REGISTERS_15_29_port, REGISTERS_15_28_port, REGISTERS_15_27_port, 
      REGISTERS_15_26_port, REGISTERS_15_25_port, REGISTERS_15_24_port, 
      REGISTERS_15_23_port, REGISTERS_15_22_port, REGISTERS_15_21_port, 
      REGISTERS_15_20_port, REGISTERS_15_19_port, REGISTERS_15_18_port, 
      REGISTERS_15_17_port, REGISTERS_15_16_port, REGISTERS_15_15_port, 
      REGISTERS_15_14_port, REGISTERS_15_13_port, REGISTERS_15_12_port, 
      REGISTERS_15_11_port, REGISTERS_15_10_port, REGISTERS_15_9_port, 
      REGISTERS_15_8_port, REGISTERS_15_7_port, REGISTERS_15_6_port, 
      REGISTERS_15_5_port, REGISTERS_15_4_port, REGISTERS_15_3_port, 
      REGISTERS_15_2_port, REGISTERS_15_1_port, REGISTERS_15_0_port, 
      REGISTERS_16_31_port, REGISTERS_16_30_port, REGISTERS_16_29_port, 
      REGISTERS_16_28_port, REGISTERS_16_27_port, REGISTERS_16_26_port, 
      REGISTERS_16_25_port, REGISTERS_16_24_port, REGISTERS_16_23_port, 
      REGISTERS_16_22_port, REGISTERS_16_21_port, REGISTERS_16_20_port, 
      REGISTERS_16_19_port, REGISTERS_16_18_port, REGISTERS_16_17_port, 
      REGISTERS_16_16_port, REGISTERS_16_15_port, REGISTERS_16_14_port, 
      REGISTERS_16_13_port, REGISTERS_16_12_port, REGISTERS_16_11_port, 
      REGISTERS_16_10_port, REGISTERS_16_9_port, REGISTERS_16_8_port, 
      REGISTERS_16_7_port, REGISTERS_16_6_port, REGISTERS_16_5_port, 
      REGISTERS_16_4_port, REGISTERS_16_3_port, REGISTERS_16_2_port, 
      REGISTERS_16_1_port, REGISTERS_16_0_port, REGISTERS_17_31_port, 
      REGISTERS_17_30_port, REGISTERS_17_29_port, REGISTERS_17_28_port, 
      REGISTERS_17_27_port, REGISTERS_17_26_port, REGISTERS_17_25_port, 
      REGISTERS_17_24_port, REGISTERS_17_23_port, REGISTERS_17_22_port, 
      REGISTERS_17_21_port, REGISTERS_17_20_port, REGISTERS_17_19_port, 
      REGISTERS_17_18_port, REGISTERS_17_17_port, REGISTERS_17_16_port, 
      REGISTERS_17_15_port, REGISTERS_17_14_port, REGISTERS_17_13_port, 
      REGISTERS_17_12_port, REGISTERS_17_11_port, REGISTERS_17_10_port, 
      REGISTERS_17_9_port, REGISTERS_17_8_port, REGISTERS_17_7_port, 
      REGISTERS_17_6_port, REGISTERS_17_5_port, REGISTERS_17_4_port, 
      REGISTERS_17_3_port, REGISTERS_17_2_port, REGISTERS_17_1_port, 
      REGISTERS_17_0_port, REGISTERS_18_31_port, REGISTERS_18_30_port, 
      REGISTERS_18_29_port, REGISTERS_18_28_port, REGISTERS_18_27_port, 
      REGISTERS_18_26_port, REGISTERS_18_25_port, REGISTERS_18_24_port, 
      REGISTERS_18_23_port, REGISTERS_18_22_port, REGISTERS_18_21_port, 
      REGISTERS_18_20_port, REGISTERS_18_19_port, REGISTERS_18_18_port, 
      REGISTERS_18_17_port, REGISTERS_18_16_port, REGISTERS_18_15_port, 
      REGISTERS_18_14_port, REGISTERS_18_13_port, REGISTERS_18_12_port, 
      REGISTERS_18_11_port, REGISTERS_18_10_port, REGISTERS_18_9_port, 
      REGISTERS_18_8_port, REGISTERS_18_7_port, REGISTERS_18_6_port, 
      REGISTERS_18_5_port, REGISTERS_18_4_port, REGISTERS_18_3_port, 
      REGISTERS_18_2_port, REGISTERS_18_1_port, REGISTERS_18_0_port, 
      REGISTERS_19_31_port, REGISTERS_19_30_port, REGISTERS_19_29_port, 
      REGISTERS_19_28_port, REGISTERS_19_27_port, REGISTERS_19_26_port, 
      REGISTERS_19_25_port, REGISTERS_19_24_port, REGISTERS_19_23_port, 
      REGISTERS_19_22_port, REGISTERS_19_21_port, REGISTERS_19_20_port, 
      REGISTERS_19_19_port, REGISTERS_19_18_port, REGISTERS_19_17_port, 
      REGISTERS_19_16_port, REGISTERS_19_15_port, REGISTERS_19_14_port, 
      REGISTERS_19_13_port, REGISTERS_19_12_port, REGISTERS_19_11_port, 
      REGISTERS_19_10_port, REGISTERS_19_9_port, REGISTERS_19_8_port, 
      REGISTERS_19_7_port, REGISTERS_19_6_port, REGISTERS_19_5_port, 
      REGISTERS_19_4_port, REGISTERS_19_3_port, REGISTERS_19_2_port, 
      REGISTERS_19_1_port, REGISTERS_19_0_port, REGISTERS_20_31_port, 
      REGISTERS_20_30_port, REGISTERS_20_29_port, REGISTERS_20_28_port, 
      REGISTERS_20_27_port, REGISTERS_20_26_port, REGISTERS_20_25_port, 
      REGISTERS_20_24_port, REGISTERS_20_23_port, REGISTERS_20_22_port, 
      REGISTERS_20_21_port, REGISTERS_20_20_port, REGISTERS_20_19_port, 
      REGISTERS_20_18_port, REGISTERS_20_17_port, REGISTERS_20_16_port, 
      REGISTERS_20_15_port, REGISTERS_20_14_port, REGISTERS_20_13_port, 
      REGISTERS_20_12_port, REGISTERS_20_11_port, REGISTERS_20_10_port, 
      REGISTERS_20_9_port, REGISTERS_20_8_port, REGISTERS_20_7_port, 
      REGISTERS_20_6_port, REGISTERS_20_5_port, REGISTERS_20_4_port, 
      REGISTERS_20_3_port, REGISTERS_20_2_port, REGISTERS_20_1_port, 
      REGISTERS_20_0_port, REGISTERS_21_31_port, REGISTERS_21_30_port, 
      REGISTERS_21_29_port, REGISTERS_21_28_port, REGISTERS_21_27_port, 
      REGISTERS_21_26_port, REGISTERS_21_25_port, REGISTERS_21_24_port, 
      REGISTERS_21_23_port, REGISTERS_21_22_port, REGISTERS_21_21_port, 
      REGISTERS_21_20_port, REGISTERS_21_19_port, REGISTERS_21_18_port, 
      REGISTERS_21_17_port, REGISTERS_21_16_port, REGISTERS_21_15_port, 
      REGISTERS_21_14_port, REGISTERS_21_13_port, REGISTERS_21_12_port, 
      REGISTERS_21_11_port, REGISTERS_21_10_port, REGISTERS_21_9_port, 
      REGISTERS_21_8_port, REGISTERS_21_7_port, REGISTERS_21_6_port, 
      REGISTERS_21_5_port, REGISTERS_21_4_port, REGISTERS_21_3_port, 
      REGISTERS_21_2_port, REGISTERS_21_1_port, REGISTERS_21_0_port, 
      REGISTERS_22_31_port, REGISTERS_22_30_port, REGISTERS_22_29_port, 
      REGISTERS_22_28_port, REGISTERS_22_27_port, REGISTERS_22_26_port, 
      REGISTERS_22_25_port, REGISTERS_22_24_port, REGISTERS_22_23_port, 
      REGISTERS_22_22_port, REGISTERS_22_21_port, REGISTERS_22_20_port, 
      REGISTERS_22_19_port, REGISTERS_22_18_port, REGISTERS_22_17_port, 
      REGISTERS_22_16_port, REGISTERS_22_15_port, REGISTERS_22_14_port, 
      REGISTERS_22_13_port, REGISTERS_22_12_port, REGISTERS_22_11_port, 
      REGISTERS_22_10_port, REGISTERS_22_9_port, REGISTERS_22_8_port, 
      REGISTERS_22_7_port, REGISTERS_22_6_port, REGISTERS_22_5_port, 
      REGISTERS_22_4_port, REGISTERS_22_3_port, REGISTERS_22_2_port, 
      REGISTERS_22_1_port, REGISTERS_22_0_port, REGISTERS_23_31_port, 
      REGISTERS_23_30_port, REGISTERS_23_29_port, REGISTERS_23_28_port, 
      REGISTERS_23_27_port, REGISTERS_23_26_port, REGISTERS_23_25_port, 
      REGISTERS_23_24_port, REGISTERS_23_23_port, REGISTERS_23_22_port, 
      REGISTERS_23_21_port, REGISTERS_23_20_port, REGISTERS_23_19_port, 
      REGISTERS_23_18_port, REGISTERS_23_17_port, REGISTERS_23_16_port, 
      REGISTERS_23_15_port, REGISTERS_23_14_port, REGISTERS_23_13_port, 
      REGISTERS_23_12_port, REGISTERS_23_11_port, REGISTERS_23_10_port, 
      REGISTERS_23_9_port, REGISTERS_23_8_port, REGISTERS_23_7_port, 
      REGISTERS_23_6_port, REGISTERS_23_5_port, REGISTERS_23_4_port, 
      REGISTERS_23_3_port, REGISTERS_23_2_port, REGISTERS_23_1_port, 
      REGISTERS_23_0_port, REGISTERS_24_31_port, REGISTERS_24_30_port, 
      REGISTERS_24_29_port, REGISTERS_24_28_port, REGISTERS_24_27_port, 
      REGISTERS_24_26_port, REGISTERS_24_25_port, REGISTERS_24_24_port, 
      REGISTERS_24_23_port, REGISTERS_24_22_port, REGISTERS_24_21_port, 
      REGISTERS_24_20_port, REGISTERS_24_19_port, REGISTERS_24_18_port, 
      REGISTERS_24_17_port, REGISTERS_24_16_port, REGISTERS_24_15_port, 
      REGISTERS_24_14_port, REGISTERS_24_13_port, REGISTERS_24_12_port, 
      REGISTERS_24_11_port, REGISTERS_24_10_port, REGISTERS_24_9_port, 
      REGISTERS_24_8_port, REGISTERS_24_7_port, REGISTERS_24_6_port, 
      REGISTERS_24_5_port, REGISTERS_24_4_port, REGISTERS_24_3_port, 
      REGISTERS_24_2_port, REGISTERS_24_1_port, REGISTERS_24_0_port, 
      REGISTERS_25_31_port, REGISTERS_25_30_port, REGISTERS_25_29_port, 
      REGISTERS_25_28_port, REGISTERS_25_27_port, REGISTERS_25_26_port, 
      REGISTERS_25_25_port, REGISTERS_25_24_port, REGISTERS_25_23_port, 
      REGISTERS_25_22_port, REGISTERS_25_21_port, REGISTERS_25_20_port, 
      REGISTERS_25_19_port, REGISTERS_25_18_port, REGISTERS_25_17_port, 
      REGISTERS_25_16_port, REGISTERS_25_15_port, REGISTERS_25_14_port, 
      REGISTERS_25_13_port, REGISTERS_25_12_port, REGISTERS_25_11_port, 
      REGISTERS_25_10_port, REGISTERS_25_9_port, REGISTERS_25_8_port, 
      REGISTERS_25_7_port, REGISTERS_25_6_port, REGISTERS_25_5_port, 
      REGISTERS_25_4_port, REGISTERS_25_3_port, REGISTERS_25_2_port, 
      REGISTERS_25_1_port, REGISTERS_25_0_port, REGISTERS_26_31_port, 
      REGISTERS_26_30_port, REGISTERS_26_29_port, REGISTERS_26_28_port, 
      REGISTERS_26_27_port, REGISTERS_26_26_port, REGISTERS_26_25_port, 
      REGISTERS_26_24_port, REGISTERS_26_23_port, REGISTERS_26_22_port, 
      REGISTERS_26_21_port, REGISTERS_26_20_port, REGISTERS_26_19_port, 
      REGISTERS_26_18_port, REGISTERS_26_17_port, REGISTERS_26_16_port, 
      REGISTERS_26_15_port, REGISTERS_26_14_port, REGISTERS_26_13_port, 
      REGISTERS_26_12_port, REGISTERS_26_11_port, REGISTERS_26_10_port, 
      REGISTERS_26_9_port, REGISTERS_26_8_port, REGISTERS_26_7_port, 
      REGISTERS_26_6_port, REGISTERS_26_5_port, REGISTERS_26_4_port, 
      REGISTERS_26_3_port, REGISTERS_26_2_port, REGISTERS_26_1_port, 
      REGISTERS_26_0_port, REGISTERS_27_31_port, REGISTERS_27_30_port, 
      REGISTERS_27_29_port, REGISTERS_27_28_port, REGISTERS_27_27_port, 
      REGISTERS_27_26_port, REGISTERS_27_25_port, REGISTERS_27_24_port, 
      REGISTERS_27_23_port, REGISTERS_27_22_port, REGISTERS_27_21_port, 
      REGISTERS_27_20_port, REGISTERS_27_19_port, REGISTERS_27_18_port, 
      REGISTERS_27_17_port, REGISTERS_27_16_port, REGISTERS_27_15_port, 
      REGISTERS_27_14_port, REGISTERS_27_13_port, REGISTERS_27_12_port, 
      REGISTERS_27_11_port, REGISTERS_27_10_port, REGISTERS_27_9_port, 
      REGISTERS_27_8_port, REGISTERS_27_7_port, REGISTERS_27_6_port, 
      REGISTERS_27_5_port, REGISTERS_27_4_port, REGISTERS_27_3_port, 
      REGISTERS_27_2_port, REGISTERS_27_1_port, REGISTERS_27_0_port, 
      REGISTERS_28_31_port, REGISTERS_28_30_port, REGISTERS_28_29_port, 
      REGISTERS_28_28_port, REGISTERS_28_27_port, REGISTERS_28_26_port, 
      REGISTERS_28_25_port, REGISTERS_28_24_port, REGISTERS_28_23_port, 
      REGISTERS_28_22_port, REGISTERS_28_21_port, REGISTERS_28_20_port, 
      REGISTERS_28_19_port, REGISTERS_28_18_port, REGISTERS_28_17_port, 
      REGISTERS_28_16_port, REGISTERS_28_15_port, REGISTERS_28_14_port, 
      REGISTERS_28_13_port, REGISTERS_28_12_port, REGISTERS_28_11_port, 
      REGISTERS_28_10_port, REGISTERS_28_9_port, REGISTERS_28_8_port, 
      REGISTERS_28_7_port, REGISTERS_28_6_port, REGISTERS_28_5_port, 
      REGISTERS_28_4_port, REGISTERS_28_3_port, REGISTERS_28_2_port, 
      REGISTERS_28_1_port, REGISTERS_28_0_port, REGISTERS_29_31_port, 
      REGISTERS_29_30_port, REGISTERS_29_29_port, REGISTERS_29_28_port, 
      REGISTERS_29_27_port, REGISTERS_29_26_port, REGISTERS_29_25_port, 
      REGISTERS_29_24_port, REGISTERS_29_23_port, REGISTERS_29_22_port, 
      REGISTERS_29_21_port, REGISTERS_29_20_port, REGISTERS_29_19_port, 
      REGISTERS_29_18_port, REGISTERS_29_17_port, REGISTERS_29_16_port, 
      REGISTERS_29_15_port, REGISTERS_29_14_port, REGISTERS_29_13_port, 
      REGISTERS_29_12_port, REGISTERS_29_11_port, REGISTERS_29_10_port, 
      REGISTERS_29_9_port, REGISTERS_29_8_port, REGISTERS_29_7_port, 
      REGISTERS_29_6_port, REGISTERS_29_5_port, REGISTERS_29_4_port, 
      REGISTERS_29_3_port, REGISTERS_29_2_port, REGISTERS_29_1_port, 
      REGISTERS_29_0_port, REGISTERS_30_31_port, REGISTERS_30_30_port, 
      REGISTERS_30_29_port, REGISTERS_30_28_port, REGISTERS_30_27_port, 
      REGISTERS_30_26_port, REGISTERS_30_25_port, REGISTERS_30_24_port, 
      REGISTERS_30_23_port, REGISTERS_30_22_port, REGISTERS_30_21_port, 
      REGISTERS_30_20_port, REGISTERS_30_19_port, REGISTERS_30_18_port, 
      REGISTERS_30_17_port, REGISTERS_30_16_port, REGISTERS_30_15_port, 
      REGISTERS_30_14_port, REGISTERS_30_13_port, REGISTERS_30_12_port, 
      REGISTERS_30_11_port, REGISTERS_30_10_port, REGISTERS_30_9_port, 
      REGISTERS_30_8_port, REGISTERS_30_7_port, REGISTERS_30_6_port, 
      REGISTERS_30_5_port, REGISTERS_30_4_port, REGISTERS_30_3_port, 
      REGISTERS_30_2_port, REGISTERS_30_1_port, REGISTERS_30_0_port, 
      REGISTERS_31_31_port, REGISTERS_31_30_port, REGISTERS_31_29_port, 
      REGISTERS_31_28_port, REGISTERS_31_27_port, REGISTERS_31_26_port, 
      REGISTERS_31_25_port, REGISTERS_31_24_port, REGISTERS_31_23_port, 
      REGISTERS_31_22_port, REGISTERS_31_21_port, REGISTERS_31_20_port, 
      REGISTERS_31_19_port, REGISTERS_31_18_port, REGISTERS_31_17_port, 
      REGISTERS_31_16_port, REGISTERS_31_15_port, REGISTERS_31_14_port, 
      REGISTERS_31_13_port, REGISTERS_31_12_port, REGISTERS_31_11_port, 
      REGISTERS_31_10_port, REGISTERS_31_9_port, REGISTERS_31_8_port, 
      REGISTERS_31_7_port, REGISTERS_31_6_port, REGISTERS_31_5_port, 
      REGISTERS_31_4_port, REGISTERS_31_3_port, REGISTERS_31_2_port, 
      REGISTERS_31_1_port, REGISTERS_31_0_port, N2163, N2227, N2291, N2355, 
      N2419, N2483, N2547, N2611, N2675, N2739, N2803, N2867, N2931, N2995, 
      N3059, N3123, N3187, N3251, N3315, N3379, N3443, N3507, N3571, N3635, 
      N3699, N3763, N3827, N3891, N3955, N4019, N4083, N4086, N4088, N4090, 
      N4092, N4094, N4096, N4098, N4100, N4102, N4104, N4106, N4108, N4110, 
      N4112, N4114, N4116, N4118, N4120, N4122, N4124, N4126, N4128, N4130, 
      N4132, N4134, N4136, N4138, N4140, N4142, N4144, N4146, N4148, N4215, 
      N4216, N4217, N4218, N4219, N4220, N4221, N4222, N4223, N4224, N4225, 
      N4226, N4227, N4228, N4229, N4230, N4231, N4232, N4233, N4234, N4235, 
      N4236, N4237, N4238, N4239, N4240, N4241, N4242, N4243, N4244, N4245, 
      N4246, N4278, N4344, N4345, N4346, N4347, N4348, N4349, N4350, N4351, 
      N4352, N4353, N4354, N4355, N4356, N4357, N4358, N4359, N4360, N4361, 
      N4362, N4363, N4364, N4365, N4366, N4367, N4368, N4369, N4370, N4371, 
      N4372, N4373, N4374, N4375, N4407, n2, n3, n4, n5, n6, n7, n8, n9, n10, 
      n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25
      , n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, 
      n40, n41, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56
      , n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, 
      n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85
      , n86, n87, n88, n89, n90, n92, n93, n94, n95, n96, n97, n98, n99, n100, 
      n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, 
      n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, 
      n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, 
      n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n160, n161, n162, 
      n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, 
      n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, 
      n187, n188, n189, n190, n191, n192, n194, n195, n196, n197, n198, n199, 
      n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
      n224, n225, n226, n228, n229, n230, n231, n232, n233, n234, n235, n236, 
      n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, 
      n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, 
      n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, 
      n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, 
      n286, n287, n288, n289, n290, n291, n292, n293, n294, n296, n297, n298, 
      n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, 
      n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, 
      n323, n324, n325, n326, n327, n328, n330, n331, n332, n333, n334, n335, 
      n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, 
      n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, 
      n360, n361, n362, n364, n365, n366, n367, n368, n369, n370, n371, n372, 
      n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, 
      n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, 
      n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, 
      n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, 
      n422, n423, n424, n425, n426, n427, n428, n429, n430, n432, n433, n434, 
      n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, 
      n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, 
      n459, n460, n461, n462, n463, n464, n466, n467, n468, n469, n470, n471, 
      n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, 
      n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, 
      n496, n497, n498, n500, n501, n502, n503, n504, n505, n506, n507, n508, 
      n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, 
      n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, 
      n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, 
      n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, 
      n558, n559, n560, n561, n562, n563, n564, n565, n566, n568, n569, n570, 
      n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, 
      n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, 
      n595, n596, n597, n598, n599, n600, n602, n603, n604, n605, n606, n607, 
      n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, 
      n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, 
      n632, n633, n634, n636, n637, n638, n639, n640, n641, n642, n643, n644, 
      n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, 
      n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, 
      n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, 
      n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, 
      n694, n695, n696, n697, n698, n699, n700, n701, n702, n704, n705, n706, 
      n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, 
      n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, 
      n731, n732, n733, n734, n735, n736, n738, n739, n740, n741, n742, n743, 
      n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, 
      n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, 
      n768, n769, n770, n772, n773, n774, n775, n776, n777, n778, n779, n780, 
      n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, 
      n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, 
      n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, 
      n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, 
      n830, n831, n832, n833, n834, n835, n836, n837, n838, n840, n841, n842, 
      n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, 
      n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, 
      n867, n868, n869, n870, n871, n872, n874, n875, n876, n877, n878, n879, 
      n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, 
      n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, 
      n904, n905, n906, n908, n909, n910, n911, n912, n913, n914, n915, n916, 
      n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, 
      n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, 
      n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, 
      n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, 
      n966, n967, n968, n969, n970, n971, n972, n973, n974, n976, n977, n978, 
      n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, 
      n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002
      , n1003, n1004, n1005, n1006, n1007, n1008, n1010, n1011, n1012, n1013, 
      n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, 
      n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, 
      n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1044, 
      n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, 
      n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, 
      n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, 
      n1075, n1076, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, 
      n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, 
      n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, 
      n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, 
      n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1124, n1125, n1126, 
      n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, 
      n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, 
      n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, 
      n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, 
      n1167, n1168, n1169, n1170, n1171, n1172, n1174, n1175, n1176, n1177, 
      n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, 
      n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, 
      n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, 
      n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, 
      n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, 
      n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, 
      n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, 
      n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, 
      n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, 
      n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, 
      n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, 
      n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, 
      n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, 
      n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, 
      n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, 
      n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, 
      n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, 
      n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, 
      n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, 
      n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, 
      n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, 
      n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, 
      n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, 
      n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, 
      n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, 
      n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, 
      n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, 
      n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, 
      n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, 
      n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, 
      n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, 
      n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, 
      n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, 
      n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, 
      n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, 
      n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, 
      n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, 
      n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, 
      n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, 
      n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, 
      n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, 
      n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, 
      n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, 
      n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, 
      n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, 
      n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, 
      n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, 
      n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, 
      n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, 
      n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, 
      n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, 
      n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, 
      n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, 
      n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, 
      n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, 
      n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, 
      n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, 
      n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, 
      n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, 
      n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, 
      n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, 
      n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, 
      n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, 
      n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1,
      n193, n227, n261, n295, n329 : std_logic;

begin
   
   REGISTERS_reg_1_31_inst : DLH_X1 port map( G => N4083, D => N4148, Q => 
                           REGISTERS_1_31_port);
   REGISTERS_reg_1_30_inst : DLH_X1 port map( G => N4083, D => N4146, Q => 
                           REGISTERS_1_30_port);
   REGISTERS_reg_1_29_inst : DLH_X1 port map( G => N4083, D => N4144, Q => 
                           REGISTERS_1_29_port);
   REGISTERS_reg_1_28_inst : DLH_X1 port map( G => N4083, D => N4142, Q => 
                           REGISTERS_1_28_port);
   REGISTERS_reg_1_27_inst : DLH_X1 port map( G => N4083, D => N4140, Q => 
                           REGISTERS_1_27_port);
   REGISTERS_reg_1_26_inst : DLH_X1 port map( G => N4083, D => N4138, Q => 
                           REGISTERS_1_26_port);
   REGISTERS_reg_1_25_inst : DLH_X1 port map( G => N4083, D => N4136, Q => 
                           REGISTERS_1_25_port);
   REGISTERS_reg_1_24_inst : DLH_X1 port map( G => N4083, D => N4134, Q => 
                           REGISTERS_1_24_port);
   REGISTERS_reg_1_23_inst : DLH_X1 port map( G => N4083, D => N4132, Q => 
                           REGISTERS_1_23_port);
   REGISTERS_reg_1_22_inst : DLH_X1 port map( G => N4083, D => N4130, Q => 
                           REGISTERS_1_22_port);
   REGISTERS_reg_1_21_inst : DLH_X1 port map( G => N4083, D => N4128, Q => 
                           REGISTERS_1_21_port);
   REGISTERS_reg_1_20_inst : DLH_X1 port map( G => N4083, D => N4126, Q => 
                           REGISTERS_1_20_port);
   REGISTERS_reg_1_19_inst : DLH_X1 port map( G => N4083, D => N4124, Q => 
                           REGISTERS_1_19_port);
   REGISTERS_reg_1_18_inst : DLH_X1 port map( G => N4083, D => N4122, Q => 
                           REGISTERS_1_18_port);
   REGISTERS_reg_1_17_inst : DLH_X1 port map( G => N4083, D => N4120, Q => 
                           REGISTERS_1_17_port);
   REGISTERS_reg_1_16_inst : DLH_X1 port map( G => N4083, D => N4118, Q => 
                           REGISTERS_1_16_port);
   REGISTERS_reg_1_15_inst : DLH_X1 port map( G => N4083, D => N4116, Q => 
                           REGISTERS_1_15_port);
   REGISTERS_reg_1_14_inst : DLH_X1 port map( G => N4083, D => N4114, Q => 
                           REGISTERS_1_14_port);
   REGISTERS_reg_1_13_inst : DLH_X1 port map( G => N4083, D => N4112, Q => 
                           REGISTERS_1_13_port);
   REGISTERS_reg_1_12_inst : DLH_X1 port map( G => N4083, D => N4110, Q => 
                           REGISTERS_1_12_port);
   REGISTERS_reg_1_11_inst : DLH_X1 port map( G => N4083, D => N4108, Q => 
                           REGISTERS_1_11_port);
   REGISTERS_reg_1_10_inst : DLH_X1 port map( G => N4083, D => N4106, Q => 
                           REGISTERS_1_10_port);
   REGISTERS_reg_1_9_inst : DLH_X1 port map( G => N4083, D => N4104, Q => 
                           REGISTERS_1_9_port);
   REGISTERS_reg_1_8_inst : DLH_X1 port map( G => N4083, D => N4102, Q => 
                           REGISTERS_1_8_port);
   REGISTERS_reg_1_7_inst : DLH_X1 port map( G => N4083, D => N4100, Q => 
                           REGISTERS_1_7_port);
   REGISTERS_reg_1_6_inst : DLH_X1 port map( G => N4083, D => N4098, Q => 
                           REGISTERS_1_6_port);
   REGISTERS_reg_1_5_inst : DLH_X1 port map( G => N4083, D => N4096, Q => 
                           REGISTERS_1_5_port);
   REGISTERS_reg_1_4_inst : DLH_X1 port map( G => N4083, D => N4094, Q => 
                           REGISTERS_1_4_port);
   REGISTERS_reg_1_3_inst : DLH_X1 port map( G => N4083, D => N4092, Q => 
                           REGISTERS_1_3_port);
   REGISTERS_reg_1_2_inst : DLH_X1 port map( G => N4083, D => N4090, Q => 
                           REGISTERS_1_2_port);
   REGISTERS_reg_1_1_inst : DLH_X1 port map( G => N4083, D => N4088, Q => 
                           REGISTERS_1_1_port);
   REGISTERS_reg_1_0_inst : DLH_X1 port map( G => N4083, D => N4086, Q => 
                           REGISTERS_1_0_port);
   REGISTERS_reg_2_31_inst : DLH_X1 port map( G => N4019, D => N4148, Q => 
                           REGISTERS_2_31_port);
   REGISTERS_reg_2_30_inst : DLH_X1 port map( G => N4019, D => N4146, Q => 
                           REGISTERS_2_30_port);
   REGISTERS_reg_2_29_inst : DLH_X1 port map( G => N4019, D => N4144, Q => 
                           REGISTERS_2_29_port);
   REGISTERS_reg_2_28_inst : DLH_X1 port map( G => N4019, D => N4142, Q => 
                           REGISTERS_2_28_port);
   REGISTERS_reg_2_27_inst : DLH_X1 port map( G => N4019, D => N4140, Q => 
                           REGISTERS_2_27_port);
   REGISTERS_reg_2_26_inst : DLH_X1 port map( G => N4019, D => N4138, Q => 
                           REGISTERS_2_26_port);
   REGISTERS_reg_2_25_inst : DLH_X1 port map( G => N4019, D => N4136, Q => 
                           REGISTERS_2_25_port);
   REGISTERS_reg_2_24_inst : DLH_X1 port map( G => N4019, D => N4134, Q => 
                           REGISTERS_2_24_port);
   REGISTERS_reg_2_23_inst : DLH_X1 port map( G => N4019, D => N4132, Q => 
                           REGISTERS_2_23_port);
   REGISTERS_reg_2_22_inst : DLH_X1 port map( G => N4019, D => N4130, Q => 
                           REGISTERS_2_22_port);
   REGISTERS_reg_2_21_inst : DLH_X1 port map( G => N4019, D => N4128, Q => 
                           REGISTERS_2_21_port);
   REGISTERS_reg_2_20_inst : DLH_X1 port map( G => N4019, D => N4126, Q => 
                           REGISTERS_2_20_port);
   REGISTERS_reg_2_19_inst : DLH_X1 port map( G => N4019, D => N4124, Q => 
                           REGISTERS_2_19_port);
   REGISTERS_reg_2_18_inst : DLH_X1 port map( G => N4019, D => N4122, Q => 
                           REGISTERS_2_18_port);
   REGISTERS_reg_2_17_inst : DLH_X1 port map( G => N4019, D => N4120, Q => 
                           REGISTERS_2_17_port);
   REGISTERS_reg_2_16_inst : DLH_X1 port map( G => N4019, D => N4118, Q => 
                           REGISTERS_2_16_port);
   REGISTERS_reg_2_15_inst : DLH_X1 port map( G => N4019, D => N4116, Q => 
                           REGISTERS_2_15_port);
   REGISTERS_reg_2_14_inst : DLH_X1 port map( G => N4019, D => N4114, Q => 
                           REGISTERS_2_14_port);
   REGISTERS_reg_2_13_inst : DLH_X1 port map( G => N4019, D => N4112, Q => 
                           REGISTERS_2_13_port);
   REGISTERS_reg_2_12_inst : DLH_X1 port map( G => N4019, D => N4110, Q => 
                           REGISTERS_2_12_port);
   REGISTERS_reg_2_11_inst : DLH_X1 port map( G => N4019, D => N4108, Q => 
                           REGISTERS_2_11_port);
   REGISTERS_reg_2_10_inst : DLH_X1 port map( G => N4019, D => N4106, Q => 
                           REGISTERS_2_10_port);
   REGISTERS_reg_2_9_inst : DLH_X1 port map( G => N4019, D => N4104, Q => 
                           REGISTERS_2_9_port);
   REGISTERS_reg_2_8_inst : DLH_X1 port map( G => N4019, D => N4102, Q => 
                           REGISTERS_2_8_port);
   REGISTERS_reg_2_7_inst : DLH_X1 port map( G => N4019, D => N4100, Q => 
                           REGISTERS_2_7_port);
   REGISTERS_reg_2_6_inst : DLH_X1 port map( G => N4019, D => N4098, Q => 
                           REGISTERS_2_6_port);
   REGISTERS_reg_2_5_inst : DLH_X1 port map( G => N4019, D => N4096, Q => 
                           REGISTERS_2_5_port);
   REGISTERS_reg_2_4_inst : DLH_X1 port map( G => N4019, D => N4094, Q => 
                           REGISTERS_2_4_port);
   REGISTERS_reg_2_3_inst : DLH_X1 port map( G => N4019, D => N4092, Q => 
                           REGISTERS_2_3_port);
   REGISTERS_reg_2_2_inst : DLH_X1 port map( G => N4019, D => N4090, Q => 
                           REGISTERS_2_2_port);
   REGISTERS_reg_2_1_inst : DLH_X1 port map( G => N4019, D => N4088, Q => 
                           REGISTERS_2_1_port);
   REGISTERS_reg_2_0_inst : DLH_X1 port map( G => N4019, D => N4086, Q => 
                           REGISTERS_2_0_port);
   REGISTERS_reg_3_31_inst : DLH_X1 port map( G => N3955, D => N4148, Q => 
                           REGISTERS_3_31_port);
   REGISTERS_reg_3_30_inst : DLH_X1 port map( G => N3955, D => N4146, Q => 
                           REGISTERS_3_30_port);
   REGISTERS_reg_3_29_inst : DLH_X1 port map( G => N3955, D => N4144, Q => 
                           REGISTERS_3_29_port);
   REGISTERS_reg_3_28_inst : DLH_X1 port map( G => N3955, D => N4142, Q => 
                           REGISTERS_3_28_port);
   REGISTERS_reg_3_27_inst : DLH_X1 port map( G => N3955, D => N4140, Q => 
                           REGISTERS_3_27_port);
   REGISTERS_reg_3_26_inst : DLH_X1 port map( G => N3955, D => N4138, Q => 
                           REGISTERS_3_26_port);
   REGISTERS_reg_3_25_inst : DLH_X1 port map( G => N3955, D => N4136, Q => 
                           REGISTERS_3_25_port);
   REGISTERS_reg_3_24_inst : DLH_X1 port map( G => N3955, D => N4134, Q => 
                           REGISTERS_3_24_port);
   REGISTERS_reg_3_23_inst : DLH_X1 port map( G => N3955, D => N4132, Q => 
                           REGISTERS_3_23_port);
   REGISTERS_reg_3_22_inst : DLH_X1 port map( G => N3955, D => N4130, Q => 
                           REGISTERS_3_22_port);
   REGISTERS_reg_3_21_inst : DLH_X1 port map( G => N3955, D => N4128, Q => 
                           REGISTERS_3_21_port);
   REGISTERS_reg_3_20_inst : DLH_X1 port map( G => N3955, D => N4126, Q => 
                           REGISTERS_3_20_port);
   REGISTERS_reg_3_19_inst : DLH_X1 port map( G => N3955, D => N4124, Q => 
                           REGISTERS_3_19_port);
   REGISTERS_reg_3_18_inst : DLH_X1 port map( G => N3955, D => N4122, Q => 
                           REGISTERS_3_18_port);
   REGISTERS_reg_3_17_inst : DLH_X1 port map( G => N3955, D => N4120, Q => 
                           REGISTERS_3_17_port);
   REGISTERS_reg_3_16_inst : DLH_X1 port map( G => N3955, D => N4118, Q => 
                           REGISTERS_3_16_port);
   REGISTERS_reg_3_15_inst : DLH_X1 port map( G => N3955, D => N4116, Q => 
                           REGISTERS_3_15_port);
   REGISTERS_reg_3_14_inst : DLH_X1 port map( G => N3955, D => N4114, Q => 
                           REGISTERS_3_14_port);
   REGISTERS_reg_3_13_inst : DLH_X1 port map( G => N3955, D => N4112, Q => 
                           REGISTERS_3_13_port);
   REGISTERS_reg_3_12_inst : DLH_X1 port map( G => N3955, D => N4110, Q => 
                           REGISTERS_3_12_port);
   REGISTERS_reg_3_11_inst : DLH_X1 port map( G => N3955, D => N4108, Q => 
                           REGISTERS_3_11_port);
   REGISTERS_reg_3_10_inst : DLH_X1 port map( G => N3955, D => N4106, Q => 
                           REGISTERS_3_10_port);
   REGISTERS_reg_3_9_inst : DLH_X1 port map( G => N3955, D => N4104, Q => 
                           REGISTERS_3_9_port);
   REGISTERS_reg_3_8_inst : DLH_X1 port map( G => N3955, D => N4102, Q => 
                           REGISTERS_3_8_port);
   REGISTERS_reg_3_7_inst : DLH_X1 port map( G => N3955, D => N4100, Q => 
                           REGISTERS_3_7_port);
   REGISTERS_reg_3_6_inst : DLH_X1 port map( G => N3955, D => N4098, Q => 
                           REGISTERS_3_6_port);
   REGISTERS_reg_3_5_inst : DLH_X1 port map( G => N3955, D => N4096, Q => 
                           REGISTERS_3_5_port);
   REGISTERS_reg_3_4_inst : DLH_X1 port map( G => N3955, D => N4094, Q => 
                           REGISTERS_3_4_port);
   REGISTERS_reg_3_3_inst : DLH_X1 port map( G => N3955, D => N4092, Q => 
                           REGISTERS_3_3_port);
   REGISTERS_reg_3_2_inst : DLH_X1 port map( G => N3955, D => N4090, Q => 
                           REGISTERS_3_2_port);
   REGISTERS_reg_3_1_inst : DLH_X1 port map( G => N3955, D => N4088, Q => 
                           REGISTERS_3_1_port);
   REGISTERS_reg_3_0_inst : DLH_X1 port map( G => N3955, D => N4086, Q => 
                           REGISTERS_3_0_port);
   REGISTERS_reg_4_31_inst : DLH_X1 port map( G => N3891, D => N4148, Q => 
                           REGISTERS_4_31_port);
   REGISTERS_reg_4_30_inst : DLH_X1 port map( G => N3891, D => N4146, Q => 
                           REGISTERS_4_30_port);
   REGISTERS_reg_4_29_inst : DLH_X1 port map( G => N3891, D => N4144, Q => 
                           REGISTERS_4_29_port);
   REGISTERS_reg_4_28_inst : DLH_X1 port map( G => N3891, D => N4142, Q => 
                           REGISTERS_4_28_port);
   REGISTERS_reg_4_27_inst : DLH_X1 port map( G => N3891, D => N4140, Q => 
                           REGISTERS_4_27_port);
   REGISTERS_reg_4_26_inst : DLH_X1 port map( G => N3891, D => N4138, Q => 
                           REGISTERS_4_26_port);
   REGISTERS_reg_4_25_inst : DLH_X1 port map( G => N3891, D => N4136, Q => 
                           REGISTERS_4_25_port);
   REGISTERS_reg_4_24_inst : DLH_X1 port map( G => N3891, D => N4134, Q => 
                           REGISTERS_4_24_port);
   REGISTERS_reg_4_23_inst : DLH_X1 port map( G => N3891, D => N4132, Q => 
                           REGISTERS_4_23_port);
   REGISTERS_reg_4_22_inst : DLH_X1 port map( G => N3891, D => N4130, Q => 
                           REGISTERS_4_22_port);
   REGISTERS_reg_4_21_inst : DLH_X1 port map( G => N3891, D => N4128, Q => 
                           REGISTERS_4_21_port);
   REGISTERS_reg_4_20_inst : DLH_X1 port map( G => N3891, D => N4126, Q => 
                           REGISTERS_4_20_port);
   REGISTERS_reg_4_19_inst : DLH_X1 port map( G => N3891, D => N4124, Q => 
                           REGISTERS_4_19_port);
   REGISTERS_reg_4_18_inst : DLH_X1 port map( G => N3891, D => N4122, Q => 
                           REGISTERS_4_18_port);
   REGISTERS_reg_4_17_inst : DLH_X1 port map( G => N3891, D => N4120, Q => 
                           REGISTERS_4_17_port);
   REGISTERS_reg_4_16_inst : DLH_X1 port map( G => N3891, D => N4118, Q => 
                           REGISTERS_4_16_port);
   REGISTERS_reg_4_15_inst : DLH_X1 port map( G => N3891, D => N4116, Q => 
                           REGISTERS_4_15_port);
   REGISTERS_reg_4_14_inst : DLH_X1 port map( G => N3891, D => N4114, Q => 
                           REGISTERS_4_14_port);
   REGISTERS_reg_4_13_inst : DLH_X1 port map( G => N3891, D => N4112, Q => 
                           REGISTERS_4_13_port);
   REGISTERS_reg_4_12_inst : DLH_X1 port map( G => N3891, D => N4110, Q => 
                           REGISTERS_4_12_port);
   REGISTERS_reg_4_11_inst : DLH_X1 port map( G => N3891, D => N4108, Q => 
                           REGISTERS_4_11_port);
   REGISTERS_reg_4_10_inst : DLH_X1 port map( G => N3891, D => N4106, Q => 
                           REGISTERS_4_10_port);
   REGISTERS_reg_4_9_inst : DLH_X1 port map( G => N3891, D => N4104, Q => 
                           REGISTERS_4_9_port);
   REGISTERS_reg_4_8_inst : DLH_X1 port map( G => N3891, D => N4102, Q => 
                           REGISTERS_4_8_port);
   REGISTERS_reg_4_7_inst : DLH_X1 port map( G => N3891, D => N4100, Q => 
                           REGISTERS_4_7_port);
   REGISTERS_reg_4_6_inst : DLH_X1 port map( G => N3891, D => N4098, Q => 
                           REGISTERS_4_6_port);
   REGISTERS_reg_4_5_inst : DLH_X1 port map( G => N3891, D => N4096, Q => 
                           REGISTERS_4_5_port);
   REGISTERS_reg_4_4_inst : DLH_X1 port map( G => N3891, D => N4094, Q => 
                           REGISTERS_4_4_port);
   REGISTERS_reg_4_3_inst : DLH_X1 port map( G => N3891, D => N4092, Q => 
                           REGISTERS_4_3_port);
   REGISTERS_reg_4_2_inst : DLH_X1 port map( G => N3891, D => N4090, Q => 
                           REGISTERS_4_2_port);
   REGISTERS_reg_4_1_inst : DLH_X1 port map( G => N3891, D => N4088, Q => 
                           REGISTERS_4_1_port);
   REGISTERS_reg_4_0_inst : DLH_X1 port map( G => N3891, D => N4086, Q => 
                           REGISTERS_4_0_port);
   REGISTERS_reg_5_31_inst : DLH_X1 port map( G => N3827, D => N4148, Q => 
                           REGISTERS_5_31_port);
   REGISTERS_reg_5_30_inst : DLH_X1 port map( G => N3827, D => N4146, Q => 
                           REGISTERS_5_30_port);
   REGISTERS_reg_5_29_inst : DLH_X1 port map( G => N3827, D => N4144, Q => 
                           REGISTERS_5_29_port);
   REGISTERS_reg_5_28_inst : DLH_X1 port map( G => N3827, D => N4142, Q => 
                           REGISTERS_5_28_port);
   REGISTERS_reg_5_27_inst : DLH_X1 port map( G => N3827, D => N4140, Q => 
                           REGISTERS_5_27_port);
   REGISTERS_reg_5_26_inst : DLH_X1 port map( G => N3827, D => N4138, Q => 
                           REGISTERS_5_26_port);
   REGISTERS_reg_5_25_inst : DLH_X1 port map( G => N3827, D => N4136, Q => 
                           REGISTERS_5_25_port);
   REGISTERS_reg_5_24_inst : DLH_X1 port map( G => N3827, D => N4134, Q => 
                           REGISTERS_5_24_port);
   REGISTERS_reg_5_23_inst : DLH_X1 port map( G => N3827, D => N4132, Q => 
                           REGISTERS_5_23_port);
   REGISTERS_reg_5_22_inst : DLH_X1 port map( G => N3827, D => N4130, Q => 
                           REGISTERS_5_22_port);
   REGISTERS_reg_5_21_inst : DLH_X1 port map( G => N3827, D => N4128, Q => 
                           REGISTERS_5_21_port);
   REGISTERS_reg_5_20_inst : DLH_X1 port map( G => N3827, D => N4126, Q => 
                           REGISTERS_5_20_port);
   REGISTERS_reg_5_19_inst : DLH_X1 port map( G => N3827, D => N4124, Q => 
                           REGISTERS_5_19_port);
   REGISTERS_reg_5_18_inst : DLH_X1 port map( G => N3827, D => N4122, Q => 
                           REGISTERS_5_18_port);
   REGISTERS_reg_5_17_inst : DLH_X1 port map( G => N3827, D => N4120, Q => 
                           REGISTERS_5_17_port);
   REGISTERS_reg_5_16_inst : DLH_X1 port map( G => N3827, D => N4118, Q => 
                           REGISTERS_5_16_port);
   REGISTERS_reg_5_15_inst : DLH_X1 port map( G => N3827, D => N4116, Q => 
                           REGISTERS_5_15_port);
   REGISTERS_reg_5_14_inst : DLH_X1 port map( G => N3827, D => N4114, Q => 
                           REGISTERS_5_14_port);
   REGISTERS_reg_5_13_inst : DLH_X1 port map( G => N3827, D => N4112, Q => 
                           REGISTERS_5_13_port);
   REGISTERS_reg_5_12_inst : DLH_X1 port map( G => N3827, D => N4110, Q => 
                           REGISTERS_5_12_port);
   REGISTERS_reg_5_11_inst : DLH_X1 port map( G => N3827, D => N4108, Q => 
                           REGISTERS_5_11_port);
   REGISTERS_reg_5_10_inst : DLH_X1 port map( G => N3827, D => N4106, Q => 
                           REGISTERS_5_10_port);
   REGISTERS_reg_5_9_inst : DLH_X1 port map( G => N3827, D => N4104, Q => 
                           REGISTERS_5_9_port);
   REGISTERS_reg_5_8_inst : DLH_X1 port map( G => N3827, D => N4102, Q => 
                           REGISTERS_5_8_port);
   REGISTERS_reg_5_7_inst : DLH_X1 port map( G => N3827, D => N4100, Q => 
                           REGISTERS_5_7_port);
   REGISTERS_reg_5_6_inst : DLH_X1 port map( G => N3827, D => N4098, Q => 
                           REGISTERS_5_6_port);
   REGISTERS_reg_5_5_inst : DLH_X1 port map( G => N3827, D => N4096, Q => 
                           REGISTERS_5_5_port);
   REGISTERS_reg_5_4_inst : DLH_X1 port map( G => N3827, D => N4094, Q => 
                           REGISTERS_5_4_port);
   REGISTERS_reg_5_3_inst : DLH_X1 port map( G => N3827, D => N4092, Q => 
                           REGISTERS_5_3_port);
   REGISTERS_reg_5_2_inst : DLH_X1 port map( G => N3827, D => N4090, Q => 
                           REGISTERS_5_2_port);
   REGISTERS_reg_5_1_inst : DLH_X1 port map( G => N3827, D => N4088, Q => 
                           REGISTERS_5_1_port);
   REGISTERS_reg_5_0_inst : DLH_X1 port map( G => N3827, D => N4086, Q => 
                           REGISTERS_5_0_port);
   REGISTERS_reg_6_31_inst : DLH_X1 port map( G => N3763, D => N4148, Q => 
                           REGISTERS_6_31_port);
   REGISTERS_reg_6_30_inst : DLH_X1 port map( G => N3763, D => N4146, Q => 
                           REGISTERS_6_30_port);
   REGISTERS_reg_6_29_inst : DLH_X1 port map( G => N3763, D => N4144, Q => 
                           REGISTERS_6_29_port);
   REGISTERS_reg_6_28_inst : DLH_X1 port map( G => N3763, D => N4142, Q => 
                           REGISTERS_6_28_port);
   REGISTERS_reg_6_27_inst : DLH_X1 port map( G => N3763, D => N4140, Q => 
                           REGISTERS_6_27_port);
   REGISTERS_reg_6_26_inst : DLH_X1 port map( G => N3763, D => N4138, Q => 
                           REGISTERS_6_26_port);
   REGISTERS_reg_6_25_inst : DLH_X1 port map( G => N3763, D => N4136, Q => 
                           REGISTERS_6_25_port);
   REGISTERS_reg_6_24_inst : DLH_X1 port map( G => N3763, D => N4134, Q => 
                           REGISTERS_6_24_port);
   REGISTERS_reg_6_23_inst : DLH_X1 port map( G => N3763, D => N4132, Q => 
                           REGISTERS_6_23_port);
   REGISTERS_reg_6_22_inst : DLH_X1 port map( G => N3763, D => N4130, Q => 
                           REGISTERS_6_22_port);
   REGISTERS_reg_6_21_inst : DLH_X1 port map( G => N3763, D => N4128, Q => 
                           REGISTERS_6_21_port);
   REGISTERS_reg_6_20_inst : DLH_X1 port map( G => N3763, D => N4126, Q => 
                           REGISTERS_6_20_port);
   REGISTERS_reg_6_19_inst : DLH_X1 port map( G => N3763, D => N4124, Q => 
                           REGISTERS_6_19_port);
   REGISTERS_reg_6_18_inst : DLH_X1 port map( G => N3763, D => N4122, Q => 
                           REGISTERS_6_18_port);
   REGISTERS_reg_6_17_inst : DLH_X1 port map( G => N3763, D => N4120, Q => 
                           REGISTERS_6_17_port);
   REGISTERS_reg_6_16_inst : DLH_X1 port map( G => N3763, D => N4118, Q => 
                           REGISTERS_6_16_port);
   REGISTERS_reg_6_15_inst : DLH_X1 port map( G => N3763, D => N4116, Q => 
                           REGISTERS_6_15_port);
   REGISTERS_reg_6_14_inst : DLH_X1 port map( G => N3763, D => N4114, Q => 
                           REGISTERS_6_14_port);
   REGISTERS_reg_6_13_inst : DLH_X1 port map( G => N3763, D => N4112, Q => 
                           REGISTERS_6_13_port);
   REGISTERS_reg_6_12_inst : DLH_X1 port map( G => N3763, D => N4110, Q => 
                           REGISTERS_6_12_port);
   REGISTERS_reg_6_11_inst : DLH_X1 port map( G => N3763, D => N4108, Q => 
                           REGISTERS_6_11_port);
   REGISTERS_reg_6_10_inst : DLH_X1 port map( G => N3763, D => N4106, Q => 
                           REGISTERS_6_10_port);
   REGISTERS_reg_6_9_inst : DLH_X1 port map( G => N3763, D => N4104, Q => 
                           REGISTERS_6_9_port);
   REGISTERS_reg_6_8_inst : DLH_X1 port map( G => N3763, D => N4102, Q => 
                           REGISTERS_6_8_port);
   REGISTERS_reg_6_7_inst : DLH_X1 port map( G => N3763, D => N4100, Q => 
                           REGISTERS_6_7_port);
   REGISTERS_reg_6_6_inst : DLH_X1 port map( G => N3763, D => N4098, Q => 
                           REGISTERS_6_6_port);
   REGISTERS_reg_6_5_inst : DLH_X1 port map( G => N3763, D => N4096, Q => 
                           REGISTERS_6_5_port);
   REGISTERS_reg_6_4_inst : DLH_X1 port map( G => N3763, D => N4094, Q => 
                           REGISTERS_6_4_port);
   REGISTERS_reg_6_3_inst : DLH_X1 port map( G => N3763, D => N4092, Q => 
                           REGISTERS_6_3_port);
   REGISTERS_reg_6_2_inst : DLH_X1 port map( G => N3763, D => N4090, Q => 
                           REGISTERS_6_2_port);
   REGISTERS_reg_6_1_inst : DLH_X1 port map( G => N3763, D => N4088, Q => 
                           REGISTERS_6_1_port);
   REGISTERS_reg_6_0_inst : DLH_X1 port map( G => N3763, D => N4086, Q => 
                           REGISTERS_6_0_port);
   REGISTERS_reg_7_31_inst : DLH_X1 port map( G => N3699, D => N4148, Q => 
                           REGISTERS_7_31_port);
   REGISTERS_reg_7_30_inst : DLH_X1 port map( G => N3699, D => N4146, Q => 
                           REGISTERS_7_30_port);
   REGISTERS_reg_7_29_inst : DLH_X1 port map( G => N3699, D => N4144, Q => 
                           REGISTERS_7_29_port);
   REGISTERS_reg_7_28_inst : DLH_X1 port map( G => N3699, D => N4142, Q => 
                           REGISTERS_7_28_port);
   REGISTERS_reg_7_27_inst : DLH_X1 port map( G => N3699, D => N4140, Q => 
                           REGISTERS_7_27_port);
   REGISTERS_reg_7_26_inst : DLH_X1 port map( G => N3699, D => N4138, Q => 
                           REGISTERS_7_26_port);
   REGISTERS_reg_7_25_inst : DLH_X1 port map( G => N3699, D => N4136, Q => 
                           REGISTERS_7_25_port);
   REGISTERS_reg_7_24_inst : DLH_X1 port map( G => N3699, D => N4134, Q => 
                           REGISTERS_7_24_port);
   REGISTERS_reg_7_23_inst : DLH_X1 port map( G => N3699, D => N4132, Q => 
                           REGISTERS_7_23_port);
   REGISTERS_reg_7_22_inst : DLH_X1 port map( G => N3699, D => N4130, Q => 
                           REGISTERS_7_22_port);
   REGISTERS_reg_7_21_inst : DLH_X1 port map( G => N3699, D => N4128, Q => 
                           REGISTERS_7_21_port);
   REGISTERS_reg_7_20_inst : DLH_X1 port map( G => N3699, D => N4126, Q => 
                           REGISTERS_7_20_port);
   REGISTERS_reg_7_19_inst : DLH_X1 port map( G => N3699, D => N4124, Q => 
                           REGISTERS_7_19_port);
   REGISTERS_reg_7_18_inst : DLH_X1 port map( G => N3699, D => N4122, Q => 
                           REGISTERS_7_18_port);
   REGISTERS_reg_7_17_inst : DLH_X1 port map( G => N3699, D => N4120, Q => 
                           REGISTERS_7_17_port);
   REGISTERS_reg_7_16_inst : DLH_X1 port map( G => N3699, D => N4118, Q => 
                           REGISTERS_7_16_port);
   REGISTERS_reg_7_15_inst : DLH_X1 port map( G => N3699, D => N4116, Q => 
                           REGISTERS_7_15_port);
   REGISTERS_reg_7_14_inst : DLH_X1 port map( G => N3699, D => N4114, Q => 
                           REGISTERS_7_14_port);
   REGISTERS_reg_7_13_inst : DLH_X1 port map( G => N3699, D => N4112, Q => 
                           REGISTERS_7_13_port);
   REGISTERS_reg_7_12_inst : DLH_X1 port map( G => N3699, D => N4110, Q => 
                           REGISTERS_7_12_port);
   REGISTERS_reg_7_11_inst : DLH_X1 port map( G => N3699, D => N4108, Q => 
                           REGISTERS_7_11_port);
   REGISTERS_reg_7_10_inst : DLH_X1 port map( G => N3699, D => N4106, Q => 
                           REGISTERS_7_10_port);
   REGISTERS_reg_7_9_inst : DLH_X1 port map( G => N3699, D => N4104, Q => 
                           REGISTERS_7_9_port);
   REGISTERS_reg_7_8_inst : DLH_X1 port map( G => N3699, D => N4102, Q => 
                           REGISTERS_7_8_port);
   REGISTERS_reg_7_7_inst : DLH_X1 port map( G => N3699, D => N4100, Q => 
                           REGISTERS_7_7_port);
   REGISTERS_reg_7_6_inst : DLH_X1 port map( G => N3699, D => N4098, Q => 
                           REGISTERS_7_6_port);
   REGISTERS_reg_7_5_inst : DLH_X1 port map( G => N3699, D => N4096, Q => 
                           REGISTERS_7_5_port);
   REGISTERS_reg_7_4_inst : DLH_X1 port map( G => N3699, D => N4094, Q => 
                           REGISTERS_7_4_port);
   REGISTERS_reg_7_3_inst : DLH_X1 port map( G => N3699, D => N4092, Q => 
                           REGISTERS_7_3_port);
   REGISTERS_reg_7_2_inst : DLH_X1 port map( G => N3699, D => N4090, Q => 
                           REGISTERS_7_2_port);
   REGISTERS_reg_7_1_inst : DLH_X1 port map( G => N3699, D => N4088, Q => 
                           REGISTERS_7_1_port);
   REGISTERS_reg_7_0_inst : DLH_X1 port map( G => N3699, D => N4086, Q => 
                           REGISTERS_7_0_port);
   REGISTERS_reg_8_31_inst : DLH_X1 port map( G => N3635, D => N4148, Q => 
                           REGISTERS_8_31_port);
   REGISTERS_reg_8_30_inst : DLH_X1 port map( G => N3635, D => N4146, Q => 
                           REGISTERS_8_30_port);
   REGISTERS_reg_8_29_inst : DLH_X1 port map( G => N3635, D => N4144, Q => 
                           REGISTERS_8_29_port);
   REGISTERS_reg_8_28_inst : DLH_X1 port map( G => N3635, D => N4142, Q => 
                           REGISTERS_8_28_port);
   REGISTERS_reg_8_27_inst : DLH_X1 port map( G => N3635, D => N4140, Q => 
                           REGISTERS_8_27_port);
   REGISTERS_reg_8_26_inst : DLH_X1 port map( G => N3635, D => N4138, Q => 
                           REGISTERS_8_26_port);
   REGISTERS_reg_8_25_inst : DLH_X1 port map( G => N3635, D => N4136, Q => 
                           REGISTERS_8_25_port);
   REGISTERS_reg_8_24_inst : DLH_X1 port map( G => N3635, D => N4134, Q => 
                           REGISTERS_8_24_port);
   REGISTERS_reg_8_23_inst : DLH_X1 port map( G => N3635, D => N4132, Q => 
                           REGISTERS_8_23_port);
   REGISTERS_reg_8_22_inst : DLH_X1 port map( G => N3635, D => N4130, Q => 
                           REGISTERS_8_22_port);
   REGISTERS_reg_8_21_inst : DLH_X1 port map( G => N3635, D => N4128, Q => 
                           REGISTERS_8_21_port);
   REGISTERS_reg_8_20_inst : DLH_X1 port map( G => N3635, D => N4126, Q => 
                           REGISTERS_8_20_port);
   REGISTERS_reg_8_19_inst : DLH_X1 port map( G => N3635, D => N4124, Q => 
                           REGISTERS_8_19_port);
   REGISTERS_reg_8_18_inst : DLH_X1 port map( G => N3635, D => N4122, Q => 
                           REGISTERS_8_18_port);
   REGISTERS_reg_8_17_inst : DLH_X1 port map( G => N3635, D => N4120, Q => 
                           REGISTERS_8_17_port);
   REGISTERS_reg_8_16_inst : DLH_X1 port map( G => N3635, D => N4118, Q => 
                           REGISTERS_8_16_port);
   REGISTERS_reg_8_15_inst : DLH_X1 port map( G => N3635, D => N4116, Q => 
                           REGISTERS_8_15_port);
   REGISTERS_reg_8_14_inst : DLH_X1 port map( G => N3635, D => N4114, Q => 
                           REGISTERS_8_14_port);
   REGISTERS_reg_8_13_inst : DLH_X1 port map( G => N3635, D => N4112, Q => 
                           REGISTERS_8_13_port);
   REGISTERS_reg_8_12_inst : DLH_X1 port map( G => N3635, D => N4110, Q => 
                           REGISTERS_8_12_port);
   REGISTERS_reg_8_11_inst : DLH_X1 port map( G => N3635, D => N4108, Q => 
                           REGISTERS_8_11_port);
   REGISTERS_reg_8_10_inst : DLH_X1 port map( G => N3635, D => N4106, Q => 
                           REGISTERS_8_10_port);
   REGISTERS_reg_8_9_inst : DLH_X1 port map( G => N3635, D => N4104, Q => 
                           REGISTERS_8_9_port);
   REGISTERS_reg_8_8_inst : DLH_X1 port map( G => N3635, D => N4102, Q => 
                           REGISTERS_8_8_port);
   REGISTERS_reg_8_7_inst : DLH_X1 port map( G => N3635, D => N4100, Q => 
                           REGISTERS_8_7_port);
   REGISTERS_reg_8_6_inst : DLH_X1 port map( G => N3635, D => N4098, Q => 
                           REGISTERS_8_6_port);
   REGISTERS_reg_8_5_inst : DLH_X1 port map( G => N3635, D => N4096, Q => 
                           REGISTERS_8_5_port);
   REGISTERS_reg_8_4_inst : DLH_X1 port map( G => N3635, D => N4094, Q => 
                           REGISTERS_8_4_port);
   REGISTERS_reg_8_3_inst : DLH_X1 port map( G => N3635, D => N4092, Q => 
                           REGISTERS_8_3_port);
   REGISTERS_reg_8_2_inst : DLH_X1 port map( G => N3635, D => N4090, Q => 
                           REGISTERS_8_2_port);
   REGISTERS_reg_8_1_inst : DLH_X1 port map( G => N3635, D => N4088, Q => 
                           REGISTERS_8_1_port);
   REGISTERS_reg_8_0_inst : DLH_X1 port map( G => N3635, D => N4086, Q => 
                           REGISTERS_8_0_port);
   REGISTERS_reg_9_31_inst : DLH_X1 port map( G => N3571, D => N4148, Q => 
                           REGISTERS_9_31_port);
   REGISTERS_reg_9_30_inst : DLH_X1 port map( G => N3571, D => N4146, Q => 
                           REGISTERS_9_30_port);
   REGISTERS_reg_9_29_inst : DLH_X1 port map( G => N3571, D => N4144, Q => 
                           REGISTERS_9_29_port);
   REGISTERS_reg_9_28_inst : DLH_X1 port map( G => N3571, D => N4142, Q => 
                           REGISTERS_9_28_port);
   REGISTERS_reg_9_27_inst : DLH_X1 port map( G => N3571, D => N4140, Q => 
                           REGISTERS_9_27_port);
   REGISTERS_reg_9_26_inst : DLH_X1 port map( G => N3571, D => N4138, Q => 
                           REGISTERS_9_26_port);
   REGISTERS_reg_9_25_inst : DLH_X1 port map( G => N3571, D => N4136, Q => 
                           REGISTERS_9_25_port);
   REGISTERS_reg_9_24_inst : DLH_X1 port map( G => N3571, D => N4134, Q => 
                           REGISTERS_9_24_port);
   REGISTERS_reg_9_23_inst : DLH_X1 port map( G => N3571, D => N4132, Q => 
                           REGISTERS_9_23_port);
   REGISTERS_reg_9_22_inst : DLH_X1 port map( G => N3571, D => N4130, Q => 
                           REGISTERS_9_22_port);
   REGISTERS_reg_9_21_inst : DLH_X1 port map( G => N3571, D => N4128, Q => 
                           REGISTERS_9_21_port);
   REGISTERS_reg_9_20_inst : DLH_X1 port map( G => N3571, D => N4126, Q => 
                           REGISTERS_9_20_port);
   REGISTERS_reg_9_19_inst : DLH_X1 port map( G => N3571, D => N4124, Q => 
                           REGISTERS_9_19_port);
   REGISTERS_reg_9_18_inst : DLH_X1 port map( G => N3571, D => N4122, Q => 
                           REGISTERS_9_18_port);
   REGISTERS_reg_9_17_inst : DLH_X1 port map( G => N3571, D => N4120, Q => 
                           REGISTERS_9_17_port);
   REGISTERS_reg_9_16_inst : DLH_X1 port map( G => N3571, D => N4118, Q => 
                           REGISTERS_9_16_port);
   REGISTERS_reg_9_15_inst : DLH_X1 port map( G => N3571, D => N4116, Q => 
                           REGISTERS_9_15_port);
   REGISTERS_reg_9_14_inst : DLH_X1 port map( G => N3571, D => N4114, Q => 
                           REGISTERS_9_14_port);
   REGISTERS_reg_9_13_inst : DLH_X1 port map( G => N3571, D => N4112, Q => 
                           REGISTERS_9_13_port);
   REGISTERS_reg_9_12_inst : DLH_X1 port map( G => N3571, D => N4110, Q => 
                           REGISTERS_9_12_port);
   REGISTERS_reg_9_11_inst : DLH_X1 port map( G => N3571, D => N4108, Q => 
                           REGISTERS_9_11_port);
   REGISTERS_reg_9_10_inst : DLH_X1 port map( G => N3571, D => N4106, Q => 
                           REGISTERS_9_10_port);
   REGISTERS_reg_9_9_inst : DLH_X1 port map( G => N3571, D => N4104, Q => 
                           REGISTERS_9_9_port);
   REGISTERS_reg_9_8_inst : DLH_X1 port map( G => N3571, D => N4102, Q => 
                           REGISTERS_9_8_port);
   REGISTERS_reg_9_7_inst : DLH_X1 port map( G => N3571, D => N4100, Q => 
                           REGISTERS_9_7_port);
   REGISTERS_reg_9_6_inst : DLH_X1 port map( G => N3571, D => N4098, Q => 
                           REGISTERS_9_6_port);
   REGISTERS_reg_9_5_inst : DLH_X1 port map( G => N3571, D => N4096, Q => 
                           REGISTERS_9_5_port);
   REGISTERS_reg_9_4_inst : DLH_X1 port map( G => N3571, D => N4094, Q => 
                           REGISTERS_9_4_port);
   REGISTERS_reg_9_3_inst : DLH_X1 port map( G => N3571, D => N4092, Q => 
                           REGISTERS_9_3_port);
   REGISTERS_reg_9_2_inst : DLH_X1 port map( G => N3571, D => N4090, Q => 
                           REGISTERS_9_2_port);
   REGISTERS_reg_9_1_inst : DLH_X1 port map( G => N3571, D => N4088, Q => 
                           REGISTERS_9_1_port);
   REGISTERS_reg_9_0_inst : DLH_X1 port map( G => N3571, D => N4086, Q => 
                           REGISTERS_9_0_port);
   REGISTERS_reg_10_31_inst : DLH_X1 port map( G => N3507, D => N4148, Q => 
                           REGISTERS_10_31_port);
   REGISTERS_reg_10_30_inst : DLH_X1 port map( G => N3507, D => N4146, Q => 
                           REGISTERS_10_30_port);
   REGISTERS_reg_10_29_inst : DLH_X1 port map( G => N3507, D => N4144, Q => 
                           REGISTERS_10_29_port);
   REGISTERS_reg_10_28_inst : DLH_X1 port map( G => N3507, D => N4142, Q => 
                           REGISTERS_10_28_port);
   REGISTERS_reg_10_27_inst : DLH_X1 port map( G => N3507, D => N4140, Q => 
                           REGISTERS_10_27_port);
   REGISTERS_reg_10_26_inst : DLH_X1 port map( G => N3507, D => N4138, Q => 
                           REGISTERS_10_26_port);
   REGISTERS_reg_10_25_inst : DLH_X1 port map( G => N3507, D => N4136, Q => 
                           REGISTERS_10_25_port);
   REGISTERS_reg_10_24_inst : DLH_X1 port map( G => N3507, D => N4134, Q => 
                           REGISTERS_10_24_port);
   REGISTERS_reg_10_23_inst : DLH_X1 port map( G => N3507, D => N4132, Q => 
                           REGISTERS_10_23_port);
   REGISTERS_reg_10_22_inst : DLH_X1 port map( G => N3507, D => N4130, Q => 
                           REGISTERS_10_22_port);
   REGISTERS_reg_10_21_inst : DLH_X1 port map( G => N3507, D => N4128, Q => 
                           REGISTERS_10_21_port);
   REGISTERS_reg_10_20_inst : DLH_X1 port map( G => N3507, D => N4126, Q => 
                           REGISTERS_10_20_port);
   REGISTERS_reg_10_19_inst : DLH_X1 port map( G => N3507, D => N4124, Q => 
                           REGISTERS_10_19_port);
   REGISTERS_reg_10_18_inst : DLH_X1 port map( G => N3507, D => N4122, Q => 
                           REGISTERS_10_18_port);
   REGISTERS_reg_10_17_inst : DLH_X1 port map( G => N3507, D => N4120, Q => 
                           REGISTERS_10_17_port);
   REGISTERS_reg_10_16_inst : DLH_X1 port map( G => N3507, D => N4118, Q => 
                           REGISTERS_10_16_port);
   REGISTERS_reg_10_15_inst : DLH_X1 port map( G => N3507, D => N4116, Q => 
                           REGISTERS_10_15_port);
   REGISTERS_reg_10_14_inst : DLH_X1 port map( G => N3507, D => N4114, Q => 
                           REGISTERS_10_14_port);
   REGISTERS_reg_10_13_inst : DLH_X1 port map( G => N3507, D => N4112, Q => 
                           REGISTERS_10_13_port);
   REGISTERS_reg_10_12_inst : DLH_X1 port map( G => N3507, D => N4110, Q => 
                           REGISTERS_10_12_port);
   REGISTERS_reg_10_11_inst : DLH_X1 port map( G => N3507, D => N4108, Q => 
                           REGISTERS_10_11_port);
   REGISTERS_reg_10_10_inst : DLH_X1 port map( G => N3507, D => N4106, Q => 
                           REGISTERS_10_10_port);
   REGISTERS_reg_10_9_inst : DLH_X1 port map( G => N3507, D => N4104, Q => 
                           REGISTERS_10_9_port);
   REGISTERS_reg_10_8_inst : DLH_X1 port map( G => N3507, D => N4102, Q => 
                           REGISTERS_10_8_port);
   REGISTERS_reg_10_7_inst : DLH_X1 port map( G => N3507, D => N4100, Q => 
                           REGISTERS_10_7_port);
   REGISTERS_reg_10_6_inst : DLH_X1 port map( G => N3507, D => N4098, Q => 
                           REGISTERS_10_6_port);
   REGISTERS_reg_10_5_inst : DLH_X1 port map( G => N3507, D => N4096, Q => 
                           REGISTERS_10_5_port);
   REGISTERS_reg_10_4_inst : DLH_X1 port map( G => N3507, D => N4094, Q => 
                           REGISTERS_10_4_port);
   REGISTERS_reg_10_3_inst : DLH_X1 port map( G => N3507, D => N4092, Q => 
                           REGISTERS_10_3_port);
   REGISTERS_reg_10_2_inst : DLH_X1 port map( G => N3507, D => N4090, Q => 
                           REGISTERS_10_2_port);
   REGISTERS_reg_10_1_inst : DLH_X1 port map( G => N3507, D => N4088, Q => 
                           REGISTERS_10_1_port);
   REGISTERS_reg_10_0_inst : DLH_X1 port map( G => N3507, D => N4086, Q => 
                           REGISTERS_10_0_port);
   REGISTERS_reg_11_31_inst : DLH_X1 port map( G => N3443, D => N4148, Q => 
                           REGISTERS_11_31_port);
   REGISTERS_reg_11_30_inst : DLH_X1 port map( G => N3443, D => N4146, Q => 
                           REGISTERS_11_30_port);
   REGISTERS_reg_11_29_inst : DLH_X1 port map( G => N3443, D => N4144, Q => 
                           REGISTERS_11_29_port);
   REGISTERS_reg_11_28_inst : DLH_X1 port map( G => N3443, D => N4142, Q => 
                           REGISTERS_11_28_port);
   REGISTERS_reg_11_27_inst : DLH_X1 port map( G => N3443, D => N4140, Q => 
                           REGISTERS_11_27_port);
   REGISTERS_reg_11_26_inst : DLH_X1 port map( G => N3443, D => N4138, Q => 
                           REGISTERS_11_26_port);
   REGISTERS_reg_11_25_inst : DLH_X1 port map( G => N3443, D => N4136, Q => 
                           REGISTERS_11_25_port);
   REGISTERS_reg_11_24_inst : DLH_X1 port map( G => N3443, D => N4134, Q => 
                           REGISTERS_11_24_port);
   REGISTERS_reg_11_23_inst : DLH_X1 port map( G => N3443, D => N4132, Q => 
                           REGISTERS_11_23_port);
   REGISTERS_reg_11_22_inst : DLH_X1 port map( G => N3443, D => N4130, Q => 
                           REGISTERS_11_22_port);
   REGISTERS_reg_11_21_inst : DLH_X1 port map( G => N3443, D => N4128, Q => 
                           REGISTERS_11_21_port);
   REGISTERS_reg_11_20_inst : DLH_X1 port map( G => N3443, D => N4126, Q => 
                           REGISTERS_11_20_port);
   REGISTERS_reg_11_19_inst : DLH_X1 port map( G => N3443, D => N4124, Q => 
                           REGISTERS_11_19_port);
   REGISTERS_reg_11_18_inst : DLH_X1 port map( G => N3443, D => N4122, Q => 
                           REGISTERS_11_18_port);
   REGISTERS_reg_11_17_inst : DLH_X1 port map( G => N3443, D => N4120, Q => 
                           REGISTERS_11_17_port);
   REGISTERS_reg_11_16_inst : DLH_X1 port map( G => N3443, D => N4118, Q => 
                           REGISTERS_11_16_port);
   REGISTERS_reg_11_15_inst : DLH_X1 port map( G => N3443, D => N4116, Q => 
                           REGISTERS_11_15_port);
   REGISTERS_reg_11_14_inst : DLH_X1 port map( G => N3443, D => N4114, Q => 
                           REGISTERS_11_14_port);
   REGISTERS_reg_11_13_inst : DLH_X1 port map( G => N3443, D => N4112, Q => 
                           REGISTERS_11_13_port);
   REGISTERS_reg_11_12_inst : DLH_X1 port map( G => N3443, D => N4110, Q => 
                           REGISTERS_11_12_port);
   REGISTERS_reg_11_11_inst : DLH_X1 port map( G => N3443, D => N4108, Q => 
                           REGISTERS_11_11_port);
   REGISTERS_reg_11_10_inst : DLH_X1 port map( G => N3443, D => N4106, Q => 
                           REGISTERS_11_10_port);
   REGISTERS_reg_11_9_inst : DLH_X1 port map( G => N3443, D => N4104, Q => 
                           REGISTERS_11_9_port);
   REGISTERS_reg_11_8_inst : DLH_X1 port map( G => N3443, D => N4102, Q => 
                           REGISTERS_11_8_port);
   REGISTERS_reg_11_7_inst : DLH_X1 port map( G => N3443, D => N4100, Q => 
                           REGISTERS_11_7_port);
   REGISTERS_reg_11_6_inst : DLH_X1 port map( G => N3443, D => N4098, Q => 
                           REGISTERS_11_6_port);
   REGISTERS_reg_11_5_inst : DLH_X1 port map( G => N3443, D => N4096, Q => 
                           REGISTERS_11_5_port);
   REGISTERS_reg_11_4_inst : DLH_X1 port map( G => N3443, D => N4094, Q => 
                           REGISTERS_11_4_port);
   REGISTERS_reg_11_3_inst : DLH_X1 port map( G => N3443, D => N4092, Q => 
                           REGISTERS_11_3_port);
   REGISTERS_reg_11_2_inst : DLH_X1 port map( G => N3443, D => N4090, Q => 
                           REGISTERS_11_2_port);
   REGISTERS_reg_11_1_inst : DLH_X1 port map( G => N3443, D => N4088, Q => 
                           REGISTERS_11_1_port);
   REGISTERS_reg_11_0_inst : DLH_X1 port map( G => N3443, D => N4086, Q => 
                           REGISTERS_11_0_port);
   REGISTERS_reg_12_31_inst : DLH_X1 port map( G => N3379, D => N4148, Q => 
                           REGISTERS_12_31_port);
   REGISTERS_reg_12_30_inst : DLH_X1 port map( G => N3379, D => N4146, Q => 
                           REGISTERS_12_30_port);
   REGISTERS_reg_12_29_inst : DLH_X1 port map( G => N3379, D => N4144, Q => 
                           REGISTERS_12_29_port);
   REGISTERS_reg_12_28_inst : DLH_X1 port map( G => N3379, D => N4142, Q => 
                           REGISTERS_12_28_port);
   REGISTERS_reg_12_27_inst : DLH_X1 port map( G => N3379, D => N4140, Q => 
                           REGISTERS_12_27_port);
   REGISTERS_reg_12_26_inst : DLH_X1 port map( G => N3379, D => N4138, Q => 
                           REGISTERS_12_26_port);
   REGISTERS_reg_12_25_inst : DLH_X1 port map( G => N3379, D => N4136, Q => 
                           REGISTERS_12_25_port);
   REGISTERS_reg_12_24_inst : DLH_X1 port map( G => N3379, D => N4134, Q => 
                           REGISTERS_12_24_port);
   REGISTERS_reg_12_23_inst : DLH_X1 port map( G => N3379, D => N4132, Q => 
                           REGISTERS_12_23_port);
   REGISTERS_reg_12_22_inst : DLH_X1 port map( G => N3379, D => N4130, Q => 
                           REGISTERS_12_22_port);
   REGISTERS_reg_12_21_inst : DLH_X1 port map( G => N3379, D => N4128, Q => 
                           REGISTERS_12_21_port);
   REGISTERS_reg_12_20_inst : DLH_X1 port map( G => N3379, D => N4126, Q => 
                           REGISTERS_12_20_port);
   REGISTERS_reg_12_19_inst : DLH_X1 port map( G => N3379, D => N4124, Q => 
                           REGISTERS_12_19_port);
   REGISTERS_reg_12_18_inst : DLH_X1 port map( G => N3379, D => N4122, Q => 
                           REGISTERS_12_18_port);
   REGISTERS_reg_12_17_inst : DLH_X1 port map( G => N3379, D => N4120, Q => 
                           REGISTERS_12_17_port);
   REGISTERS_reg_12_16_inst : DLH_X1 port map( G => N3379, D => N4118, Q => 
                           REGISTERS_12_16_port);
   REGISTERS_reg_12_15_inst : DLH_X1 port map( G => N3379, D => N4116, Q => 
                           REGISTERS_12_15_port);
   REGISTERS_reg_12_14_inst : DLH_X1 port map( G => N3379, D => N4114, Q => 
                           REGISTERS_12_14_port);
   REGISTERS_reg_12_13_inst : DLH_X1 port map( G => N3379, D => N4112, Q => 
                           REGISTERS_12_13_port);
   REGISTERS_reg_12_12_inst : DLH_X1 port map( G => N3379, D => N4110, Q => 
                           REGISTERS_12_12_port);
   REGISTERS_reg_12_11_inst : DLH_X1 port map( G => N3379, D => N4108, Q => 
                           REGISTERS_12_11_port);
   REGISTERS_reg_12_10_inst : DLH_X1 port map( G => N3379, D => N4106, Q => 
                           REGISTERS_12_10_port);
   REGISTERS_reg_12_9_inst : DLH_X1 port map( G => N3379, D => N4104, Q => 
                           REGISTERS_12_9_port);
   REGISTERS_reg_12_8_inst : DLH_X1 port map( G => N3379, D => N4102, Q => 
                           REGISTERS_12_8_port);
   REGISTERS_reg_12_7_inst : DLH_X1 port map( G => N3379, D => N4100, Q => 
                           REGISTERS_12_7_port);
   REGISTERS_reg_12_6_inst : DLH_X1 port map( G => N3379, D => N4098, Q => 
                           REGISTERS_12_6_port);
   REGISTERS_reg_12_5_inst : DLH_X1 port map( G => N3379, D => N4096, Q => 
                           REGISTERS_12_5_port);
   REGISTERS_reg_12_4_inst : DLH_X1 port map( G => N3379, D => N4094, Q => 
                           REGISTERS_12_4_port);
   REGISTERS_reg_12_3_inst : DLH_X1 port map( G => N3379, D => N4092, Q => 
                           REGISTERS_12_3_port);
   REGISTERS_reg_12_2_inst : DLH_X1 port map( G => N3379, D => N4090, Q => 
                           REGISTERS_12_2_port);
   REGISTERS_reg_12_1_inst : DLH_X1 port map( G => N3379, D => N4088, Q => 
                           REGISTERS_12_1_port);
   REGISTERS_reg_12_0_inst : DLH_X1 port map( G => N3379, D => N4086, Q => 
                           REGISTERS_12_0_port);
   REGISTERS_reg_13_31_inst : DLH_X1 port map( G => N3315, D => N4148, Q => 
                           REGISTERS_13_31_port);
   REGISTERS_reg_13_30_inst : DLH_X1 port map( G => N3315, D => N4146, Q => 
                           REGISTERS_13_30_port);
   REGISTERS_reg_13_29_inst : DLH_X1 port map( G => N3315, D => N4144, Q => 
                           REGISTERS_13_29_port);
   REGISTERS_reg_13_28_inst : DLH_X1 port map( G => N3315, D => N4142, Q => 
                           REGISTERS_13_28_port);
   REGISTERS_reg_13_27_inst : DLH_X1 port map( G => N3315, D => N4140, Q => 
                           REGISTERS_13_27_port);
   REGISTERS_reg_13_26_inst : DLH_X1 port map( G => N3315, D => N4138, Q => 
                           REGISTERS_13_26_port);
   REGISTERS_reg_13_25_inst : DLH_X1 port map( G => N3315, D => N4136, Q => 
                           REGISTERS_13_25_port);
   REGISTERS_reg_13_24_inst : DLH_X1 port map( G => N3315, D => N4134, Q => 
                           REGISTERS_13_24_port);
   REGISTERS_reg_13_23_inst : DLH_X1 port map( G => N3315, D => N4132, Q => 
                           REGISTERS_13_23_port);
   REGISTERS_reg_13_22_inst : DLH_X1 port map( G => N3315, D => N4130, Q => 
                           REGISTERS_13_22_port);
   REGISTERS_reg_13_21_inst : DLH_X1 port map( G => N3315, D => N4128, Q => 
                           REGISTERS_13_21_port);
   REGISTERS_reg_13_20_inst : DLH_X1 port map( G => N3315, D => N4126, Q => 
                           REGISTERS_13_20_port);
   REGISTERS_reg_13_19_inst : DLH_X1 port map( G => N3315, D => N4124, Q => 
                           REGISTERS_13_19_port);
   REGISTERS_reg_13_18_inst : DLH_X1 port map( G => N3315, D => N4122, Q => 
                           REGISTERS_13_18_port);
   REGISTERS_reg_13_17_inst : DLH_X1 port map( G => N3315, D => N4120, Q => 
                           REGISTERS_13_17_port);
   REGISTERS_reg_13_16_inst : DLH_X1 port map( G => N3315, D => N4118, Q => 
                           REGISTERS_13_16_port);
   REGISTERS_reg_13_15_inst : DLH_X1 port map( G => N3315, D => N4116, Q => 
                           REGISTERS_13_15_port);
   REGISTERS_reg_13_14_inst : DLH_X1 port map( G => N3315, D => N4114, Q => 
                           REGISTERS_13_14_port);
   REGISTERS_reg_13_13_inst : DLH_X1 port map( G => N3315, D => N4112, Q => 
                           REGISTERS_13_13_port);
   REGISTERS_reg_13_12_inst : DLH_X1 port map( G => N3315, D => N4110, Q => 
                           REGISTERS_13_12_port);
   REGISTERS_reg_13_11_inst : DLH_X1 port map( G => N3315, D => N4108, Q => 
                           REGISTERS_13_11_port);
   REGISTERS_reg_13_10_inst : DLH_X1 port map( G => N3315, D => N4106, Q => 
                           REGISTERS_13_10_port);
   REGISTERS_reg_13_9_inst : DLH_X1 port map( G => N3315, D => N4104, Q => 
                           REGISTERS_13_9_port);
   REGISTERS_reg_13_8_inst : DLH_X1 port map( G => N3315, D => N4102, Q => 
                           REGISTERS_13_8_port);
   REGISTERS_reg_13_7_inst : DLH_X1 port map( G => N3315, D => N4100, Q => 
                           REGISTERS_13_7_port);
   REGISTERS_reg_13_6_inst : DLH_X1 port map( G => N3315, D => N4098, Q => 
                           REGISTERS_13_6_port);
   REGISTERS_reg_13_5_inst : DLH_X1 port map( G => N3315, D => N4096, Q => 
                           REGISTERS_13_5_port);
   REGISTERS_reg_13_4_inst : DLH_X1 port map( G => N3315, D => N4094, Q => 
                           REGISTERS_13_4_port);
   REGISTERS_reg_13_3_inst : DLH_X1 port map( G => N3315, D => N4092, Q => 
                           REGISTERS_13_3_port);
   REGISTERS_reg_13_2_inst : DLH_X1 port map( G => N3315, D => N4090, Q => 
                           REGISTERS_13_2_port);
   REGISTERS_reg_13_1_inst : DLH_X1 port map( G => N3315, D => N4088, Q => 
                           REGISTERS_13_1_port);
   REGISTERS_reg_13_0_inst : DLH_X1 port map( G => N3315, D => N4086, Q => 
                           REGISTERS_13_0_port);
   REGISTERS_reg_14_31_inst : DLH_X1 port map( G => N3251, D => N4148, Q => 
                           REGISTERS_14_31_port);
   REGISTERS_reg_14_30_inst : DLH_X1 port map( G => N3251, D => N4146, Q => 
                           REGISTERS_14_30_port);
   REGISTERS_reg_14_29_inst : DLH_X1 port map( G => N3251, D => N4144, Q => 
                           REGISTERS_14_29_port);
   REGISTERS_reg_14_28_inst : DLH_X1 port map( G => N3251, D => N4142, Q => 
                           REGISTERS_14_28_port);
   REGISTERS_reg_14_27_inst : DLH_X1 port map( G => N3251, D => N4140, Q => 
                           REGISTERS_14_27_port);
   REGISTERS_reg_14_26_inst : DLH_X1 port map( G => N3251, D => N4138, Q => 
                           REGISTERS_14_26_port);
   REGISTERS_reg_14_25_inst : DLH_X1 port map( G => N3251, D => N4136, Q => 
                           REGISTERS_14_25_port);
   REGISTERS_reg_14_24_inst : DLH_X1 port map( G => N3251, D => N4134, Q => 
                           REGISTERS_14_24_port);
   REGISTERS_reg_14_23_inst : DLH_X1 port map( G => N3251, D => N4132, Q => 
                           REGISTERS_14_23_port);
   REGISTERS_reg_14_22_inst : DLH_X1 port map( G => N3251, D => N4130, Q => 
                           REGISTERS_14_22_port);
   REGISTERS_reg_14_21_inst : DLH_X1 port map( G => N3251, D => N4128, Q => 
                           REGISTERS_14_21_port);
   REGISTERS_reg_14_20_inst : DLH_X1 port map( G => N3251, D => N4126, Q => 
                           REGISTERS_14_20_port);
   REGISTERS_reg_14_19_inst : DLH_X1 port map( G => N3251, D => N4124, Q => 
                           REGISTERS_14_19_port);
   REGISTERS_reg_14_18_inst : DLH_X1 port map( G => N3251, D => N4122, Q => 
                           REGISTERS_14_18_port);
   REGISTERS_reg_14_17_inst : DLH_X1 port map( G => N3251, D => N4120, Q => 
                           REGISTERS_14_17_port);
   REGISTERS_reg_14_16_inst : DLH_X1 port map( G => N3251, D => N4118, Q => 
                           REGISTERS_14_16_port);
   REGISTERS_reg_14_15_inst : DLH_X1 port map( G => N3251, D => N4116, Q => 
                           REGISTERS_14_15_port);
   REGISTERS_reg_14_14_inst : DLH_X1 port map( G => N3251, D => N4114, Q => 
                           REGISTERS_14_14_port);
   REGISTERS_reg_14_13_inst : DLH_X1 port map( G => N3251, D => N4112, Q => 
                           REGISTERS_14_13_port);
   REGISTERS_reg_14_12_inst : DLH_X1 port map( G => N3251, D => N4110, Q => 
                           REGISTERS_14_12_port);
   REGISTERS_reg_14_11_inst : DLH_X1 port map( G => N3251, D => N4108, Q => 
                           REGISTERS_14_11_port);
   REGISTERS_reg_14_10_inst : DLH_X1 port map( G => N3251, D => N4106, Q => 
                           REGISTERS_14_10_port);
   REGISTERS_reg_14_9_inst : DLH_X1 port map( G => N3251, D => N4104, Q => 
                           REGISTERS_14_9_port);
   REGISTERS_reg_14_8_inst : DLH_X1 port map( G => N3251, D => N4102, Q => 
                           REGISTERS_14_8_port);
   REGISTERS_reg_14_7_inst : DLH_X1 port map( G => N3251, D => N4100, Q => 
                           REGISTERS_14_7_port);
   REGISTERS_reg_14_6_inst : DLH_X1 port map( G => N3251, D => N4098, Q => 
                           REGISTERS_14_6_port);
   REGISTERS_reg_14_5_inst : DLH_X1 port map( G => N3251, D => N4096, Q => 
                           REGISTERS_14_5_port);
   REGISTERS_reg_14_4_inst : DLH_X1 port map( G => N3251, D => N4094, Q => 
                           REGISTERS_14_4_port);
   REGISTERS_reg_14_3_inst : DLH_X1 port map( G => N3251, D => N4092, Q => 
                           REGISTERS_14_3_port);
   REGISTERS_reg_14_2_inst : DLH_X1 port map( G => N3251, D => N4090, Q => 
                           REGISTERS_14_2_port);
   REGISTERS_reg_14_1_inst : DLH_X1 port map( G => N3251, D => N4088, Q => 
                           REGISTERS_14_1_port);
   REGISTERS_reg_14_0_inst : DLH_X1 port map( G => N3251, D => N4086, Q => 
                           REGISTERS_14_0_port);
   REGISTERS_reg_15_31_inst : DLH_X1 port map( G => N3187, D => N4148, Q => 
                           REGISTERS_15_31_port);
   REGISTERS_reg_15_30_inst : DLH_X1 port map( G => N3187, D => N4146, Q => 
                           REGISTERS_15_30_port);
   REGISTERS_reg_15_29_inst : DLH_X1 port map( G => N3187, D => N4144, Q => 
                           REGISTERS_15_29_port);
   REGISTERS_reg_15_28_inst : DLH_X1 port map( G => N3187, D => N4142, Q => 
                           REGISTERS_15_28_port);
   REGISTERS_reg_15_27_inst : DLH_X1 port map( G => N3187, D => N4140, Q => 
                           REGISTERS_15_27_port);
   REGISTERS_reg_15_26_inst : DLH_X1 port map( G => N3187, D => N4138, Q => 
                           REGISTERS_15_26_port);
   REGISTERS_reg_15_25_inst : DLH_X1 port map( G => N3187, D => N4136, Q => 
                           REGISTERS_15_25_port);
   REGISTERS_reg_15_24_inst : DLH_X1 port map( G => N3187, D => N4134, Q => 
                           REGISTERS_15_24_port);
   REGISTERS_reg_15_23_inst : DLH_X1 port map( G => N3187, D => N4132, Q => 
                           REGISTERS_15_23_port);
   REGISTERS_reg_15_22_inst : DLH_X1 port map( G => N3187, D => N4130, Q => 
                           REGISTERS_15_22_port);
   REGISTERS_reg_15_21_inst : DLH_X1 port map( G => N3187, D => N4128, Q => 
                           REGISTERS_15_21_port);
   REGISTERS_reg_15_20_inst : DLH_X1 port map( G => N3187, D => N4126, Q => 
                           REGISTERS_15_20_port);
   REGISTERS_reg_15_19_inst : DLH_X1 port map( G => N3187, D => N4124, Q => 
                           REGISTERS_15_19_port);
   REGISTERS_reg_15_18_inst : DLH_X1 port map( G => N3187, D => N4122, Q => 
                           REGISTERS_15_18_port);
   REGISTERS_reg_15_17_inst : DLH_X1 port map( G => N3187, D => N4120, Q => 
                           REGISTERS_15_17_port);
   REGISTERS_reg_15_16_inst : DLH_X1 port map( G => N3187, D => N4118, Q => 
                           REGISTERS_15_16_port);
   REGISTERS_reg_15_15_inst : DLH_X1 port map( G => N3187, D => N4116, Q => 
                           REGISTERS_15_15_port);
   REGISTERS_reg_15_14_inst : DLH_X1 port map( G => N3187, D => N4114, Q => 
                           REGISTERS_15_14_port);
   REGISTERS_reg_15_13_inst : DLH_X1 port map( G => N3187, D => N4112, Q => 
                           REGISTERS_15_13_port);
   REGISTERS_reg_15_12_inst : DLH_X1 port map( G => N3187, D => N4110, Q => 
                           REGISTERS_15_12_port);
   REGISTERS_reg_15_11_inst : DLH_X1 port map( G => N3187, D => N4108, Q => 
                           REGISTERS_15_11_port);
   REGISTERS_reg_15_10_inst : DLH_X1 port map( G => N3187, D => N4106, Q => 
                           REGISTERS_15_10_port);
   REGISTERS_reg_15_9_inst : DLH_X1 port map( G => N3187, D => N4104, Q => 
                           REGISTERS_15_9_port);
   REGISTERS_reg_15_8_inst : DLH_X1 port map( G => N3187, D => N4102, Q => 
                           REGISTERS_15_8_port);
   REGISTERS_reg_15_7_inst : DLH_X1 port map( G => N3187, D => N4100, Q => 
                           REGISTERS_15_7_port);
   REGISTERS_reg_15_6_inst : DLH_X1 port map( G => N3187, D => N4098, Q => 
                           REGISTERS_15_6_port);
   REGISTERS_reg_15_5_inst : DLH_X1 port map( G => N3187, D => N4096, Q => 
                           REGISTERS_15_5_port);
   REGISTERS_reg_15_4_inst : DLH_X1 port map( G => N3187, D => N4094, Q => 
                           REGISTERS_15_4_port);
   REGISTERS_reg_15_3_inst : DLH_X1 port map( G => N3187, D => N4092, Q => 
                           REGISTERS_15_3_port);
   REGISTERS_reg_15_2_inst : DLH_X1 port map( G => N3187, D => N4090, Q => 
                           REGISTERS_15_2_port);
   REGISTERS_reg_15_1_inst : DLH_X1 port map( G => N3187, D => N4088, Q => 
                           REGISTERS_15_1_port);
   REGISTERS_reg_15_0_inst : DLH_X1 port map( G => N3187, D => N4086, Q => 
                           REGISTERS_15_0_port);
   REGISTERS_reg_16_31_inst : DLH_X1 port map( G => N3123, D => N4148, Q => 
                           REGISTERS_16_31_port);
   REGISTERS_reg_16_30_inst : DLH_X1 port map( G => N3123, D => N4146, Q => 
                           REGISTERS_16_30_port);
   REGISTERS_reg_16_29_inst : DLH_X1 port map( G => N3123, D => N4144, Q => 
                           REGISTERS_16_29_port);
   REGISTERS_reg_16_28_inst : DLH_X1 port map( G => N3123, D => N4142, Q => 
                           REGISTERS_16_28_port);
   REGISTERS_reg_16_27_inst : DLH_X1 port map( G => N3123, D => N4140, Q => 
                           REGISTERS_16_27_port);
   REGISTERS_reg_16_26_inst : DLH_X1 port map( G => N3123, D => N4138, Q => 
                           REGISTERS_16_26_port);
   REGISTERS_reg_16_25_inst : DLH_X1 port map( G => N3123, D => N4136, Q => 
                           REGISTERS_16_25_port);
   REGISTERS_reg_16_24_inst : DLH_X1 port map( G => N3123, D => N4134, Q => 
                           REGISTERS_16_24_port);
   REGISTERS_reg_16_23_inst : DLH_X1 port map( G => N3123, D => N4132, Q => 
                           REGISTERS_16_23_port);
   REGISTERS_reg_16_22_inst : DLH_X1 port map( G => N3123, D => N4130, Q => 
                           REGISTERS_16_22_port);
   REGISTERS_reg_16_21_inst : DLH_X1 port map( G => N3123, D => N4128, Q => 
                           REGISTERS_16_21_port);
   REGISTERS_reg_16_20_inst : DLH_X1 port map( G => N3123, D => N4126, Q => 
                           REGISTERS_16_20_port);
   REGISTERS_reg_16_19_inst : DLH_X1 port map( G => N3123, D => N4124, Q => 
                           REGISTERS_16_19_port);
   REGISTERS_reg_16_18_inst : DLH_X1 port map( G => N3123, D => N4122, Q => 
                           REGISTERS_16_18_port);
   REGISTERS_reg_16_17_inst : DLH_X1 port map( G => N3123, D => N4120, Q => 
                           REGISTERS_16_17_port);
   REGISTERS_reg_16_16_inst : DLH_X1 port map( G => N3123, D => N4118, Q => 
                           REGISTERS_16_16_port);
   REGISTERS_reg_16_15_inst : DLH_X1 port map( G => N3123, D => N4116, Q => 
                           REGISTERS_16_15_port);
   REGISTERS_reg_16_14_inst : DLH_X1 port map( G => N3123, D => N4114, Q => 
                           REGISTERS_16_14_port);
   REGISTERS_reg_16_13_inst : DLH_X1 port map( G => N3123, D => N4112, Q => 
                           REGISTERS_16_13_port);
   REGISTERS_reg_16_12_inst : DLH_X1 port map( G => N3123, D => N4110, Q => 
                           REGISTERS_16_12_port);
   REGISTERS_reg_16_11_inst : DLH_X1 port map( G => N3123, D => N4108, Q => 
                           REGISTERS_16_11_port);
   REGISTERS_reg_16_10_inst : DLH_X1 port map( G => N3123, D => N4106, Q => 
                           REGISTERS_16_10_port);
   REGISTERS_reg_16_9_inst : DLH_X1 port map( G => N3123, D => N4104, Q => 
                           REGISTERS_16_9_port);
   REGISTERS_reg_16_8_inst : DLH_X1 port map( G => N3123, D => N4102, Q => 
                           REGISTERS_16_8_port);
   REGISTERS_reg_16_7_inst : DLH_X1 port map( G => N3123, D => N4100, Q => 
                           REGISTERS_16_7_port);
   REGISTERS_reg_16_6_inst : DLH_X1 port map( G => N3123, D => N4098, Q => 
                           REGISTERS_16_6_port);
   REGISTERS_reg_16_5_inst : DLH_X1 port map( G => N3123, D => N4096, Q => 
                           REGISTERS_16_5_port);
   REGISTERS_reg_16_4_inst : DLH_X1 port map( G => N3123, D => N4094, Q => 
                           REGISTERS_16_4_port);
   REGISTERS_reg_16_3_inst : DLH_X1 port map( G => N3123, D => N4092, Q => 
                           REGISTERS_16_3_port);
   REGISTERS_reg_16_2_inst : DLH_X1 port map( G => N3123, D => N4090, Q => 
                           REGISTERS_16_2_port);
   REGISTERS_reg_16_1_inst : DLH_X1 port map( G => N3123, D => N4088, Q => 
                           REGISTERS_16_1_port);
   REGISTERS_reg_16_0_inst : DLH_X1 port map( G => N3123, D => N4086, Q => 
                           REGISTERS_16_0_port);
   REGISTERS_reg_17_31_inst : DLH_X1 port map( G => N3059, D => N4148, Q => 
                           REGISTERS_17_31_port);
   REGISTERS_reg_17_30_inst : DLH_X1 port map( G => N3059, D => N4146, Q => 
                           REGISTERS_17_30_port);
   REGISTERS_reg_17_29_inst : DLH_X1 port map( G => N3059, D => N4144, Q => 
                           REGISTERS_17_29_port);
   REGISTERS_reg_17_28_inst : DLH_X1 port map( G => N3059, D => N4142, Q => 
                           REGISTERS_17_28_port);
   REGISTERS_reg_17_27_inst : DLH_X1 port map( G => N3059, D => N4140, Q => 
                           REGISTERS_17_27_port);
   REGISTERS_reg_17_26_inst : DLH_X1 port map( G => N3059, D => N4138, Q => 
                           REGISTERS_17_26_port);
   REGISTERS_reg_17_25_inst : DLH_X1 port map( G => N3059, D => N4136, Q => 
                           REGISTERS_17_25_port);
   REGISTERS_reg_17_24_inst : DLH_X1 port map( G => N3059, D => N4134, Q => 
                           REGISTERS_17_24_port);
   REGISTERS_reg_17_23_inst : DLH_X1 port map( G => N3059, D => N4132, Q => 
                           REGISTERS_17_23_port);
   REGISTERS_reg_17_22_inst : DLH_X1 port map( G => N3059, D => N4130, Q => 
                           REGISTERS_17_22_port);
   REGISTERS_reg_17_21_inst : DLH_X1 port map( G => N3059, D => N4128, Q => 
                           REGISTERS_17_21_port);
   REGISTERS_reg_17_20_inst : DLH_X1 port map( G => N3059, D => N4126, Q => 
                           REGISTERS_17_20_port);
   REGISTERS_reg_17_19_inst : DLH_X1 port map( G => N3059, D => N4124, Q => 
                           REGISTERS_17_19_port);
   REGISTERS_reg_17_18_inst : DLH_X1 port map( G => N3059, D => N4122, Q => 
                           REGISTERS_17_18_port);
   REGISTERS_reg_17_17_inst : DLH_X1 port map( G => N3059, D => N4120, Q => 
                           REGISTERS_17_17_port);
   REGISTERS_reg_17_16_inst : DLH_X1 port map( G => N3059, D => N4118, Q => 
                           REGISTERS_17_16_port);
   REGISTERS_reg_17_15_inst : DLH_X1 port map( G => N3059, D => N4116, Q => 
                           REGISTERS_17_15_port);
   REGISTERS_reg_17_14_inst : DLH_X1 port map( G => N3059, D => N4114, Q => 
                           REGISTERS_17_14_port);
   REGISTERS_reg_17_13_inst : DLH_X1 port map( G => N3059, D => N4112, Q => 
                           REGISTERS_17_13_port);
   REGISTERS_reg_17_12_inst : DLH_X1 port map( G => N3059, D => N4110, Q => 
                           REGISTERS_17_12_port);
   REGISTERS_reg_17_11_inst : DLH_X1 port map( G => N3059, D => N4108, Q => 
                           REGISTERS_17_11_port);
   REGISTERS_reg_17_10_inst : DLH_X1 port map( G => N3059, D => N4106, Q => 
                           REGISTERS_17_10_port);
   REGISTERS_reg_17_9_inst : DLH_X1 port map( G => N3059, D => N4104, Q => 
                           REGISTERS_17_9_port);
   REGISTERS_reg_17_8_inst : DLH_X1 port map( G => N3059, D => N4102, Q => 
                           REGISTERS_17_8_port);
   REGISTERS_reg_17_7_inst : DLH_X1 port map( G => N3059, D => N4100, Q => 
                           REGISTERS_17_7_port);
   REGISTERS_reg_17_6_inst : DLH_X1 port map( G => N3059, D => N4098, Q => 
                           REGISTERS_17_6_port);
   REGISTERS_reg_17_5_inst : DLH_X1 port map( G => N3059, D => N4096, Q => 
                           REGISTERS_17_5_port);
   REGISTERS_reg_17_4_inst : DLH_X1 port map( G => N3059, D => N4094, Q => 
                           REGISTERS_17_4_port);
   REGISTERS_reg_17_3_inst : DLH_X1 port map( G => N3059, D => N4092, Q => 
                           REGISTERS_17_3_port);
   REGISTERS_reg_17_2_inst : DLH_X1 port map( G => N3059, D => N4090, Q => 
                           REGISTERS_17_2_port);
   REGISTERS_reg_17_1_inst : DLH_X1 port map( G => N3059, D => N4088, Q => 
                           REGISTERS_17_1_port);
   REGISTERS_reg_17_0_inst : DLH_X1 port map( G => N3059, D => N4086, Q => 
                           REGISTERS_17_0_port);
   REGISTERS_reg_18_31_inst : DLH_X1 port map( G => N2995, D => N4148, Q => 
                           REGISTERS_18_31_port);
   REGISTERS_reg_18_30_inst : DLH_X1 port map( G => N2995, D => N4146, Q => 
                           REGISTERS_18_30_port);
   REGISTERS_reg_18_29_inst : DLH_X1 port map( G => N2995, D => N4144, Q => 
                           REGISTERS_18_29_port);
   REGISTERS_reg_18_28_inst : DLH_X1 port map( G => N2995, D => N4142, Q => 
                           REGISTERS_18_28_port);
   REGISTERS_reg_18_27_inst : DLH_X1 port map( G => N2995, D => N4140, Q => 
                           REGISTERS_18_27_port);
   REGISTERS_reg_18_26_inst : DLH_X1 port map( G => N2995, D => N4138, Q => 
                           REGISTERS_18_26_port);
   REGISTERS_reg_18_25_inst : DLH_X1 port map( G => N2995, D => N4136, Q => 
                           REGISTERS_18_25_port);
   REGISTERS_reg_18_24_inst : DLH_X1 port map( G => N2995, D => N4134, Q => 
                           REGISTERS_18_24_port);
   REGISTERS_reg_18_23_inst : DLH_X1 port map( G => N2995, D => N4132, Q => 
                           REGISTERS_18_23_port);
   REGISTERS_reg_18_22_inst : DLH_X1 port map( G => N2995, D => N4130, Q => 
                           REGISTERS_18_22_port);
   REGISTERS_reg_18_21_inst : DLH_X1 port map( G => N2995, D => N4128, Q => 
                           REGISTERS_18_21_port);
   REGISTERS_reg_18_20_inst : DLH_X1 port map( G => N2995, D => N4126, Q => 
                           REGISTERS_18_20_port);
   REGISTERS_reg_18_19_inst : DLH_X1 port map( G => N2995, D => N4124, Q => 
                           REGISTERS_18_19_port);
   REGISTERS_reg_18_18_inst : DLH_X1 port map( G => N2995, D => N4122, Q => 
                           REGISTERS_18_18_port);
   REGISTERS_reg_18_17_inst : DLH_X1 port map( G => N2995, D => N4120, Q => 
                           REGISTERS_18_17_port);
   REGISTERS_reg_18_16_inst : DLH_X1 port map( G => N2995, D => N4118, Q => 
                           REGISTERS_18_16_port);
   REGISTERS_reg_18_15_inst : DLH_X1 port map( G => N2995, D => N4116, Q => 
                           REGISTERS_18_15_port);
   REGISTERS_reg_18_14_inst : DLH_X1 port map( G => N2995, D => N4114, Q => 
                           REGISTERS_18_14_port);
   REGISTERS_reg_18_13_inst : DLH_X1 port map( G => N2995, D => N4112, Q => 
                           REGISTERS_18_13_port);
   REGISTERS_reg_18_12_inst : DLH_X1 port map( G => N2995, D => N4110, Q => 
                           REGISTERS_18_12_port);
   REGISTERS_reg_18_11_inst : DLH_X1 port map( G => N2995, D => N4108, Q => 
                           REGISTERS_18_11_port);
   REGISTERS_reg_18_10_inst : DLH_X1 port map( G => N2995, D => N4106, Q => 
                           REGISTERS_18_10_port);
   REGISTERS_reg_18_9_inst : DLH_X1 port map( G => N2995, D => N4104, Q => 
                           REGISTERS_18_9_port);
   REGISTERS_reg_18_8_inst : DLH_X1 port map( G => N2995, D => N4102, Q => 
                           REGISTERS_18_8_port);
   REGISTERS_reg_18_7_inst : DLH_X1 port map( G => N2995, D => N4100, Q => 
                           REGISTERS_18_7_port);
   REGISTERS_reg_18_6_inst : DLH_X1 port map( G => N2995, D => N4098, Q => 
                           REGISTERS_18_6_port);
   REGISTERS_reg_18_5_inst : DLH_X1 port map( G => N2995, D => N4096, Q => 
                           REGISTERS_18_5_port);
   REGISTERS_reg_18_4_inst : DLH_X1 port map( G => N2995, D => N4094, Q => 
                           REGISTERS_18_4_port);
   REGISTERS_reg_18_3_inst : DLH_X1 port map( G => N2995, D => N4092, Q => 
                           REGISTERS_18_3_port);
   REGISTERS_reg_18_2_inst : DLH_X1 port map( G => N2995, D => N4090, Q => 
                           REGISTERS_18_2_port);
   REGISTERS_reg_18_1_inst : DLH_X1 port map( G => N2995, D => N4088, Q => 
                           REGISTERS_18_1_port);
   REGISTERS_reg_18_0_inst : DLH_X1 port map( G => N2995, D => N4086, Q => 
                           REGISTERS_18_0_port);
   REGISTERS_reg_19_31_inst : DLH_X1 port map( G => N2931, D => N4148, Q => 
                           REGISTERS_19_31_port);
   REGISTERS_reg_19_30_inst : DLH_X1 port map( G => N2931, D => N4146, Q => 
                           REGISTERS_19_30_port);
   REGISTERS_reg_19_29_inst : DLH_X1 port map( G => N2931, D => N4144, Q => 
                           REGISTERS_19_29_port);
   REGISTERS_reg_19_28_inst : DLH_X1 port map( G => N2931, D => N4142, Q => 
                           REGISTERS_19_28_port);
   REGISTERS_reg_19_27_inst : DLH_X1 port map( G => N2931, D => N4140, Q => 
                           REGISTERS_19_27_port);
   REGISTERS_reg_19_26_inst : DLH_X1 port map( G => N2931, D => N4138, Q => 
                           REGISTERS_19_26_port);
   REGISTERS_reg_19_25_inst : DLH_X1 port map( G => N2931, D => N4136, Q => 
                           REGISTERS_19_25_port);
   REGISTERS_reg_19_24_inst : DLH_X1 port map( G => N2931, D => N4134, Q => 
                           REGISTERS_19_24_port);
   REGISTERS_reg_19_23_inst : DLH_X1 port map( G => N2931, D => N4132, Q => 
                           REGISTERS_19_23_port);
   REGISTERS_reg_19_22_inst : DLH_X1 port map( G => N2931, D => N4130, Q => 
                           REGISTERS_19_22_port);
   REGISTERS_reg_19_21_inst : DLH_X1 port map( G => N2931, D => N4128, Q => 
                           REGISTERS_19_21_port);
   REGISTERS_reg_19_20_inst : DLH_X1 port map( G => N2931, D => N4126, Q => 
                           REGISTERS_19_20_port);
   REGISTERS_reg_19_19_inst : DLH_X1 port map( G => N2931, D => N4124, Q => 
                           REGISTERS_19_19_port);
   REGISTERS_reg_19_18_inst : DLH_X1 port map( G => N2931, D => N4122, Q => 
                           REGISTERS_19_18_port);
   REGISTERS_reg_19_17_inst : DLH_X1 port map( G => N2931, D => N4120, Q => 
                           REGISTERS_19_17_port);
   REGISTERS_reg_19_16_inst : DLH_X1 port map( G => N2931, D => N4118, Q => 
                           REGISTERS_19_16_port);
   REGISTERS_reg_19_15_inst : DLH_X1 port map( G => N2931, D => N4116, Q => 
                           REGISTERS_19_15_port);
   REGISTERS_reg_19_14_inst : DLH_X1 port map( G => N2931, D => N4114, Q => 
                           REGISTERS_19_14_port);
   REGISTERS_reg_19_13_inst : DLH_X1 port map( G => N2931, D => N4112, Q => 
                           REGISTERS_19_13_port);
   REGISTERS_reg_19_12_inst : DLH_X1 port map( G => N2931, D => N4110, Q => 
                           REGISTERS_19_12_port);
   REGISTERS_reg_19_11_inst : DLH_X1 port map( G => N2931, D => N4108, Q => 
                           REGISTERS_19_11_port);
   REGISTERS_reg_19_10_inst : DLH_X1 port map( G => N2931, D => N4106, Q => 
                           REGISTERS_19_10_port);
   REGISTERS_reg_19_9_inst : DLH_X1 port map( G => N2931, D => N4104, Q => 
                           REGISTERS_19_9_port);
   REGISTERS_reg_19_8_inst : DLH_X1 port map( G => N2931, D => N4102, Q => 
                           REGISTERS_19_8_port);
   REGISTERS_reg_19_7_inst : DLH_X1 port map( G => N2931, D => N4100, Q => 
                           REGISTERS_19_7_port);
   REGISTERS_reg_19_6_inst : DLH_X1 port map( G => N2931, D => N4098, Q => 
                           REGISTERS_19_6_port);
   REGISTERS_reg_19_5_inst : DLH_X1 port map( G => N2931, D => N4096, Q => 
                           REGISTERS_19_5_port);
   REGISTERS_reg_19_4_inst : DLH_X1 port map( G => N2931, D => N4094, Q => 
                           REGISTERS_19_4_port);
   REGISTERS_reg_19_3_inst : DLH_X1 port map( G => N2931, D => N4092, Q => 
                           REGISTERS_19_3_port);
   REGISTERS_reg_19_2_inst : DLH_X1 port map( G => N2931, D => N4090, Q => 
                           REGISTERS_19_2_port);
   REGISTERS_reg_19_1_inst : DLH_X1 port map( G => N2931, D => N4088, Q => 
                           REGISTERS_19_1_port);
   REGISTERS_reg_19_0_inst : DLH_X1 port map( G => N2931, D => N4086, Q => 
                           REGISTERS_19_0_port);
   REGISTERS_reg_20_31_inst : DLH_X1 port map( G => N2867, D => N4148, Q => 
                           REGISTERS_20_31_port);
   REGISTERS_reg_20_30_inst : DLH_X1 port map( G => N2867, D => N4146, Q => 
                           REGISTERS_20_30_port);
   REGISTERS_reg_20_29_inst : DLH_X1 port map( G => N2867, D => N4144, Q => 
                           REGISTERS_20_29_port);
   REGISTERS_reg_20_28_inst : DLH_X1 port map( G => N2867, D => N4142, Q => 
                           REGISTERS_20_28_port);
   REGISTERS_reg_20_27_inst : DLH_X1 port map( G => N2867, D => N4140, Q => 
                           REGISTERS_20_27_port);
   REGISTERS_reg_20_26_inst : DLH_X1 port map( G => N2867, D => N4138, Q => 
                           REGISTERS_20_26_port);
   REGISTERS_reg_20_25_inst : DLH_X1 port map( G => N2867, D => N4136, Q => 
                           REGISTERS_20_25_port);
   REGISTERS_reg_20_24_inst : DLH_X1 port map( G => N2867, D => N4134, Q => 
                           REGISTERS_20_24_port);
   REGISTERS_reg_20_23_inst : DLH_X1 port map( G => N2867, D => N4132, Q => 
                           REGISTERS_20_23_port);
   REGISTERS_reg_20_22_inst : DLH_X1 port map( G => N2867, D => N4130, Q => 
                           REGISTERS_20_22_port);
   REGISTERS_reg_20_21_inst : DLH_X1 port map( G => N2867, D => N4128, Q => 
                           REGISTERS_20_21_port);
   REGISTERS_reg_20_20_inst : DLH_X1 port map( G => N2867, D => N4126, Q => 
                           REGISTERS_20_20_port);
   REGISTERS_reg_20_19_inst : DLH_X1 port map( G => N2867, D => N4124, Q => 
                           REGISTERS_20_19_port);
   REGISTERS_reg_20_18_inst : DLH_X1 port map( G => N2867, D => N4122, Q => 
                           REGISTERS_20_18_port);
   REGISTERS_reg_20_17_inst : DLH_X1 port map( G => N2867, D => N4120, Q => 
                           REGISTERS_20_17_port);
   REGISTERS_reg_20_16_inst : DLH_X1 port map( G => N2867, D => N4118, Q => 
                           REGISTERS_20_16_port);
   REGISTERS_reg_20_15_inst : DLH_X1 port map( G => N2867, D => N4116, Q => 
                           REGISTERS_20_15_port);
   REGISTERS_reg_20_14_inst : DLH_X1 port map( G => N2867, D => N4114, Q => 
                           REGISTERS_20_14_port);
   REGISTERS_reg_20_13_inst : DLH_X1 port map( G => N2867, D => N4112, Q => 
                           REGISTERS_20_13_port);
   REGISTERS_reg_20_12_inst : DLH_X1 port map( G => N2867, D => N4110, Q => 
                           REGISTERS_20_12_port);
   REGISTERS_reg_20_11_inst : DLH_X1 port map( G => N2867, D => N4108, Q => 
                           REGISTERS_20_11_port);
   REGISTERS_reg_20_10_inst : DLH_X1 port map( G => N2867, D => N4106, Q => 
                           REGISTERS_20_10_port);
   REGISTERS_reg_20_9_inst : DLH_X1 port map( G => N2867, D => N4104, Q => 
                           REGISTERS_20_9_port);
   REGISTERS_reg_20_8_inst : DLH_X1 port map( G => N2867, D => N4102, Q => 
                           REGISTERS_20_8_port);
   REGISTERS_reg_20_7_inst : DLH_X1 port map( G => N2867, D => N4100, Q => 
                           REGISTERS_20_7_port);
   REGISTERS_reg_20_6_inst : DLH_X1 port map( G => N2867, D => N4098, Q => 
                           REGISTERS_20_6_port);
   REGISTERS_reg_20_5_inst : DLH_X1 port map( G => N2867, D => N4096, Q => 
                           REGISTERS_20_5_port);
   REGISTERS_reg_20_4_inst : DLH_X1 port map( G => N2867, D => N4094, Q => 
                           REGISTERS_20_4_port);
   REGISTERS_reg_20_3_inst : DLH_X1 port map( G => N2867, D => N4092, Q => 
                           REGISTERS_20_3_port);
   REGISTERS_reg_20_2_inst : DLH_X1 port map( G => N2867, D => N4090, Q => 
                           REGISTERS_20_2_port);
   REGISTERS_reg_20_1_inst : DLH_X1 port map( G => N2867, D => N4088, Q => 
                           REGISTERS_20_1_port);
   REGISTERS_reg_20_0_inst : DLH_X1 port map( G => N2867, D => N4086, Q => 
                           REGISTERS_20_0_port);
   REGISTERS_reg_21_31_inst : DLH_X1 port map( G => N2803, D => N4148, Q => 
                           REGISTERS_21_31_port);
   REGISTERS_reg_21_30_inst : DLH_X1 port map( G => N2803, D => N4146, Q => 
                           REGISTERS_21_30_port);
   REGISTERS_reg_21_29_inst : DLH_X1 port map( G => N2803, D => N4144, Q => 
                           REGISTERS_21_29_port);
   REGISTERS_reg_21_28_inst : DLH_X1 port map( G => N2803, D => N4142, Q => 
                           REGISTERS_21_28_port);
   REGISTERS_reg_21_27_inst : DLH_X1 port map( G => N2803, D => N4140, Q => 
                           REGISTERS_21_27_port);
   REGISTERS_reg_21_26_inst : DLH_X1 port map( G => N2803, D => N4138, Q => 
                           REGISTERS_21_26_port);
   REGISTERS_reg_21_25_inst : DLH_X1 port map( G => N2803, D => N4136, Q => 
                           REGISTERS_21_25_port);
   REGISTERS_reg_21_24_inst : DLH_X1 port map( G => N2803, D => N4134, Q => 
                           REGISTERS_21_24_port);
   REGISTERS_reg_21_23_inst : DLH_X1 port map( G => N2803, D => N4132, Q => 
                           REGISTERS_21_23_port);
   REGISTERS_reg_21_22_inst : DLH_X1 port map( G => N2803, D => N4130, Q => 
                           REGISTERS_21_22_port);
   REGISTERS_reg_21_21_inst : DLH_X1 port map( G => N2803, D => N4128, Q => 
                           REGISTERS_21_21_port);
   REGISTERS_reg_21_20_inst : DLH_X1 port map( G => N2803, D => N4126, Q => 
                           REGISTERS_21_20_port);
   REGISTERS_reg_21_19_inst : DLH_X1 port map( G => N2803, D => N4124, Q => 
                           REGISTERS_21_19_port);
   REGISTERS_reg_21_18_inst : DLH_X1 port map( G => N2803, D => N4122, Q => 
                           REGISTERS_21_18_port);
   REGISTERS_reg_21_17_inst : DLH_X1 port map( G => N2803, D => N4120, Q => 
                           REGISTERS_21_17_port);
   REGISTERS_reg_21_16_inst : DLH_X1 port map( G => N2803, D => N4118, Q => 
                           REGISTERS_21_16_port);
   REGISTERS_reg_21_15_inst : DLH_X1 port map( G => N2803, D => N4116, Q => 
                           REGISTERS_21_15_port);
   REGISTERS_reg_21_14_inst : DLH_X1 port map( G => N2803, D => N4114, Q => 
                           REGISTERS_21_14_port);
   REGISTERS_reg_21_13_inst : DLH_X1 port map( G => N2803, D => N4112, Q => 
                           REGISTERS_21_13_port);
   REGISTERS_reg_21_12_inst : DLH_X1 port map( G => N2803, D => N4110, Q => 
                           REGISTERS_21_12_port);
   REGISTERS_reg_21_11_inst : DLH_X1 port map( G => N2803, D => N4108, Q => 
                           REGISTERS_21_11_port);
   REGISTERS_reg_21_10_inst : DLH_X1 port map( G => N2803, D => N4106, Q => 
                           REGISTERS_21_10_port);
   REGISTERS_reg_21_9_inst : DLH_X1 port map( G => N2803, D => N4104, Q => 
                           REGISTERS_21_9_port);
   REGISTERS_reg_21_8_inst : DLH_X1 port map( G => N2803, D => N4102, Q => 
                           REGISTERS_21_8_port);
   REGISTERS_reg_21_7_inst : DLH_X1 port map( G => N2803, D => N4100, Q => 
                           REGISTERS_21_7_port);
   REGISTERS_reg_21_6_inst : DLH_X1 port map( G => N2803, D => N4098, Q => 
                           REGISTERS_21_6_port);
   REGISTERS_reg_21_5_inst : DLH_X1 port map( G => N2803, D => N4096, Q => 
                           REGISTERS_21_5_port);
   REGISTERS_reg_21_4_inst : DLH_X1 port map( G => N2803, D => N4094, Q => 
                           REGISTERS_21_4_port);
   REGISTERS_reg_21_3_inst : DLH_X1 port map( G => N2803, D => N4092, Q => 
                           REGISTERS_21_3_port);
   REGISTERS_reg_21_2_inst : DLH_X1 port map( G => N2803, D => N4090, Q => 
                           REGISTERS_21_2_port);
   REGISTERS_reg_21_1_inst : DLH_X1 port map( G => N2803, D => N4088, Q => 
                           REGISTERS_21_1_port);
   REGISTERS_reg_21_0_inst : DLH_X1 port map( G => N2803, D => N4086, Q => 
                           REGISTERS_21_0_port);
   REGISTERS_reg_22_31_inst : DLH_X1 port map( G => N2739, D => N4148, Q => 
                           REGISTERS_22_31_port);
   REGISTERS_reg_22_30_inst : DLH_X1 port map( G => N2739, D => N4146, Q => 
                           REGISTERS_22_30_port);
   REGISTERS_reg_22_29_inst : DLH_X1 port map( G => N2739, D => N4144, Q => 
                           REGISTERS_22_29_port);
   REGISTERS_reg_22_28_inst : DLH_X1 port map( G => N2739, D => N4142, Q => 
                           REGISTERS_22_28_port);
   REGISTERS_reg_22_27_inst : DLH_X1 port map( G => N2739, D => N4140, Q => 
                           REGISTERS_22_27_port);
   REGISTERS_reg_22_26_inst : DLH_X1 port map( G => N2739, D => N4138, Q => 
                           REGISTERS_22_26_port);
   REGISTERS_reg_22_25_inst : DLH_X1 port map( G => N2739, D => N4136, Q => 
                           REGISTERS_22_25_port);
   REGISTERS_reg_22_24_inst : DLH_X1 port map( G => N2739, D => N4134, Q => 
                           REGISTERS_22_24_port);
   REGISTERS_reg_22_23_inst : DLH_X1 port map( G => N2739, D => N4132, Q => 
                           REGISTERS_22_23_port);
   REGISTERS_reg_22_22_inst : DLH_X1 port map( G => N2739, D => N4130, Q => 
                           REGISTERS_22_22_port);
   REGISTERS_reg_22_21_inst : DLH_X1 port map( G => N2739, D => N4128, Q => 
                           REGISTERS_22_21_port);
   REGISTERS_reg_22_20_inst : DLH_X1 port map( G => N2739, D => N4126, Q => 
                           REGISTERS_22_20_port);
   REGISTERS_reg_22_19_inst : DLH_X1 port map( G => N2739, D => N4124, Q => 
                           REGISTERS_22_19_port);
   REGISTERS_reg_22_18_inst : DLH_X1 port map( G => N2739, D => N4122, Q => 
                           REGISTERS_22_18_port);
   REGISTERS_reg_22_17_inst : DLH_X1 port map( G => N2739, D => N4120, Q => 
                           REGISTERS_22_17_port);
   REGISTERS_reg_22_16_inst : DLH_X1 port map( G => N2739, D => N4118, Q => 
                           REGISTERS_22_16_port);
   REGISTERS_reg_22_15_inst : DLH_X1 port map( G => N2739, D => N4116, Q => 
                           REGISTERS_22_15_port);
   REGISTERS_reg_22_14_inst : DLH_X1 port map( G => N2739, D => N4114, Q => 
                           REGISTERS_22_14_port);
   REGISTERS_reg_22_13_inst : DLH_X1 port map( G => N2739, D => N4112, Q => 
                           REGISTERS_22_13_port);
   REGISTERS_reg_22_12_inst : DLH_X1 port map( G => N2739, D => N4110, Q => 
                           REGISTERS_22_12_port);
   REGISTERS_reg_22_11_inst : DLH_X1 port map( G => N2739, D => N4108, Q => 
                           REGISTERS_22_11_port);
   REGISTERS_reg_22_10_inst : DLH_X1 port map( G => N2739, D => N4106, Q => 
                           REGISTERS_22_10_port);
   REGISTERS_reg_22_9_inst : DLH_X1 port map( G => N2739, D => N4104, Q => 
                           REGISTERS_22_9_port);
   REGISTERS_reg_22_8_inst : DLH_X1 port map( G => N2739, D => N4102, Q => 
                           REGISTERS_22_8_port);
   REGISTERS_reg_22_7_inst : DLH_X1 port map( G => N2739, D => N4100, Q => 
                           REGISTERS_22_7_port);
   REGISTERS_reg_22_6_inst : DLH_X1 port map( G => N2739, D => N4098, Q => 
                           REGISTERS_22_6_port);
   REGISTERS_reg_22_5_inst : DLH_X1 port map( G => N2739, D => N4096, Q => 
                           REGISTERS_22_5_port);
   REGISTERS_reg_22_4_inst : DLH_X1 port map( G => N2739, D => N4094, Q => 
                           REGISTERS_22_4_port);
   REGISTERS_reg_22_3_inst : DLH_X1 port map( G => N2739, D => N4092, Q => 
                           REGISTERS_22_3_port);
   REGISTERS_reg_22_2_inst : DLH_X1 port map( G => N2739, D => N4090, Q => 
                           REGISTERS_22_2_port);
   REGISTERS_reg_22_1_inst : DLH_X1 port map( G => N2739, D => N4088, Q => 
                           REGISTERS_22_1_port);
   REGISTERS_reg_22_0_inst : DLH_X1 port map( G => N2739, D => N4086, Q => 
                           REGISTERS_22_0_port);
   REGISTERS_reg_23_31_inst : DLH_X1 port map( G => N2675, D => N4148, Q => 
                           REGISTERS_23_31_port);
   REGISTERS_reg_23_30_inst : DLH_X1 port map( G => N2675, D => N4146, Q => 
                           REGISTERS_23_30_port);
   REGISTERS_reg_23_29_inst : DLH_X1 port map( G => N2675, D => N4144, Q => 
                           REGISTERS_23_29_port);
   REGISTERS_reg_23_28_inst : DLH_X1 port map( G => N2675, D => N4142, Q => 
                           REGISTERS_23_28_port);
   REGISTERS_reg_23_27_inst : DLH_X1 port map( G => N2675, D => N4140, Q => 
                           REGISTERS_23_27_port);
   REGISTERS_reg_23_26_inst : DLH_X1 port map( G => N2675, D => N4138, Q => 
                           REGISTERS_23_26_port);
   REGISTERS_reg_23_25_inst : DLH_X1 port map( G => N2675, D => N4136, Q => 
                           REGISTERS_23_25_port);
   REGISTERS_reg_23_24_inst : DLH_X1 port map( G => N2675, D => N4134, Q => 
                           REGISTERS_23_24_port);
   REGISTERS_reg_23_23_inst : DLH_X1 port map( G => N2675, D => N4132, Q => 
                           REGISTERS_23_23_port);
   REGISTERS_reg_23_22_inst : DLH_X1 port map( G => N2675, D => N4130, Q => 
                           REGISTERS_23_22_port);
   REGISTERS_reg_23_21_inst : DLH_X1 port map( G => N2675, D => N4128, Q => 
                           REGISTERS_23_21_port);
   REGISTERS_reg_23_20_inst : DLH_X1 port map( G => N2675, D => N4126, Q => 
                           REGISTERS_23_20_port);
   REGISTERS_reg_23_19_inst : DLH_X1 port map( G => N2675, D => N4124, Q => 
                           REGISTERS_23_19_port);
   REGISTERS_reg_23_18_inst : DLH_X1 port map( G => N2675, D => N4122, Q => 
                           REGISTERS_23_18_port);
   REGISTERS_reg_23_17_inst : DLH_X1 port map( G => N2675, D => N4120, Q => 
                           REGISTERS_23_17_port);
   REGISTERS_reg_23_16_inst : DLH_X1 port map( G => N2675, D => N4118, Q => 
                           REGISTERS_23_16_port);
   REGISTERS_reg_23_15_inst : DLH_X1 port map( G => N2675, D => N4116, Q => 
                           REGISTERS_23_15_port);
   REGISTERS_reg_23_14_inst : DLH_X1 port map( G => N2675, D => N4114, Q => 
                           REGISTERS_23_14_port);
   REGISTERS_reg_23_13_inst : DLH_X1 port map( G => N2675, D => N4112, Q => 
                           REGISTERS_23_13_port);
   REGISTERS_reg_23_12_inst : DLH_X1 port map( G => N2675, D => N4110, Q => 
                           REGISTERS_23_12_port);
   REGISTERS_reg_23_11_inst : DLH_X1 port map( G => N2675, D => N4108, Q => 
                           REGISTERS_23_11_port);
   REGISTERS_reg_23_10_inst : DLH_X1 port map( G => N2675, D => N4106, Q => 
                           REGISTERS_23_10_port);
   REGISTERS_reg_23_9_inst : DLH_X1 port map( G => N2675, D => N4104, Q => 
                           REGISTERS_23_9_port);
   REGISTERS_reg_23_8_inst : DLH_X1 port map( G => N2675, D => N4102, Q => 
                           REGISTERS_23_8_port);
   REGISTERS_reg_23_7_inst : DLH_X1 port map( G => N2675, D => N4100, Q => 
                           REGISTERS_23_7_port);
   REGISTERS_reg_23_6_inst : DLH_X1 port map( G => N2675, D => N4098, Q => 
                           REGISTERS_23_6_port);
   REGISTERS_reg_23_5_inst : DLH_X1 port map( G => N2675, D => N4096, Q => 
                           REGISTERS_23_5_port);
   REGISTERS_reg_23_4_inst : DLH_X1 port map( G => N2675, D => N4094, Q => 
                           REGISTERS_23_4_port);
   REGISTERS_reg_23_3_inst : DLH_X1 port map( G => N2675, D => N4092, Q => 
                           REGISTERS_23_3_port);
   REGISTERS_reg_23_2_inst : DLH_X1 port map( G => N2675, D => N4090, Q => 
                           REGISTERS_23_2_port);
   REGISTERS_reg_23_1_inst : DLH_X1 port map( G => N2675, D => N4088, Q => 
                           REGISTERS_23_1_port);
   REGISTERS_reg_23_0_inst : DLH_X1 port map( G => N2675, D => N4086, Q => 
                           REGISTERS_23_0_port);
   REGISTERS_reg_24_31_inst : DLH_X1 port map( G => N2611, D => N4148, Q => 
                           REGISTERS_24_31_port);
   REGISTERS_reg_24_30_inst : DLH_X1 port map( G => N2611, D => N4146, Q => 
                           REGISTERS_24_30_port);
   REGISTERS_reg_24_29_inst : DLH_X1 port map( G => N2611, D => N4144, Q => 
                           REGISTERS_24_29_port);
   REGISTERS_reg_24_28_inst : DLH_X1 port map( G => N2611, D => N4142, Q => 
                           REGISTERS_24_28_port);
   REGISTERS_reg_24_27_inst : DLH_X1 port map( G => N2611, D => N4140, Q => 
                           REGISTERS_24_27_port);
   REGISTERS_reg_24_26_inst : DLH_X1 port map( G => N2611, D => N4138, Q => 
                           REGISTERS_24_26_port);
   REGISTERS_reg_24_25_inst : DLH_X1 port map( G => N2611, D => N4136, Q => 
                           REGISTERS_24_25_port);
   REGISTERS_reg_24_24_inst : DLH_X1 port map( G => N2611, D => N4134, Q => 
                           REGISTERS_24_24_port);
   REGISTERS_reg_24_23_inst : DLH_X1 port map( G => N2611, D => N4132, Q => 
                           REGISTERS_24_23_port);
   REGISTERS_reg_24_22_inst : DLH_X1 port map( G => N2611, D => N4130, Q => 
                           REGISTERS_24_22_port);
   REGISTERS_reg_24_21_inst : DLH_X1 port map( G => N2611, D => N4128, Q => 
                           REGISTERS_24_21_port);
   REGISTERS_reg_24_20_inst : DLH_X1 port map( G => N2611, D => N4126, Q => 
                           REGISTERS_24_20_port);
   REGISTERS_reg_24_19_inst : DLH_X1 port map( G => N2611, D => N4124, Q => 
                           REGISTERS_24_19_port);
   REGISTERS_reg_24_18_inst : DLH_X1 port map( G => N2611, D => N4122, Q => 
                           REGISTERS_24_18_port);
   REGISTERS_reg_24_17_inst : DLH_X1 port map( G => N2611, D => N4120, Q => 
                           REGISTERS_24_17_port);
   REGISTERS_reg_24_16_inst : DLH_X1 port map( G => N2611, D => N4118, Q => 
                           REGISTERS_24_16_port);
   REGISTERS_reg_24_15_inst : DLH_X1 port map( G => N2611, D => N4116, Q => 
                           REGISTERS_24_15_port);
   REGISTERS_reg_24_14_inst : DLH_X1 port map( G => N2611, D => N4114, Q => 
                           REGISTERS_24_14_port);
   REGISTERS_reg_24_13_inst : DLH_X1 port map( G => N2611, D => N4112, Q => 
                           REGISTERS_24_13_port);
   REGISTERS_reg_24_12_inst : DLH_X1 port map( G => N2611, D => N4110, Q => 
                           REGISTERS_24_12_port);
   REGISTERS_reg_24_11_inst : DLH_X1 port map( G => N2611, D => N4108, Q => 
                           REGISTERS_24_11_port);
   REGISTERS_reg_24_10_inst : DLH_X1 port map( G => N2611, D => N4106, Q => 
                           REGISTERS_24_10_port);
   REGISTERS_reg_24_9_inst : DLH_X1 port map( G => N2611, D => N4104, Q => 
                           REGISTERS_24_9_port);
   REGISTERS_reg_24_8_inst : DLH_X1 port map( G => N2611, D => N4102, Q => 
                           REGISTERS_24_8_port);
   REGISTERS_reg_24_7_inst : DLH_X1 port map( G => N2611, D => N4100, Q => 
                           REGISTERS_24_7_port);
   REGISTERS_reg_24_6_inst : DLH_X1 port map( G => N2611, D => N4098, Q => 
                           REGISTERS_24_6_port);
   REGISTERS_reg_24_5_inst : DLH_X1 port map( G => N2611, D => N4096, Q => 
                           REGISTERS_24_5_port);
   REGISTERS_reg_24_4_inst : DLH_X1 port map( G => N2611, D => N4094, Q => 
                           REGISTERS_24_4_port);
   REGISTERS_reg_24_3_inst : DLH_X1 port map( G => N2611, D => N4092, Q => 
                           REGISTERS_24_3_port);
   REGISTERS_reg_24_2_inst : DLH_X1 port map( G => N2611, D => N4090, Q => 
                           REGISTERS_24_2_port);
   REGISTERS_reg_24_1_inst : DLH_X1 port map( G => N2611, D => N4088, Q => 
                           REGISTERS_24_1_port);
   REGISTERS_reg_24_0_inst : DLH_X1 port map( G => N2611, D => N4086, Q => 
                           REGISTERS_24_0_port);
   REGISTERS_reg_25_31_inst : DLH_X1 port map( G => N2547, D => N4148, Q => 
                           REGISTERS_25_31_port);
   REGISTERS_reg_25_30_inst : DLH_X1 port map( G => N2547, D => N4146, Q => 
                           REGISTERS_25_30_port);
   REGISTERS_reg_25_29_inst : DLH_X1 port map( G => N2547, D => N4144, Q => 
                           REGISTERS_25_29_port);
   REGISTERS_reg_25_28_inst : DLH_X1 port map( G => N2547, D => N4142, Q => 
                           REGISTERS_25_28_port);
   REGISTERS_reg_25_27_inst : DLH_X1 port map( G => N2547, D => N4140, Q => 
                           REGISTERS_25_27_port);
   REGISTERS_reg_25_26_inst : DLH_X1 port map( G => N2547, D => N4138, Q => 
                           REGISTERS_25_26_port);
   REGISTERS_reg_25_25_inst : DLH_X1 port map( G => N2547, D => N4136, Q => 
                           REGISTERS_25_25_port);
   REGISTERS_reg_25_24_inst : DLH_X1 port map( G => N2547, D => N4134, Q => 
                           REGISTERS_25_24_port);
   REGISTERS_reg_25_23_inst : DLH_X1 port map( G => N2547, D => N4132, Q => 
                           REGISTERS_25_23_port);
   REGISTERS_reg_25_22_inst : DLH_X1 port map( G => N2547, D => N4130, Q => 
                           REGISTERS_25_22_port);
   REGISTERS_reg_25_21_inst : DLH_X1 port map( G => N2547, D => N4128, Q => 
                           REGISTERS_25_21_port);
   REGISTERS_reg_25_20_inst : DLH_X1 port map( G => N2547, D => N4126, Q => 
                           REGISTERS_25_20_port);
   REGISTERS_reg_25_19_inst : DLH_X1 port map( G => N2547, D => N4124, Q => 
                           REGISTERS_25_19_port);
   REGISTERS_reg_25_18_inst : DLH_X1 port map( G => N2547, D => N4122, Q => 
                           REGISTERS_25_18_port);
   REGISTERS_reg_25_17_inst : DLH_X1 port map( G => N2547, D => N4120, Q => 
                           REGISTERS_25_17_port);
   REGISTERS_reg_25_16_inst : DLH_X1 port map( G => N2547, D => N4118, Q => 
                           REGISTERS_25_16_port);
   REGISTERS_reg_25_15_inst : DLH_X1 port map( G => N2547, D => N4116, Q => 
                           REGISTERS_25_15_port);
   REGISTERS_reg_25_14_inst : DLH_X1 port map( G => N2547, D => N4114, Q => 
                           REGISTERS_25_14_port);
   REGISTERS_reg_25_13_inst : DLH_X1 port map( G => N2547, D => N4112, Q => 
                           REGISTERS_25_13_port);
   REGISTERS_reg_25_12_inst : DLH_X1 port map( G => N2547, D => N4110, Q => 
                           REGISTERS_25_12_port);
   REGISTERS_reg_25_11_inst : DLH_X1 port map( G => N2547, D => N4108, Q => 
                           REGISTERS_25_11_port);
   REGISTERS_reg_25_10_inst : DLH_X1 port map( G => N2547, D => N4106, Q => 
                           REGISTERS_25_10_port);
   REGISTERS_reg_25_9_inst : DLH_X1 port map( G => N2547, D => N4104, Q => 
                           REGISTERS_25_9_port);
   REGISTERS_reg_25_8_inst : DLH_X1 port map( G => N2547, D => N4102, Q => 
                           REGISTERS_25_8_port);
   REGISTERS_reg_25_7_inst : DLH_X1 port map( G => N2547, D => N4100, Q => 
                           REGISTERS_25_7_port);
   REGISTERS_reg_25_6_inst : DLH_X1 port map( G => N2547, D => N4098, Q => 
                           REGISTERS_25_6_port);
   REGISTERS_reg_25_5_inst : DLH_X1 port map( G => N2547, D => N4096, Q => 
                           REGISTERS_25_5_port);
   REGISTERS_reg_25_4_inst : DLH_X1 port map( G => N2547, D => N4094, Q => 
                           REGISTERS_25_4_port);
   REGISTERS_reg_25_3_inst : DLH_X1 port map( G => N2547, D => N4092, Q => 
                           REGISTERS_25_3_port);
   REGISTERS_reg_25_2_inst : DLH_X1 port map( G => N2547, D => N4090, Q => 
                           REGISTERS_25_2_port);
   REGISTERS_reg_25_1_inst : DLH_X1 port map( G => N2547, D => N4088, Q => 
                           REGISTERS_25_1_port);
   REGISTERS_reg_25_0_inst : DLH_X1 port map( G => N2547, D => N4086, Q => 
                           REGISTERS_25_0_port);
   REGISTERS_reg_26_31_inst : DLH_X1 port map( G => N2483, D => N4148, Q => 
                           REGISTERS_26_31_port);
   REGISTERS_reg_26_30_inst : DLH_X1 port map( G => N2483, D => N4146, Q => 
                           REGISTERS_26_30_port);
   REGISTERS_reg_26_29_inst : DLH_X1 port map( G => N2483, D => N4144, Q => 
                           REGISTERS_26_29_port);
   REGISTERS_reg_26_28_inst : DLH_X1 port map( G => N2483, D => N4142, Q => 
                           REGISTERS_26_28_port);
   REGISTERS_reg_26_27_inst : DLH_X1 port map( G => N2483, D => N4140, Q => 
                           REGISTERS_26_27_port);
   REGISTERS_reg_26_26_inst : DLH_X1 port map( G => N2483, D => N4138, Q => 
                           REGISTERS_26_26_port);
   REGISTERS_reg_26_25_inst : DLH_X1 port map( G => N2483, D => N4136, Q => 
                           REGISTERS_26_25_port);
   REGISTERS_reg_26_24_inst : DLH_X1 port map( G => N2483, D => N4134, Q => 
                           REGISTERS_26_24_port);
   REGISTERS_reg_26_23_inst : DLH_X1 port map( G => N2483, D => N4132, Q => 
                           REGISTERS_26_23_port);
   REGISTERS_reg_26_22_inst : DLH_X1 port map( G => N2483, D => N4130, Q => 
                           REGISTERS_26_22_port);
   REGISTERS_reg_26_21_inst : DLH_X1 port map( G => N2483, D => N4128, Q => 
                           REGISTERS_26_21_port);
   REGISTERS_reg_26_20_inst : DLH_X1 port map( G => N2483, D => N4126, Q => 
                           REGISTERS_26_20_port);
   REGISTERS_reg_26_19_inst : DLH_X1 port map( G => N2483, D => N4124, Q => 
                           REGISTERS_26_19_port);
   REGISTERS_reg_26_18_inst : DLH_X1 port map( G => N2483, D => N4122, Q => 
                           REGISTERS_26_18_port);
   REGISTERS_reg_26_17_inst : DLH_X1 port map( G => N2483, D => N4120, Q => 
                           REGISTERS_26_17_port);
   REGISTERS_reg_26_16_inst : DLH_X1 port map( G => N2483, D => N4118, Q => 
                           REGISTERS_26_16_port);
   REGISTERS_reg_26_15_inst : DLH_X1 port map( G => N2483, D => N4116, Q => 
                           REGISTERS_26_15_port);
   REGISTERS_reg_26_14_inst : DLH_X1 port map( G => N2483, D => N4114, Q => 
                           REGISTERS_26_14_port);
   REGISTERS_reg_26_13_inst : DLH_X1 port map( G => N2483, D => N4112, Q => 
                           REGISTERS_26_13_port);
   REGISTERS_reg_26_12_inst : DLH_X1 port map( G => N2483, D => N4110, Q => 
                           REGISTERS_26_12_port);
   REGISTERS_reg_26_11_inst : DLH_X1 port map( G => N2483, D => N4108, Q => 
                           REGISTERS_26_11_port);
   REGISTERS_reg_26_10_inst : DLH_X1 port map( G => N2483, D => N4106, Q => 
                           REGISTERS_26_10_port);
   REGISTERS_reg_26_9_inst : DLH_X1 port map( G => N2483, D => N4104, Q => 
                           REGISTERS_26_9_port);
   REGISTERS_reg_26_8_inst : DLH_X1 port map( G => N2483, D => N4102, Q => 
                           REGISTERS_26_8_port);
   REGISTERS_reg_26_7_inst : DLH_X1 port map( G => N2483, D => N4100, Q => 
                           REGISTERS_26_7_port);
   REGISTERS_reg_26_6_inst : DLH_X1 port map( G => N2483, D => N4098, Q => 
                           REGISTERS_26_6_port);
   REGISTERS_reg_26_5_inst : DLH_X1 port map( G => N2483, D => N4096, Q => 
                           REGISTERS_26_5_port);
   REGISTERS_reg_26_4_inst : DLH_X1 port map( G => N2483, D => N4094, Q => 
                           REGISTERS_26_4_port);
   REGISTERS_reg_26_3_inst : DLH_X1 port map( G => N2483, D => N4092, Q => 
                           REGISTERS_26_3_port);
   REGISTERS_reg_26_2_inst : DLH_X1 port map( G => N2483, D => N4090, Q => 
                           REGISTERS_26_2_port);
   REGISTERS_reg_26_1_inst : DLH_X1 port map( G => N2483, D => N4088, Q => 
                           REGISTERS_26_1_port);
   REGISTERS_reg_26_0_inst : DLH_X1 port map( G => N2483, D => N4086, Q => 
                           REGISTERS_26_0_port);
   REGISTERS_reg_27_31_inst : DLH_X1 port map( G => N2419, D => N4148, Q => 
                           REGISTERS_27_31_port);
   REGISTERS_reg_27_30_inst : DLH_X1 port map( G => N2419, D => N4146, Q => 
                           REGISTERS_27_30_port);
   REGISTERS_reg_27_29_inst : DLH_X1 port map( G => N2419, D => N4144, Q => 
                           REGISTERS_27_29_port);
   REGISTERS_reg_27_28_inst : DLH_X1 port map( G => N2419, D => N4142, Q => 
                           REGISTERS_27_28_port);
   REGISTERS_reg_27_27_inst : DLH_X1 port map( G => N2419, D => N4140, Q => 
                           REGISTERS_27_27_port);
   REGISTERS_reg_27_26_inst : DLH_X1 port map( G => N2419, D => N4138, Q => 
                           REGISTERS_27_26_port);
   REGISTERS_reg_27_25_inst : DLH_X1 port map( G => N2419, D => N4136, Q => 
                           REGISTERS_27_25_port);
   REGISTERS_reg_27_24_inst : DLH_X1 port map( G => N2419, D => N4134, Q => 
                           REGISTERS_27_24_port);
   REGISTERS_reg_27_23_inst : DLH_X1 port map( G => N2419, D => N4132, Q => 
                           REGISTERS_27_23_port);
   REGISTERS_reg_27_22_inst : DLH_X1 port map( G => N2419, D => N4130, Q => 
                           REGISTERS_27_22_port);
   REGISTERS_reg_27_21_inst : DLH_X1 port map( G => N2419, D => N4128, Q => 
                           REGISTERS_27_21_port);
   REGISTERS_reg_27_20_inst : DLH_X1 port map( G => N2419, D => N4126, Q => 
                           REGISTERS_27_20_port);
   REGISTERS_reg_27_19_inst : DLH_X1 port map( G => N2419, D => N4124, Q => 
                           REGISTERS_27_19_port);
   REGISTERS_reg_27_18_inst : DLH_X1 port map( G => N2419, D => N4122, Q => 
                           REGISTERS_27_18_port);
   REGISTERS_reg_27_17_inst : DLH_X1 port map( G => N2419, D => N4120, Q => 
                           REGISTERS_27_17_port);
   REGISTERS_reg_27_16_inst : DLH_X1 port map( G => N2419, D => N4118, Q => 
                           REGISTERS_27_16_port);
   REGISTERS_reg_27_15_inst : DLH_X1 port map( G => N2419, D => N4116, Q => 
                           REGISTERS_27_15_port);
   REGISTERS_reg_27_14_inst : DLH_X1 port map( G => N2419, D => N4114, Q => 
                           REGISTERS_27_14_port);
   REGISTERS_reg_27_13_inst : DLH_X1 port map( G => N2419, D => N4112, Q => 
                           REGISTERS_27_13_port);
   REGISTERS_reg_27_12_inst : DLH_X1 port map( G => N2419, D => N4110, Q => 
                           REGISTERS_27_12_port);
   REGISTERS_reg_27_11_inst : DLH_X1 port map( G => N2419, D => N4108, Q => 
                           REGISTERS_27_11_port);
   REGISTERS_reg_27_10_inst : DLH_X1 port map( G => N2419, D => N4106, Q => 
                           REGISTERS_27_10_port);
   REGISTERS_reg_27_9_inst : DLH_X1 port map( G => N2419, D => N4104, Q => 
                           REGISTERS_27_9_port);
   REGISTERS_reg_27_8_inst : DLH_X1 port map( G => N2419, D => N4102, Q => 
                           REGISTERS_27_8_port);
   REGISTERS_reg_27_7_inst : DLH_X1 port map( G => N2419, D => N4100, Q => 
                           REGISTERS_27_7_port);
   REGISTERS_reg_27_6_inst : DLH_X1 port map( G => N2419, D => N4098, Q => 
                           REGISTERS_27_6_port);
   REGISTERS_reg_27_5_inst : DLH_X1 port map( G => N2419, D => N4096, Q => 
                           REGISTERS_27_5_port);
   REGISTERS_reg_27_4_inst : DLH_X1 port map( G => N2419, D => N4094, Q => 
                           REGISTERS_27_4_port);
   REGISTERS_reg_27_3_inst : DLH_X1 port map( G => N2419, D => N4092, Q => 
                           REGISTERS_27_3_port);
   REGISTERS_reg_27_2_inst : DLH_X1 port map( G => N2419, D => N4090, Q => 
                           REGISTERS_27_2_port);
   REGISTERS_reg_27_1_inst : DLH_X1 port map( G => N2419, D => N4088, Q => 
                           REGISTERS_27_1_port);
   REGISTERS_reg_27_0_inst : DLH_X1 port map( G => N2419, D => N4086, Q => 
                           REGISTERS_27_0_port);
   REGISTERS_reg_28_31_inst : DLH_X1 port map( G => N2355, D => N4148, Q => 
                           REGISTERS_28_31_port);
   REGISTERS_reg_28_30_inst : DLH_X1 port map( G => N2355, D => N4146, Q => 
                           REGISTERS_28_30_port);
   REGISTERS_reg_28_29_inst : DLH_X1 port map( G => N2355, D => N4144, Q => 
                           REGISTERS_28_29_port);
   REGISTERS_reg_28_28_inst : DLH_X1 port map( G => N2355, D => N4142, Q => 
                           REGISTERS_28_28_port);
   REGISTERS_reg_28_27_inst : DLH_X1 port map( G => N2355, D => N4140, Q => 
                           REGISTERS_28_27_port);
   REGISTERS_reg_28_26_inst : DLH_X1 port map( G => N2355, D => N4138, Q => 
                           REGISTERS_28_26_port);
   REGISTERS_reg_28_25_inst : DLH_X1 port map( G => N2355, D => N4136, Q => 
                           REGISTERS_28_25_port);
   REGISTERS_reg_28_24_inst : DLH_X1 port map( G => N2355, D => N4134, Q => 
                           REGISTERS_28_24_port);
   REGISTERS_reg_28_23_inst : DLH_X1 port map( G => N2355, D => N4132, Q => 
                           REGISTERS_28_23_port);
   REGISTERS_reg_28_22_inst : DLH_X1 port map( G => N2355, D => N4130, Q => 
                           REGISTERS_28_22_port);
   REGISTERS_reg_28_21_inst : DLH_X1 port map( G => N2355, D => N4128, Q => 
                           REGISTERS_28_21_port);
   REGISTERS_reg_28_20_inst : DLH_X1 port map( G => N2355, D => N4126, Q => 
                           REGISTERS_28_20_port);
   REGISTERS_reg_28_19_inst : DLH_X1 port map( G => N2355, D => N4124, Q => 
                           REGISTERS_28_19_port);
   REGISTERS_reg_28_18_inst : DLH_X1 port map( G => N2355, D => N4122, Q => 
                           REGISTERS_28_18_port);
   REGISTERS_reg_28_17_inst : DLH_X1 port map( G => N2355, D => N4120, Q => 
                           REGISTERS_28_17_port);
   REGISTERS_reg_28_16_inst : DLH_X1 port map( G => N2355, D => N4118, Q => 
                           REGISTERS_28_16_port);
   REGISTERS_reg_28_15_inst : DLH_X1 port map( G => N2355, D => N4116, Q => 
                           REGISTERS_28_15_port);
   REGISTERS_reg_28_14_inst : DLH_X1 port map( G => N2355, D => N4114, Q => 
                           REGISTERS_28_14_port);
   REGISTERS_reg_28_13_inst : DLH_X1 port map( G => N2355, D => N4112, Q => 
                           REGISTERS_28_13_port);
   REGISTERS_reg_28_12_inst : DLH_X1 port map( G => N2355, D => N4110, Q => 
                           REGISTERS_28_12_port);
   REGISTERS_reg_28_11_inst : DLH_X1 port map( G => N2355, D => N4108, Q => 
                           REGISTERS_28_11_port);
   REGISTERS_reg_28_10_inst : DLH_X1 port map( G => N2355, D => N4106, Q => 
                           REGISTERS_28_10_port);
   REGISTERS_reg_28_9_inst : DLH_X1 port map( G => N2355, D => N4104, Q => 
                           REGISTERS_28_9_port);
   REGISTERS_reg_28_8_inst : DLH_X1 port map( G => N2355, D => N4102, Q => 
                           REGISTERS_28_8_port);
   REGISTERS_reg_28_7_inst : DLH_X1 port map( G => N2355, D => N4100, Q => 
                           REGISTERS_28_7_port);
   REGISTERS_reg_28_6_inst : DLH_X1 port map( G => N2355, D => N4098, Q => 
                           REGISTERS_28_6_port);
   REGISTERS_reg_28_5_inst : DLH_X1 port map( G => N2355, D => N4096, Q => 
                           REGISTERS_28_5_port);
   REGISTERS_reg_28_4_inst : DLH_X1 port map( G => N2355, D => N4094, Q => 
                           REGISTERS_28_4_port);
   REGISTERS_reg_28_3_inst : DLH_X1 port map( G => N2355, D => N4092, Q => 
                           REGISTERS_28_3_port);
   REGISTERS_reg_28_2_inst : DLH_X1 port map( G => N2355, D => N4090, Q => 
                           REGISTERS_28_2_port);
   REGISTERS_reg_28_1_inst : DLH_X1 port map( G => N2355, D => N4088, Q => 
                           REGISTERS_28_1_port);
   REGISTERS_reg_28_0_inst : DLH_X1 port map( G => N2355, D => N4086, Q => 
                           REGISTERS_28_0_port);
   REGISTERS_reg_29_31_inst : DLH_X1 port map( G => N2291, D => N4148, Q => 
                           REGISTERS_29_31_port);
   REGISTERS_reg_29_30_inst : DLH_X1 port map( G => N2291, D => N4146, Q => 
                           REGISTERS_29_30_port);
   REGISTERS_reg_29_29_inst : DLH_X1 port map( G => N2291, D => N4144, Q => 
                           REGISTERS_29_29_port);
   REGISTERS_reg_29_28_inst : DLH_X1 port map( G => N2291, D => N4142, Q => 
                           REGISTERS_29_28_port);
   REGISTERS_reg_29_27_inst : DLH_X1 port map( G => N2291, D => N4140, Q => 
                           REGISTERS_29_27_port);
   REGISTERS_reg_29_26_inst : DLH_X1 port map( G => N2291, D => N4138, Q => 
                           REGISTERS_29_26_port);
   REGISTERS_reg_29_25_inst : DLH_X1 port map( G => N2291, D => N4136, Q => 
                           REGISTERS_29_25_port);
   REGISTERS_reg_29_24_inst : DLH_X1 port map( G => N2291, D => N4134, Q => 
                           REGISTERS_29_24_port);
   REGISTERS_reg_29_23_inst : DLH_X1 port map( G => N2291, D => N4132, Q => 
                           REGISTERS_29_23_port);
   REGISTERS_reg_29_22_inst : DLH_X1 port map( G => N2291, D => N4130, Q => 
                           REGISTERS_29_22_port);
   REGISTERS_reg_29_21_inst : DLH_X1 port map( G => N2291, D => N4128, Q => 
                           REGISTERS_29_21_port);
   REGISTERS_reg_29_20_inst : DLH_X1 port map( G => N2291, D => N4126, Q => 
                           REGISTERS_29_20_port);
   REGISTERS_reg_29_19_inst : DLH_X1 port map( G => N2291, D => N4124, Q => 
                           REGISTERS_29_19_port);
   REGISTERS_reg_29_18_inst : DLH_X1 port map( G => N2291, D => N4122, Q => 
                           REGISTERS_29_18_port);
   REGISTERS_reg_29_17_inst : DLH_X1 port map( G => N2291, D => N4120, Q => 
                           REGISTERS_29_17_port);
   REGISTERS_reg_29_16_inst : DLH_X1 port map( G => N2291, D => N4118, Q => 
                           REGISTERS_29_16_port);
   REGISTERS_reg_29_15_inst : DLH_X1 port map( G => N2291, D => N4116, Q => 
                           REGISTERS_29_15_port);
   REGISTERS_reg_29_14_inst : DLH_X1 port map( G => N2291, D => N4114, Q => 
                           REGISTERS_29_14_port);
   REGISTERS_reg_29_13_inst : DLH_X1 port map( G => N2291, D => N4112, Q => 
                           REGISTERS_29_13_port);
   REGISTERS_reg_29_12_inst : DLH_X1 port map( G => N2291, D => N4110, Q => 
                           REGISTERS_29_12_port);
   REGISTERS_reg_29_11_inst : DLH_X1 port map( G => N2291, D => N4108, Q => 
                           REGISTERS_29_11_port);
   REGISTERS_reg_29_10_inst : DLH_X1 port map( G => N2291, D => N4106, Q => 
                           REGISTERS_29_10_port);
   REGISTERS_reg_29_9_inst : DLH_X1 port map( G => N2291, D => N4104, Q => 
                           REGISTERS_29_9_port);
   REGISTERS_reg_29_8_inst : DLH_X1 port map( G => N2291, D => N4102, Q => 
                           REGISTERS_29_8_port);
   REGISTERS_reg_29_7_inst : DLH_X1 port map( G => N2291, D => N4100, Q => 
                           REGISTERS_29_7_port);
   REGISTERS_reg_29_6_inst : DLH_X1 port map( G => N2291, D => N4098, Q => 
                           REGISTERS_29_6_port);
   REGISTERS_reg_29_5_inst : DLH_X1 port map( G => N2291, D => N4096, Q => 
                           REGISTERS_29_5_port);
   REGISTERS_reg_29_4_inst : DLH_X1 port map( G => N2291, D => N4094, Q => 
                           REGISTERS_29_4_port);
   REGISTERS_reg_29_3_inst : DLH_X1 port map( G => N2291, D => N4092, Q => 
                           REGISTERS_29_3_port);
   REGISTERS_reg_29_2_inst : DLH_X1 port map( G => N2291, D => N4090, Q => 
                           REGISTERS_29_2_port);
   REGISTERS_reg_29_1_inst : DLH_X1 port map( G => N2291, D => N4088, Q => 
                           REGISTERS_29_1_port);
   REGISTERS_reg_29_0_inst : DLH_X1 port map( G => N2291, D => N4086, Q => 
                           REGISTERS_29_0_port);
   REGISTERS_reg_30_31_inst : DLH_X1 port map( G => N2227, D => N4148, Q => 
                           REGISTERS_30_31_port);
   REGISTERS_reg_30_30_inst : DLH_X1 port map( G => N2227, D => N4146, Q => 
                           REGISTERS_30_30_port);
   REGISTERS_reg_30_29_inst : DLH_X1 port map( G => N2227, D => N4144, Q => 
                           REGISTERS_30_29_port);
   REGISTERS_reg_30_28_inst : DLH_X1 port map( G => N2227, D => N4142, Q => 
                           REGISTERS_30_28_port);
   REGISTERS_reg_30_27_inst : DLH_X1 port map( G => N2227, D => N4140, Q => 
                           REGISTERS_30_27_port);
   REGISTERS_reg_30_26_inst : DLH_X1 port map( G => N2227, D => N4138, Q => 
                           REGISTERS_30_26_port);
   REGISTERS_reg_30_25_inst : DLH_X1 port map( G => N2227, D => N4136, Q => 
                           REGISTERS_30_25_port);
   REGISTERS_reg_30_24_inst : DLH_X1 port map( G => N2227, D => N4134, Q => 
                           REGISTERS_30_24_port);
   REGISTERS_reg_30_23_inst : DLH_X1 port map( G => N2227, D => N4132, Q => 
                           REGISTERS_30_23_port);
   REGISTERS_reg_30_22_inst : DLH_X1 port map( G => N2227, D => N4130, Q => 
                           REGISTERS_30_22_port);
   REGISTERS_reg_30_21_inst : DLH_X1 port map( G => N2227, D => N4128, Q => 
                           REGISTERS_30_21_port);
   REGISTERS_reg_30_20_inst : DLH_X1 port map( G => N2227, D => N4126, Q => 
                           REGISTERS_30_20_port);
   REGISTERS_reg_30_19_inst : DLH_X1 port map( G => N2227, D => N4124, Q => 
                           REGISTERS_30_19_port);
   REGISTERS_reg_30_18_inst : DLH_X1 port map( G => N2227, D => N4122, Q => 
                           REGISTERS_30_18_port);
   REGISTERS_reg_30_17_inst : DLH_X1 port map( G => N2227, D => N4120, Q => 
                           REGISTERS_30_17_port);
   REGISTERS_reg_30_16_inst : DLH_X1 port map( G => N2227, D => N4118, Q => 
                           REGISTERS_30_16_port);
   REGISTERS_reg_30_15_inst : DLH_X1 port map( G => N2227, D => N4116, Q => 
                           REGISTERS_30_15_port);
   REGISTERS_reg_30_14_inst : DLH_X1 port map( G => N2227, D => N4114, Q => 
                           REGISTERS_30_14_port);
   REGISTERS_reg_30_13_inst : DLH_X1 port map( G => N2227, D => N4112, Q => 
                           REGISTERS_30_13_port);
   REGISTERS_reg_30_12_inst : DLH_X1 port map( G => N2227, D => N4110, Q => 
                           REGISTERS_30_12_port);
   REGISTERS_reg_30_11_inst : DLH_X1 port map( G => N2227, D => N4108, Q => 
                           REGISTERS_30_11_port);
   REGISTERS_reg_30_10_inst : DLH_X1 port map( G => N2227, D => N4106, Q => 
                           REGISTERS_30_10_port);
   REGISTERS_reg_30_9_inst : DLH_X1 port map( G => N2227, D => N4104, Q => 
                           REGISTERS_30_9_port);
   REGISTERS_reg_30_8_inst : DLH_X1 port map( G => N2227, D => N4102, Q => 
                           REGISTERS_30_8_port);
   REGISTERS_reg_30_7_inst : DLH_X1 port map( G => N2227, D => N4100, Q => 
                           REGISTERS_30_7_port);
   REGISTERS_reg_30_6_inst : DLH_X1 port map( G => N2227, D => N4098, Q => 
                           REGISTERS_30_6_port);
   REGISTERS_reg_30_5_inst : DLH_X1 port map( G => N2227, D => N4096, Q => 
                           REGISTERS_30_5_port);
   REGISTERS_reg_30_4_inst : DLH_X1 port map( G => N2227, D => N4094, Q => 
                           REGISTERS_30_4_port);
   REGISTERS_reg_30_3_inst : DLH_X1 port map( G => N2227, D => N4092, Q => 
                           REGISTERS_30_3_port);
   REGISTERS_reg_30_2_inst : DLH_X1 port map( G => N2227, D => N4090, Q => 
                           REGISTERS_30_2_port);
   REGISTERS_reg_30_1_inst : DLH_X1 port map( G => N2227, D => N4088, Q => 
                           REGISTERS_30_1_port);
   REGISTERS_reg_30_0_inst : DLH_X1 port map( G => N2227, D => N4086, Q => 
                           REGISTERS_30_0_port);
   REGISTERS_reg_31_31_inst : DLH_X1 port map( G => N2163, D => N4148, Q => 
                           REGISTERS_31_31_port);
   REGISTERS_reg_31_30_inst : DLH_X1 port map( G => N2163, D => N4146, Q => 
                           REGISTERS_31_30_port);
   REGISTERS_reg_31_29_inst : DLH_X1 port map( G => N2163, D => N4144, Q => 
                           REGISTERS_31_29_port);
   REGISTERS_reg_31_28_inst : DLH_X1 port map( G => N2163, D => N4142, Q => 
                           REGISTERS_31_28_port);
   REGISTERS_reg_31_27_inst : DLH_X1 port map( G => N2163, D => N4140, Q => 
                           REGISTERS_31_27_port);
   REGISTERS_reg_31_26_inst : DLH_X1 port map( G => N2163, D => N4138, Q => 
                           REGISTERS_31_26_port);
   REGISTERS_reg_31_25_inst : DLH_X1 port map( G => N2163, D => N4136, Q => 
                           REGISTERS_31_25_port);
   REGISTERS_reg_31_24_inst : DLH_X1 port map( G => N2163, D => N4134, Q => 
                           REGISTERS_31_24_port);
   REGISTERS_reg_31_23_inst : DLH_X1 port map( G => N2163, D => N4132, Q => 
                           REGISTERS_31_23_port);
   REGISTERS_reg_31_22_inst : DLH_X1 port map( G => N2163, D => N4130, Q => 
                           REGISTERS_31_22_port);
   REGISTERS_reg_31_21_inst : DLH_X1 port map( G => N2163, D => N4128, Q => 
                           REGISTERS_31_21_port);
   REGISTERS_reg_31_20_inst : DLH_X1 port map( G => N2163, D => N4126, Q => 
                           REGISTERS_31_20_port);
   REGISTERS_reg_31_19_inst : DLH_X1 port map( G => N2163, D => N4124, Q => 
                           REGISTERS_31_19_port);
   REGISTERS_reg_31_18_inst : DLH_X1 port map( G => N2163, D => N4122, Q => 
                           REGISTERS_31_18_port);
   REGISTERS_reg_31_17_inst : DLH_X1 port map( G => N2163, D => N4120, Q => 
                           REGISTERS_31_17_port);
   REGISTERS_reg_31_16_inst : DLH_X1 port map( G => N2163, D => N4118, Q => 
                           REGISTERS_31_16_port);
   REGISTERS_reg_31_15_inst : DLH_X1 port map( G => N2163, D => N4116, Q => 
                           REGISTERS_31_15_port);
   REGISTERS_reg_31_14_inst : DLH_X1 port map( G => N2163, D => N4114, Q => 
                           REGISTERS_31_14_port);
   REGISTERS_reg_31_13_inst : DLH_X1 port map( G => N2163, D => N4112, Q => 
                           REGISTERS_31_13_port);
   REGISTERS_reg_31_12_inst : DLH_X1 port map( G => N2163, D => N4110, Q => 
                           REGISTERS_31_12_port);
   REGISTERS_reg_31_11_inst : DLH_X1 port map( G => N2163, D => N4108, Q => 
                           REGISTERS_31_11_port);
   REGISTERS_reg_31_10_inst : DLH_X1 port map( G => N2163, D => N4106, Q => 
                           REGISTERS_31_10_port);
   REGISTERS_reg_31_9_inst : DLH_X1 port map( G => N2163, D => N4104, Q => 
                           REGISTERS_31_9_port);
   REGISTERS_reg_31_8_inst : DLH_X1 port map( G => N2163, D => N4102, Q => 
                           REGISTERS_31_8_port);
   REGISTERS_reg_31_7_inst : DLH_X1 port map( G => N2163, D => N4100, Q => 
                           REGISTERS_31_7_port);
   REGISTERS_reg_31_6_inst : DLH_X1 port map( G => N2163, D => N4098, Q => 
                           REGISTERS_31_6_port);
   REGISTERS_reg_31_5_inst : DLH_X1 port map( G => N2163, D => N4096, Q => 
                           REGISTERS_31_5_port);
   REGISTERS_reg_31_4_inst : DLH_X1 port map( G => N2163, D => N4094, Q => 
                           REGISTERS_31_4_port);
   REGISTERS_reg_31_3_inst : DLH_X1 port map( G => N2163, D => N4092, Q => 
                           REGISTERS_31_3_port);
   REGISTERS_reg_31_2_inst : DLH_X1 port map( G => N2163, D => N4090, Q => 
                           REGISTERS_31_2_port);
   REGISTERS_reg_31_1_inst : DLH_X1 port map( G => N2163, D => N4088, Q => 
                           REGISTERS_31_1_port);
   REGISTERS_reg_31_0_inst : DLH_X1 port map( G => N2163, D => N4086, Q => 
                           REGISTERS_31_0_port);
   OUT1_reg_31_inst : DLH_X1 port map( G => N4278, D => N4215, Q => OUT1(31));
   OUT1_reg_30_inst : DLH_X1 port map( G => N4278, D => N4216, Q => OUT1(30));
   OUT1_reg_29_inst : DLH_X1 port map( G => N4278, D => N4217, Q => OUT1(29));
   OUT1_reg_28_inst : DLH_X1 port map( G => N4278, D => N4218, Q => OUT1(28));
   OUT1_reg_27_inst : DLH_X1 port map( G => N4278, D => N4219, Q => OUT1(27));
   OUT1_reg_26_inst : DLH_X1 port map( G => N4278, D => N4220, Q => OUT1(26));
   OUT1_reg_25_inst : DLH_X1 port map( G => N4278, D => N4221, Q => OUT1(25));
   OUT1_reg_24_inst : DLH_X1 port map( G => N4278, D => N4222, Q => OUT1(24));
   OUT1_reg_23_inst : DLH_X1 port map( G => N4278, D => N4223, Q => OUT1(23));
   OUT1_reg_22_inst : DLH_X1 port map( G => N4278, D => N4224, Q => OUT1(22));
   OUT1_reg_21_inst : DLH_X1 port map( G => N4278, D => N4225, Q => OUT1(21));
   OUT1_reg_20_inst : DLH_X1 port map( G => N4278, D => N4226, Q => OUT1(20));
   OUT1_reg_19_inst : DLH_X1 port map( G => N4278, D => N4227, Q => OUT1(19));
   OUT1_reg_18_inst : DLH_X1 port map( G => N4278, D => N4228, Q => OUT1(18));
   OUT1_reg_17_inst : DLH_X1 port map( G => N4278, D => N4229, Q => OUT1(17));
   OUT1_reg_16_inst : DLH_X1 port map( G => N4278, D => N4230, Q => OUT1(16));
   OUT1_reg_15_inst : DLH_X1 port map( G => N4278, D => N4231, Q => OUT1(15));
   OUT1_reg_14_inst : DLH_X1 port map( G => N4278, D => N4232, Q => OUT1(14));
   OUT1_reg_13_inst : DLH_X1 port map( G => N4278, D => N4233, Q => OUT1(13));
   OUT1_reg_12_inst : DLH_X1 port map( G => N4278, D => N4234, Q => OUT1(12));
   OUT1_reg_11_inst : DLH_X1 port map( G => N4278, D => N4235, Q => OUT1(11));
   OUT1_reg_10_inst : DLH_X1 port map( G => N4278, D => N4236, Q => OUT1(10));
   OUT1_reg_9_inst : DLH_X1 port map( G => N4278, D => N4237, Q => OUT1(9));
   OUT1_reg_8_inst : DLH_X1 port map( G => N4278, D => N4238, Q => OUT1(8));
   OUT1_reg_7_inst : DLH_X1 port map( G => N4278, D => N4239, Q => OUT1(7));
   OUT1_reg_6_inst : DLH_X1 port map( G => N4278, D => N4240, Q => OUT1(6));
   OUT1_reg_5_inst : DLH_X1 port map( G => N4278, D => N4241, Q => OUT1(5));
   OUT1_reg_4_inst : DLH_X1 port map( G => N4278, D => N4242, Q => OUT1(4));
   OUT1_reg_3_inst : DLH_X1 port map( G => N4278, D => N4243, Q => OUT1(3));
   OUT1_reg_2_inst : DLH_X1 port map( G => N4278, D => N4244, Q => OUT1(2));
   OUT1_reg_1_inst : DLH_X1 port map( G => N4278, D => N4245, Q => OUT1(1));
   OUT1_reg_0_inst : DLH_X1 port map( G => N4278, D => N4246, Q => OUT1(0));
   OUT2_reg_31_inst : DLH_X1 port map( G => N4407, D => N4344, Q => OUT2(31));
   OUT2_reg_30_inst : DLH_X1 port map( G => N4407, D => N4345, Q => OUT2(30));
   OUT2_reg_29_inst : DLH_X1 port map( G => N4407, D => N4346, Q => OUT2(29));
   OUT2_reg_28_inst : DLH_X1 port map( G => N4407, D => N4347, Q => OUT2(28));
   OUT2_reg_27_inst : DLH_X1 port map( G => N4407, D => N4348, Q => OUT2(27));
   OUT2_reg_26_inst : DLH_X1 port map( G => N4407, D => N4349, Q => OUT2(26));
   OUT2_reg_25_inst : DLH_X1 port map( G => N4407, D => N4350, Q => OUT2(25));
   OUT2_reg_24_inst : DLH_X1 port map( G => N4407, D => N4351, Q => OUT2(24));
   OUT2_reg_23_inst : DLH_X1 port map( G => N4407, D => N4352, Q => OUT2(23));
   OUT2_reg_22_inst : DLH_X1 port map( G => N4407, D => N4353, Q => OUT2(22));
   OUT2_reg_21_inst : DLH_X1 port map( G => N4407, D => N4354, Q => OUT2(21));
   OUT2_reg_20_inst : DLH_X1 port map( G => N4407, D => N4355, Q => OUT2(20));
   OUT2_reg_19_inst : DLH_X1 port map( G => N4407, D => N4356, Q => OUT2(19));
   OUT2_reg_18_inst : DLH_X1 port map( G => N4407, D => N4357, Q => OUT2(18));
   OUT2_reg_17_inst : DLH_X1 port map( G => N4407, D => N4358, Q => OUT2(17));
   OUT2_reg_16_inst : DLH_X1 port map( G => N4407, D => N4359, Q => OUT2(16));
   OUT2_reg_15_inst : DLH_X1 port map( G => N4407, D => N4360, Q => OUT2(15));
   OUT2_reg_14_inst : DLH_X1 port map( G => N4407, D => N4361, Q => OUT2(14));
   OUT2_reg_13_inst : DLH_X1 port map( G => N4407, D => N4362, Q => OUT2(13));
   OUT2_reg_12_inst : DLH_X1 port map( G => N4407, D => N4363, Q => OUT2(12));
   OUT2_reg_11_inst : DLH_X1 port map( G => N4407, D => N4364, Q => OUT2(11));
   OUT2_reg_10_inst : DLH_X1 port map( G => N4407, D => N4365, Q => OUT2(10));
   OUT2_reg_9_inst : DLH_X1 port map( G => N4407, D => N4366, Q => OUT2(9));
   OUT2_reg_8_inst : DLH_X1 port map( G => N4407, D => N4367, Q => OUT2(8));
   OUT2_reg_7_inst : DLH_X1 port map( G => N4407, D => N4368, Q => OUT2(7));
   OUT2_reg_6_inst : DLH_X1 port map( G => N4407, D => N4369, Q => OUT2(6));
   OUT2_reg_5_inst : DLH_X1 port map( G => N4407, D => N4370, Q => OUT2(5));
   OUT2_reg_4_inst : DLH_X1 port map( G => N4407, D => N4371, Q => OUT2(4));
   OUT2_reg_3_inst : DLH_X1 port map( G => N4407, D => N4372, Q => OUT2(3));
   OUT2_reg_2_inst : DLH_X1 port map( G => N4407, D => N4373, Q => OUT2(2));
   OUT2_reg_1_inst : DLH_X1 port map( G => N4407, D => N4374, Q => OUT2(1));
   OUT2_reg_0_inst : DLH_X1 port map( G => N4407, D => N4375, Q => OUT2(0));
   U35 : AND2_X1 port map( A1 => RD2, A2 => ENABLE, ZN => N4407);
   U36 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => N4375);
   U37 : NOR4_X1 port map( A1 => n4, A2 => n5, A3 => n6, A4 => n7, ZN => n3);
   U38 : OAI221_X1 port map( B1 => n8, B2 => n9, C1 => n10, C2 => n11, A => n12
                           , ZN => n7);
   U39 : AOI22_X1 port map( A1 => REGISTERS_19_0_port, A2 => n13, B1 => 
                           REGISTERS_18_0_port, B2 => n14, ZN => n12);
   U40 : OAI221_X1 port map( B1 => n15, B2 => n16, C1 => n17, C2 => n18, A => 
                           n19, ZN => n6);
   U41 : AOI22_X1 port map( A1 => REGISTERS_23_0_port, A2 => n20, B1 => 
                           REGISTERS_22_0_port, B2 => n21, ZN => n19);
   U42 : OAI221_X1 port map( B1 => n22, B2 => n23, C1 => n24, C2 => n25, A => 
                           n26, ZN => n5);
   U43 : AOI22_X1 port map( A1 => REGISTERS_27_0_port, A2 => n27, B1 => 
                           REGISTERS_26_0_port, B2 => n28, ZN => n26);
   U44 : OAI221_X1 port map( B1 => n29, B2 => n30, C1 => n31, C2 => n32, A => 
                           n33, ZN => n4);
   U45 : AOI22_X1 port map( A1 => REGISTERS_29_0_port, A2 => n34, B1 => 
                           REGISTERS_28_0_port, B2 => n35, ZN => n33);
   U46 : NOR4_X1 port map( A1 => n36, A2 => n37, A3 => n38, A4 => n39, ZN => n2
                           );
   U48 : AOI22_X1 port map( A1 => REGISTERS_3_0_port, A2 => n45, B1 => 
                           REGISTERS_2_0_port, B2 => n46, ZN => n44);
   U49 : OAI221_X1 port map( B1 => n47, B2 => n48, C1 => n49, C2 => n50, A => 
                           n51, ZN => n38);
   U50 : AOI22_X1 port map( A1 => REGISTERS_7_0_port, A2 => n52, B1 => 
                           REGISTERS_6_0_port, B2 => n53, ZN => n51);
   U51 : OAI221_X1 port map( B1 => n54, B2 => n55, C1 => n56, C2 => n57, A => 
                           n58, ZN => n37);
   U52 : AOI22_X1 port map( A1 => REGISTERS_11_0_port, A2 => n59, B1 => 
                           REGISTERS_10_0_port, B2 => n60, ZN => n58);
   U53 : OAI221_X1 port map( B1 => n61, B2 => n62, C1 => n63, C2 => n64, A => 
                           n65, ZN => n36);
   U54 : AOI22_X1 port map( A1 => REGISTERS_15_0_port, A2 => n66, B1 => 
                           REGISTERS_14_0_port, B2 => n67, ZN => n65);
   U55 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => N4374);
   U56 : NOR4_X1 port map( A1 => n70, A2 => n71, A3 => n72, A4 => n73, ZN => 
                           n69);
   U57 : OAI221_X1 port map( B1 => n8, B2 => n74, C1 => n10, C2 => n75, A => 
                           n76, ZN => n73);
   U58 : AOI22_X1 port map( A1 => REGISTERS_19_1_port, A2 => n13, B1 => 
                           REGISTERS_18_1_port, B2 => n14, ZN => n76);
   U59 : OAI221_X1 port map( B1 => n15, B2 => n77, C1 => n17, C2 => n78, A => 
                           n79, ZN => n72);
   U60 : AOI22_X1 port map( A1 => REGISTERS_23_1_port, A2 => n20, B1 => 
                           REGISTERS_22_1_port, B2 => n21, ZN => n79);
   U61 : OAI221_X1 port map( B1 => n22, B2 => n80, C1 => n24, C2 => n81, A => 
                           n82, ZN => n71);
   U62 : AOI22_X1 port map( A1 => REGISTERS_27_1_port, A2 => n27, B1 => 
                           REGISTERS_26_1_port, B2 => n28, ZN => n82);
   U63 : OAI221_X1 port map( B1 => n29, B2 => n83, C1 => n31, C2 => n84, A => 
                           n85, ZN => n70);
   U64 : AOI22_X1 port map( A1 => REGISTERS_29_1_port, A2 => n34, B1 => 
                           REGISTERS_28_1_port, B2 => n35, ZN => n85);
   U65 : NOR4_X1 port map( A1 => n86, A2 => n87, A3 => n88, A4 => n89, ZN => 
                           n68);
   U67 : AOI22_X1 port map( A1 => REGISTERS_3_1_port, A2 => n45, B1 => 
                           REGISTERS_2_1_port, B2 => n46, ZN => n92);
   U68 : OAI221_X1 port map( B1 => n47, B2 => n93, C1 => n49, C2 => n94, A => 
                           n95, ZN => n88);
   U69 : AOI22_X1 port map( A1 => REGISTERS_7_1_port, A2 => n52, B1 => 
                           REGISTERS_6_1_port, B2 => n53, ZN => n95);
   U70 : OAI221_X1 port map( B1 => n54, B2 => n96, C1 => n56, C2 => n97, A => 
                           n98, ZN => n87);
   U71 : AOI22_X1 port map( A1 => REGISTERS_11_1_port, A2 => n59, B1 => 
                           REGISTERS_10_1_port, B2 => n60, ZN => n98);
   U72 : OAI221_X1 port map( B1 => n61, B2 => n99, C1 => n63, C2 => n100, A => 
                           n101, ZN => n86);
   U73 : AOI22_X1 port map( A1 => REGISTERS_15_1_port, A2 => n66, B1 => 
                           REGISTERS_14_1_port, B2 => n67, ZN => n101);
   U74 : NAND2_X1 port map( A1 => n102, A2 => n103, ZN => N4373);
   U75 : NOR4_X1 port map( A1 => n104, A2 => n105, A3 => n106, A4 => n107, ZN 
                           => n103);
   U76 : OAI221_X1 port map( B1 => n8, B2 => n108, C1 => n10, C2 => n109, A => 
                           n110, ZN => n107);
   U77 : AOI22_X1 port map( A1 => REGISTERS_19_2_port, A2 => n13, B1 => 
                           REGISTERS_18_2_port, B2 => n14, ZN => n110);
   U78 : OAI221_X1 port map( B1 => n15, B2 => n111, C1 => n17, C2 => n112, A =>
                           n113, ZN => n106);
   U79 : AOI22_X1 port map( A1 => REGISTERS_23_2_port, A2 => n20, B1 => 
                           REGISTERS_22_2_port, B2 => n21, ZN => n113);
   U80 : OAI221_X1 port map( B1 => n22, B2 => n114, C1 => n24, C2 => n115, A =>
                           n116, ZN => n105);
   U81 : AOI22_X1 port map( A1 => REGISTERS_27_2_port, A2 => n27, B1 => 
                           REGISTERS_26_2_port, B2 => n28, ZN => n116);
   U82 : OAI221_X1 port map( B1 => n29, B2 => n117, C1 => n31, C2 => n118, A =>
                           n119, ZN => n104);
   U83 : AOI22_X1 port map( A1 => REGISTERS_29_2_port, A2 => n34, B1 => 
                           REGISTERS_28_2_port, B2 => n35, ZN => n119);
   U84 : NOR4_X1 port map( A1 => n120, A2 => n121, A3 => n122, A4 => n123, ZN 
                           => n102);
   U86 : AOI22_X1 port map( A1 => REGISTERS_3_2_port, A2 => n45, B1 => 
                           REGISTERS_2_2_port, B2 => n46, ZN => n126);
   U87 : OAI221_X1 port map( B1 => n47, B2 => n127, C1 => n49, C2 => n128, A =>
                           n129, ZN => n122);
   U88 : AOI22_X1 port map( A1 => REGISTERS_7_2_port, A2 => n52, B1 => 
                           REGISTERS_6_2_port, B2 => n53, ZN => n129);
   U89 : OAI221_X1 port map( B1 => n54, B2 => n130, C1 => n56, C2 => n131, A =>
                           n132, ZN => n121);
   U90 : AOI22_X1 port map( A1 => REGISTERS_11_2_port, A2 => n59, B1 => 
                           REGISTERS_10_2_port, B2 => n60, ZN => n132);
   U91 : OAI221_X1 port map( B1 => n61, B2 => n133, C1 => n63, C2 => n134, A =>
                           n135, ZN => n120);
   U92 : AOI22_X1 port map( A1 => REGISTERS_15_2_port, A2 => n66, B1 => 
                           REGISTERS_14_2_port, B2 => n67, ZN => n135);
   U93 : NAND2_X1 port map( A1 => n136, A2 => n137, ZN => N4372);
   U94 : NOR4_X1 port map( A1 => n138, A2 => n139, A3 => n140, A4 => n141, ZN 
                           => n137);
   U95 : OAI221_X1 port map( B1 => n8, B2 => n142, C1 => n10, C2 => n143, A => 
                           n144, ZN => n141);
   U96 : AOI22_X1 port map( A1 => REGISTERS_19_3_port, A2 => n13, B1 => 
                           REGISTERS_18_3_port, B2 => n14, ZN => n144);
   U97 : OAI221_X1 port map( B1 => n15, B2 => n145, C1 => n17, C2 => n146, A =>
                           n147, ZN => n140);
   U98 : AOI22_X1 port map( A1 => REGISTERS_23_3_port, A2 => n20, B1 => 
                           REGISTERS_22_3_port, B2 => n21, ZN => n147);
   U99 : OAI221_X1 port map( B1 => n22, B2 => n148, C1 => n24, C2 => n149, A =>
                           n150, ZN => n139);
   U100 : AOI22_X1 port map( A1 => REGISTERS_27_3_port, A2 => n27, B1 => 
                           REGISTERS_26_3_port, B2 => n28, ZN => n150);
   U101 : OAI221_X1 port map( B1 => n29, B2 => n151, C1 => n31, C2 => n152, A 
                           => n153, ZN => n138);
   U102 : AOI22_X1 port map( A1 => REGISTERS_29_3_port, A2 => n34, B1 => 
                           REGISTERS_28_3_port, B2 => n35, ZN => n153);
   U103 : NOR4_X1 port map( A1 => n154, A2 => n155, A3 => n156, A4 => n157, ZN 
                           => n136);
   U105 : AOI22_X1 port map( A1 => REGISTERS_3_3_port, A2 => n45, B1 => 
                           REGISTERS_2_3_port, B2 => n46, ZN => n160);
   U106 : OAI221_X1 port map( B1 => n47, B2 => n161, C1 => n49, C2 => n162, A 
                           => n163, ZN => n156);
   U107 : AOI22_X1 port map( A1 => REGISTERS_7_3_port, A2 => n52, B1 => 
                           REGISTERS_6_3_port, B2 => n53, ZN => n163);
   U108 : OAI221_X1 port map( B1 => n54, B2 => n164, C1 => n56, C2 => n165, A 
                           => n166, ZN => n155);
   U109 : AOI22_X1 port map( A1 => REGISTERS_11_3_port, A2 => n59, B1 => 
                           REGISTERS_10_3_port, B2 => n60, ZN => n166);
   U110 : OAI221_X1 port map( B1 => n61, B2 => n167, C1 => n63, C2 => n168, A 
                           => n169, ZN => n154);
   U111 : AOI22_X1 port map( A1 => REGISTERS_15_3_port, A2 => n66, B1 => 
                           REGISTERS_14_3_port, B2 => n67, ZN => n169);
   U112 : NAND2_X1 port map( A1 => n170, A2 => n171, ZN => N4371);
   U113 : NOR4_X1 port map( A1 => n172, A2 => n173, A3 => n174, A4 => n175, ZN 
                           => n171);
   U114 : OAI221_X1 port map( B1 => n8, B2 => n176, C1 => n10, C2 => n177, A =>
                           n178, ZN => n175);
   U115 : AOI22_X1 port map( A1 => REGISTERS_19_4_port, A2 => n13, B1 => 
                           REGISTERS_18_4_port, B2 => n14, ZN => n178);
   U116 : OAI221_X1 port map( B1 => n15, B2 => n179, C1 => n17, C2 => n180, A 
                           => n181, ZN => n174);
   U117 : AOI22_X1 port map( A1 => REGISTERS_23_4_port, A2 => n20, B1 => 
                           REGISTERS_22_4_port, B2 => n21, ZN => n181);
   U118 : OAI221_X1 port map( B1 => n22, B2 => n182, C1 => n24, C2 => n183, A 
                           => n184, ZN => n173);
   U119 : AOI22_X1 port map( A1 => REGISTERS_27_4_port, A2 => n27, B1 => 
                           REGISTERS_26_4_port, B2 => n28, ZN => n184);
   U120 : OAI221_X1 port map( B1 => n29, B2 => n185, C1 => n31, C2 => n186, A 
                           => n187, ZN => n172);
   U121 : AOI22_X1 port map( A1 => REGISTERS_29_4_port, A2 => n34, B1 => 
                           REGISTERS_28_4_port, B2 => n35, ZN => n187);
   U122 : NOR4_X1 port map( A1 => n188, A2 => n189, A3 => n190, A4 => n191, ZN 
                           => n170);
   U124 : AOI22_X1 port map( A1 => REGISTERS_3_4_port, A2 => n45, B1 => 
                           REGISTERS_2_4_port, B2 => n46, ZN => n194);
   U125 : OAI221_X1 port map( B1 => n47, B2 => n195, C1 => n49, C2 => n196, A 
                           => n197, ZN => n190);
   U126 : AOI22_X1 port map( A1 => REGISTERS_7_4_port, A2 => n52, B1 => 
                           REGISTERS_6_4_port, B2 => n53, ZN => n197);
   U127 : OAI221_X1 port map( B1 => n54, B2 => n198, C1 => n56, C2 => n199, A 
                           => n200, ZN => n189);
   U128 : AOI22_X1 port map( A1 => REGISTERS_11_4_port, A2 => n59, B1 => 
                           REGISTERS_10_4_port, B2 => n60, ZN => n200);
   U129 : OAI221_X1 port map( B1 => n61, B2 => n201, C1 => n63, C2 => n202, A 
                           => n203, ZN => n188);
   U130 : AOI22_X1 port map( A1 => REGISTERS_15_4_port, A2 => n66, B1 => 
                           REGISTERS_14_4_port, B2 => n67, ZN => n203);
   U131 : NAND2_X1 port map( A1 => n204, A2 => n205, ZN => N4370);
   U132 : NOR4_X1 port map( A1 => n206, A2 => n207, A3 => n208, A4 => n209, ZN 
                           => n205);
   U133 : OAI221_X1 port map( B1 => n8, B2 => n210, C1 => n10, C2 => n211, A =>
                           n212, ZN => n209);
   U134 : AOI22_X1 port map( A1 => REGISTERS_19_5_port, A2 => n13, B1 => 
                           REGISTERS_18_5_port, B2 => n14, ZN => n212);
   U135 : OAI221_X1 port map( B1 => n15, B2 => n213, C1 => n17, C2 => n214, A 
                           => n215, ZN => n208);
   U136 : AOI22_X1 port map( A1 => REGISTERS_23_5_port, A2 => n20, B1 => 
                           REGISTERS_22_5_port, B2 => n21, ZN => n215);
   U137 : OAI221_X1 port map( B1 => n22, B2 => n216, C1 => n24, C2 => n217, A 
                           => n218, ZN => n207);
   U138 : AOI22_X1 port map( A1 => REGISTERS_27_5_port, A2 => n27, B1 => 
                           REGISTERS_26_5_port, B2 => n28, ZN => n218);
   U139 : OAI221_X1 port map( B1 => n29, B2 => n219, C1 => n31, C2 => n220, A 
                           => n221, ZN => n206);
   U140 : AOI22_X1 port map( A1 => REGISTERS_29_5_port, A2 => n34, B1 => 
                           REGISTERS_28_5_port, B2 => n35, ZN => n221);
   U141 : NOR4_X1 port map( A1 => n222, A2 => n223, A3 => n224, A4 => n225, ZN 
                           => n204);
   U143 : AOI22_X1 port map( A1 => REGISTERS_3_5_port, A2 => n45, B1 => 
                           REGISTERS_2_5_port, B2 => n46, ZN => n228);
   U144 : OAI221_X1 port map( B1 => n47, B2 => n229, C1 => n49, C2 => n230, A 
                           => n231, ZN => n224);
   U145 : AOI22_X1 port map( A1 => REGISTERS_7_5_port, A2 => n52, B1 => 
                           REGISTERS_6_5_port, B2 => n53, ZN => n231);
   U146 : OAI221_X1 port map( B1 => n54, B2 => n232, C1 => n56, C2 => n233, A 
                           => n234, ZN => n223);
   U147 : AOI22_X1 port map( A1 => REGISTERS_11_5_port, A2 => n59, B1 => 
                           REGISTERS_10_5_port, B2 => n60, ZN => n234);
   U148 : OAI221_X1 port map( B1 => n61, B2 => n235, C1 => n63, C2 => n236, A 
                           => n237, ZN => n222);
   U149 : AOI22_X1 port map( A1 => REGISTERS_15_5_port, A2 => n66, B1 => 
                           REGISTERS_14_5_port, B2 => n67, ZN => n237);
   U150 : NAND2_X1 port map( A1 => n238, A2 => n239, ZN => N4369);
   U151 : NOR4_X1 port map( A1 => n240, A2 => n241, A3 => n242, A4 => n243, ZN 
                           => n239);
   U152 : OAI221_X1 port map( B1 => n8, B2 => n244, C1 => n10, C2 => n245, A =>
                           n246, ZN => n243);
   U153 : AOI22_X1 port map( A1 => REGISTERS_19_6_port, A2 => n13, B1 => 
                           REGISTERS_18_6_port, B2 => n14, ZN => n246);
   U154 : OAI221_X1 port map( B1 => n15, B2 => n247, C1 => n17, C2 => n248, A 
                           => n249, ZN => n242);
   U155 : AOI22_X1 port map( A1 => REGISTERS_23_6_port, A2 => n20, B1 => 
                           REGISTERS_22_6_port, B2 => n21, ZN => n249);
   U156 : OAI221_X1 port map( B1 => n22, B2 => n250, C1 => n24, C2 => n251, A 
                           => n252, ZN => n241);
   U157 : AOI22_X1 port map( A1 => REGISTERS_27_6_port, A2 => n27, B1 => 
                           REGISTERS_26_6_port, B2 => n28, ZN => n252);
   U158 : OAI221_X1 port map( B1 => n29, B2 => n253, C1 => n31, C2 => n254, A 
                           => n255, ZN => n240);
   U159 : AOI22_X1 port map( A1 => REGISTERS_29_6_port, A2 => n34, B1 => 
                           REGISTERS_28_6_port, B2 => n35, ZN => n255);
   U160 : NOR4_X1 port map( A1 => n256, A2 => n257, A3 => n258, A4 => n259, ZN 
                           => n238);
   U162 : AOI22_X1 port map( A1 => REGISTERS_3_6_port, A2 => n45, B1 => 
                           REGISTERS_2_6_port, B2 => n46, ZN => n262);
   U163 : OAI221_X1 port map( B1 => n47, B2 => n263, C1 => n49, C2 => n264, A 
                           => n265, ZN => n258);
   U164 : AOI22_X1 port map( A1 => REGISTERS_7_6_port, A2 => n52, B1 => 
                           REGISTERS_6_6_port, B2 => n53, ZN => n265);
   U165 : OAI221_X1 port map( B1 => n54, B2 => n266, C1 => n56, C2 => n267, A 
                           => n268, ZN => n257);
   U166 : AOI22_X1 port map( A1 => REGISTERS_11_6_port, A2 => n59, B1 => 
                           REGISTERS_10_6_port, B2 => n60, ZN => n268);
   U167 : OAI221_X1 port map( B1 => n61, B2 => n269, C1 => n63, C2 => n270, A 
                           => n271, ZN => n256);
   U168 : AOI22_X1 port map( A1 => REGISTERS_15_6_port, A2 => n66, B1 => 
                           REGISTERS_14_6_port, B2 => n67, ZN => n271);
   U169 : NAND2_X1 port map( A1 => n272, A2 => n273, ZN => N4368);
   U170 : NOR4_X1 port map( A1 => n274, A2 => n275, A3 => n276, A4 => n277, ZN 
                           => n273);
   U171 : OAI221_X1 port map( B1 => n8, B2 => n278, C1 => n10, C2 => n279, A =>
                           n280, ZN => n277);
   U172 : AOI22_X1 port map( A1 => REGISTERS_19_7_port, A2 => n13, B1 => 
                           REGISTERS_18_7_port, B2 => n14, ZN => n280);
   U173 : OAI221_X1 port map( B1 => n15, B2 => n281, C1 => n17, C2 => n282, A 
                           => n283, ZN => n276);
   U174 : AOI22_X1 port map( A1 => REGISTERS_23_7_port, A2 => n20, B1 => 
                           REGISTERS_22_7_port, B2 => n21, ZN => n283);
   U175 : OAI221_X1 port map( B1 => n22, B2 => n284, C1 => n24, C2 => n285, A 
                           => n286, ZN => n275);
   U176 : AOI22_X1 port map( A1 => REGISTERS_27_7_port, A2 => n27, B1 => 
                           REGISTERS_26_7_port, B2 => n28, ZN => n286);
   U177 : OAI221_X1 port map( B1 => n29, B2 => n287, C1 => n31, C2 => n288, A 
                           => n289, ZN => n274);
   U178 : AOI22_X1 port map( A1 => REGISTERS_29_7_port, A2 => n34, B1 => 
                           REGISTERS_28_7_port, B2 => n35, ZN => n289);
   U179 : NOR4_X1 port map( A1 => n290, A2 => n291, A3 => n292, A4 => n293, ZN 
                           => n272);
   U181 : AOI22_X1 port map( A1 => REGISTERS_3_7_port, A2 => n45, B1 => 
                           REGISTERS_2_7_port, B2 => n46, ZN => n296);
   U182 : OAI221_X1 port map( B1 => n47, B2 => n297, C1 => n49, C2 => n298, A 
                           => n299, ZN => n292);
   U183 : AOI22_X1 port map( A1 => REGISTERS_7_7_port, A2 => n52, B1 => 
                           REGISTERS_6_7_port, B2 => n53, ZN => n299);
   U184 : OAI221_X1 port map( B1 => n54, B2 => n300, C1 => n56, C2 => n301, A 
                           => n302, ZN => n291);
   U185 : AOI22_X1 port map( A1 => REGISTERS_11_7_port, A2 => n59, B1 => 
                           REGISTERS_10_7_port, B2 => n60, ZN => n302);
   U186 : OAI221_X1 port map( B1 => n61, B2 => n303, C1 => n63, C2 => n304, A 
                           => n305, ZN => n290);
   U187 : AOI22_X1 port map( A1 => REGISTERS_15_7_port, A2 => n66, B1 => 
                           REGISTERS_14_7_port, B2 => n67, ZN => n305);
   U188 : NAND2_X1 port map( A1 => n306, A2 => n307, ZN => N4367);
   U189 : NOR4_X1 port map( A1 => n308, A2 => n309, A3 => n310, A4 => n311, ZN 
                           => n307);
   U190 : OAI221_X1 port map( B1 => n8, B2 => n312, C1 => n10, C2 => n313, A =>
                           n314, ZN => n311);
   U191 : AOI22_X1 port map( A1 => REGISTERS_19_8_port, A2 => n13, B1 => 
                           REGISTERS_18_8_port, B2 => n14, ZN => n314);
   U192 : OAI221_X1 port map( B1 => n15, B2 => n315, C1 => n17, C2 => n316, A 
                           => n317, ZN => n310);
   U193 : AOI22_X1 port map( A1 => REGISTERS_23_8_port, A2 => n20, B1 => 
                           REGISTERS_22_8_port, B2 => n21, ZN => n317);
   U194 : OAI221_X1 port map( B1 => n22, B2 => n318, C1 => n24, C2 => n319, A 
                           => n320, ZN => n309);
   U195 : AOI22_X1 port map( A1 => REGISTERS_27_8_port, A2 => n27, B1 => 
                           REGISTERS_26_8_port, B2 => n28, ZN => n320);
   U196 : OAI221_X1 port map( B1 => n29, B2 => n321, C1 => n31, C2 => n322, A 
                           => n323, ZN => n308);
   U197 : AOI22_X1 port map( A1 => REGISTERS_29_8_port, A2 => n34, B1 => 
                           REGISTERS_28_8_port, B2 => n35, ZN => n323);
   U198 : NOR4_X1 port map( A1 => n324, A2 => n325, A3 => n326, A4 => n327, ZN 
                           => n306);
   U200 : AOI22_X1 port map( A1 => REGISTERS_3_8_port, A2 => n45, B1 => 
                           REGISTERS_2_8_port, B2 => n46, ZN => n330);
   U201 : OAI221_X1 port map( B1 => n47, B2 => n331, C1 => n49, C2 => n332, A 
                           => n333, ZN => n326);
   U202 : AOI22_X1 port map( A1 => REGISTERS_7_8_port, A2 => n52, B1 => 
                           REGISTERS_6_8_port, B2 => n53, ZN => n333);
   U203 : OAI221_X1 port map( B1 => n54, B2 => n334, C1 => n56, C2 => n335, A 
                           => n336, ZN => n325);
   U204 : AOI22_X1 port map( A1 => REGISTERS_11_8_port, A2 => n59, B1 => 
                           REGISTERS_10_8_port, B2 => n60, ZN => n336);
   U205 : OAI221_X1 port map( B1 => n61, B2 => n337, C1 => n63, C2 => n338, A 
                           => n339, ZN => n324);
   U206 : AOI22_X1 port map( A1 => REGISTERS_15_8_port, A2 => n66, B1 => 
                           REGISTERS_14_8_port, B2 => n67, ZN => n339);
   U207 : NAND2_X1 port map( A1 => n340, A2 => n341, ZN => N4366);
   U208 : NOR4_X1 port map( A1 => n342, A2 => n343, A3 => n344, A4 => n345, ZN 
                           => n341);
   U209 : OAI221_X1 port map( B1 => n8, B2 => n346, C1 => n10, C2 => n347, A =>
                           n348, ZN => n345);
   U210 : AOI22_X1 port map( A1 => REGISTERS_19_9_port, A2 => n13, B1 => 
                           REGISTERS_18_9_port, B2 => n14, ZN => n348);
   U211 : OAI221_X1 port map( B1 => n15, B2 => n349, C1 => n17, C2 => n350, A 
                           => n351, ZN => n344);
   U212 : AOI22_X1 port map( A1 => REGISTERS_23_9_port, A2 => n20, B1 => 
                           REGISTERS_22_9_port, B2 => n21, ZN => n351);
   U213 : OAI221_X1 port map( B1 => n22, B2 => n352, C1 => n24, C2 => n353, A 
                           => n354, ZN => n343);
   U214 : AOI22_X1 port map( A1 => REGISTERS_27_9_port, A2 => n27, B1 => 
                           REGISTERS_26_9_port, B2 => n28, ZN => n354);
   U215 : OAI221_X1 port map( B1 => n29, B2 => n355, C1 => n31, C2 => n356, A 
                           => n357, ZN => n342);
   U216 : AOI22_X1 port map( A1 => REGISTERS_29_9_port, A2 => n34, B1 => 
                           REGISTERS_28_9_port, B2 => n35, ZN => n357);
   U217 : NOR4_X1 port map( A1 => n358, A2 => n359, A3 => n360, A4 => n361, ZN 
                           => n340);
   U219 : AOI22_X1 port map( A1 => REGISTERS_3_9_port, A2 => n45, B1 => 
                           REGISTERS_2_9_port, B2 => n46, ZN => n364);
   U220 : OAI221_X1 port map( B1 => n47, B2 => n365, C1 => n49, C2 => n366, A 
                           => n367, ZN => n360);
   U221 : AOI22_X1 port map( A1 => REGISTERS_7_9_port, A2 => n52, B1 => 
                           REGISTERS_6_9_port, B2 => n53, ZN => n367);
   U222 : OAI221_X1 port map( B1 => n54, B2 => n368, C1 => n56, C2 => n369, A 
                           => n370, ZN => n359);
   U223 : AOI22_X1 port map( A1 => REGISTERS_11_9_port, A2 => n59, B1 => 
                           REGISTERS_10_9_port, B2 => n60, ZN => n370);
   U224 : OAI221_X1 port map( B1 => n61, B2 => n371, C1 => n63, C2 => n372, A 
                           => n373, ZN => n358);
   U225 : AOI22_X1 port map( A1 => REGISTERS_15_9_port, A2 => n66, B1 => 
                           REGISTERS_14_9_port, B2 => n67, ZN => n373);
   U226 : NAND2_X1 port map( A1 => n374, A2 => n375, ZN => N4365);
   U227 : NOR4_X1 port map( A1 => n376, A2 => n377, A3 => n378, A4 => n379, ZN 
                           => n375);
   U228 : OAI221_X1 port map( B1 => n8, B2 => n380, C1 => n10, C2 => n381, A =>
                           n382, ZN => n379);
   U229 : AOI22_X1 port map( A1 => REGISTERS_19_10_port, A2 => n13, B1 => 
                           REGISTERS_18_10_port, B2 => n14, ZN => n382);
   U230 : OAI221_X1 port map( B1 => n15, B2 => n383, C1 => n17, C2 => n384, A 
                           => n385, ZN => n378);
   U231 : AOI22_X1 port map( A1 => REGISTERS_23_10_port, A2 => n20, B1 => 
                           REGISTERS_22_10_port, B2 => n21, ZN => n385);
   U232 : OAI221_X1 port map( B1 => n22, B2 => n386, C1 => n24, C2 => n387, A 
                           => n388, ZN => n377);
   U233 : AOI22_X1 port map( A1 => REGISTERS_27_10_port, A2 => n27, B1 => 
                           REGISTERS_26_10_port, B2 => n28, ZN => n388);
   U234 : OAI221_X1 port map( B1 => n29, B2 => n389, C1 => n31, C2 => n390, A 
                           => n391, ZN => n376);
   U235 : AOI22_X1 port map( A1 => REGISTERS_29_10_port, A2 => n34, B1 => 
                           REGISTERS_28_10_port, B2 => n35, ZN => n391);
   U236 : NOR4_X1 port map( A1 => n392, A2 => n393, A3 => n394, A4 => n395, ZN 
                           => n374);
   U238 : AOI22_X1 port map( A1 => REGISTERS_3_10_port, A2 => n45, B1 => 
                           REGISTERS_2_10_port, B2 => n46, ZN => n398);
   U239 : OAI221_X1 port map( B1 => n47, B2 => n399, C1 => n49, C2 => n400, A 
                           => n401, ZN => n394);
   U240 : AOI22_X1 port map( A1 => REGISTERS_7_10_port, A2 => n52, B1 => 
                           REGISTERS_6_10_port, B2 => n53, ZN => n401);
   U241 : OAI221_X1 port map( B1 => n54, B2 => n402, C1 => n56, C2 => n403, A 
                           => n404, ZN => n393);
   U242 : AOI22_X1 port map( A1 => REGISTERS_11_10_port, A2 => n59, B1 => 
                           REGISTERS_10_10_port, B2 => n60, ZN => n404);
   U243 : OAI221_X1 port map( B1 => n61, B2 => n405, C1 => n63, C2 => n406, A 
                           => n407, ZN => n392);
   U244 : AOI22_X1 port map( A1 => REGISTERS_15_10_port, A2 => n66, B1 => 
                           REGISTERS_14_10_port, B2 => n67, ZN => n407);
   U245 : NAND2_X1 port map( A1 => n408, A2 => n409, ZN => N4364);
   U246 : NOR4_X1 port map( A1 => n410, A2 => n411, A3 => n412, A4 => n413, ZN 
                           => n409);
   U247 : OAI221_X1 port map( B1 => n8, B2 => n414, C1 => n10, C2 => n415, A =>
                           n416, ZN => n413);
   U248 : AOI22_X1 port map( A1 => REGISTERS_19_11_port, A2 => n13, B1 => 
                           REGISTERS_18_11_port, B2 => n14, ZN => n416);
   U249 : OAI221_X1 port map( B1 => n15, B2 => n417, C1 => n17, C2 => n418, A 
                           => n419, ZN => n412);
   U250 : AOI22_X1 port map( A1 => REGISTERS_23_11_port, A2 => n20, B1 => 
                           REGISTERS_22_11_port, B2 => n21, ZN => n419);
   U251 : OAI221_X1 port map( B1 => n22, B2 => n420, C1 => n24, C2 => n421, A 
                           => n422, ZN => n411);
   U252 : AOI22_X1 port map( A1 => REGISTERS_27_11_port, A2 => n27, B1 => 
                           REGISTERS_26_11_port, B2 => n28, ZN => n422);
   U253 : OAI221_X1 port map( B1 => n29, B2 => n423, C1 => n31, C2 => n424, A 
                           => n425, ZN => n410);
   U254 : AOI22_X1 port map( A1 => REGISTERS_29_11_port, A2 => n34, B1 => 
                           REGISTERS_28_11_port, B2 => n35, ZN => n425);
   U255 : NOR4_X1 port map( A1 => n426, A2 => n427, A3 => n428, A4 => n429, ZN 
                           => n408);
   U257 : AOI22_X1 port map( A1 => REGISTERS_3_11_port, A2 => n45, B1 => 
                           REGISTERS_2_11_port, B2 => n46, ZN => n432);
   U258 : OAI221_X1 port map( B1 => n47, B2 => n433, C1 => n49, C2 => n434, A 
                           => n435, ZN => n428);
   U259 : AOI22_X1 port map( A1 => REGISTERS_7_11_port, A2 => n52, B1 => 
                           REGISTERS_6_11_port, B2 => n53, ZN => n435);
   U260 : OAI221_X1 port map( B1 => n54, B2 => n436, C1 => n56, C2 => n437, A 
                           => n438, ZN => n427);
   U261 : AOI22_X1 port map( A1 => REGISTERS_11_11_port, A2 => n59, B1 => 
                           REGISTERS_10_11_port, B2 => n60, ZN => n438);
   U262 : OAI221_X1 port map( B1 => n61, B2 => n439, C1 => n63, C2 => n440, A 
                           => n441, ZN => n426);
   U263 : AOI22_X1 port map( A1 => REGISTERS_15_11_port, A2 => n66, B1 => 
                           REGISTERS_14_11_port, B2 => n67, ZN => n441);
   U264 : NAND2_X1 port map( A1 => n442, A2 => n443, ZN => N4363);
   U265 : NOR4_X1 port map( A1 => n444, A2 => n445, A3 => n446, A4 => n447, ZN 
                           => n443);
   U266 : OAI221_X1 port map( B1 => n8, B2 => n448, C1 => n10, C2 => n449, A =>
                           n450, ZN => n447);
   U267 : AOI22_X1 port map( A1 => REGISTERS_19_12_port, A2 => n13, B1 => 
                           REGISTERS_18_12_port, B2 => n14, ZN => n450);
   U268 : OAI221_X1 port map( B1 => n15, B2 => n451, C1 => n17, C2 => n452, A 
                           => n453, ZN => n446);
   U269 : AOI22_X1 port map( A1 => REGISTERS_23_12_port, A2 => n20, B1 => 
                           REGISTERS_22_12_port, B2 => n21, ZN => n453);
   U270 : OAI221_X1 port map( B1 => n22, B2 => n454, C1 => n24, C2 => n455, A 
                           => n456, ZN => n445);
   U271 : AOI22_X1 port map( A1 => REGISTERS_27_12_port, A2 => n27, B1 => 
                           REGISTERS_26_12_port, B2 => n28, ZN => n456);
   U272 : OAI221_X1 port map( B1 => n29, B2 => n457, C1 => n31, C2 => n458, A 
                           => n459, ZN => n444);
   U273 : AOI22_X1 port map( A1 => REGISTERS_29_12_port, A2 => n34, B1 => 
                           REGISTERS_28_12_port, B2 => n35, ZN => n459);
   U274 : NOR4_X1 port map( A1 => n460, A2 => n461, A3 => n462, A4 => n463, ZN 
                           => n442);
   U276 : AOI22_X1 port map( A1 => REGISTERS_3_12_port, A2 => n45, B1 => 
                           REGISTERS_2_12_port, B2 => n46, ZN => n466);
   U277 : OAI221_X1 port map( B1 => n47, B2 => n467, C1 => n49, C2 => n468, A 
                           => n469, ZN => n462);
   U278 : AOI22_X1 port map( A1 => REGISTERS_7_12_port, A2 => n52, B1 => 
                           REGISTERS_6_12_port, B2 => n53, ZN => n469);
   U279 : OAI221_X1 port map( B1 => n54, B2 => n470, C1 => n56, C2 => n471, A 
                           => n472, ZN => n461);
   U280 : AOI22_X1 port map( A1 => REGISTERS_11_12_port, A2 => n59, B1 => 
                           REGISTERS_10_12_port, B2 => n60, ZN => n472);
   U281 : OAI221_X1 port map( B1 => n61, B2 => n473, C1 => n63, C2 => n474, A 
                           => n475, ZN => n460);
   U282 : AOI22_X1 port map( A1 => REGISTERS_15_12_port, A2 => n66, B1 => 
                           REGISTERS_14_12_port, B2 => n67, ZN => n475);
   U283 : NAND2_X1 port map( A1 => n476, A2 => n477, ZN => N4362);
   U284 : NOR4_X1 port map( A1 => n478, A2 => n479, A3 => n480, A4 => n481, ZN 
                           => n477);
   U285 : OAI221_X1 port map( B1 => n8, B2 => n482, C1 => n10, C2 => n483, A =>
                           n484, ZN => n481);
   U286 : AOI22_X1 port map( A1 => REGISTERS_19_13_port, A2 => n13, B1 => 
                           REGISTERS_18_13_port, B2 => n14, ZN => n484);
   U287 : OAI221_X1 port map( B1 => n15, B2 => n485, C1 => n17, C2 => n486, A 
                           => n487, ZN => n480);
   U288 : AOI22_X1 port map( A1 => REGISTERS_23_13_port, A2 => n20, B1 => 
                           REGISTERS_22_13_port, B2 => n21, ZN => n487);
   U289 : OAI221_X1 port map( B1 => n22, B2 => n488, C1 => n24, C2 => n489, A 
                           => n490, ZN => n479);
   U290 : AOI22_X1 port map( A1 => REGISTERS_27_13_port, A2 => n27, B1 => 
                           REGISTERS_26_13_port, B2 => n28, ZN => n490);
   U291 : OAI221_X1 port map( B1 => n29, B2 => n491, C1 => n31, C2 => n492, A 
                           => n493, ZN => n478);
   U292 : AOI22_X1 port map( A1 => REGISTERS_29_13_port, A2 => n34, B1 => 
                           REGISTERS_28_13_port, B2 => n35, ZN => n493);
   U293 : NOR4_X1 port map( A1 => n494, A2 => n495, A3 => n496, A4 => n497, ZN 
                           => n476);
   U295 : AOI22_X1 port map( A1 => REGISTERS_3_13_port, A2 => n45, B1 => 
                           REGISTERS_2_13_port, B2 => n46, ZN => n500);
   U296 : OAI221_X1 port map( B1 => n47, B2 => n501, C1 => n49, C2 => n502, A 
                           => n503, ZN => n496);
   U297 : AOI22_X1 port map( A1 => REGISTERS_7_13_port, A2 => n52, B1 => 
                           REGISTERS_6_13_port, B2 => n53, ZN => n503);
   U298 : OAI221_X1 port map( B1 => n54, B2 => n504, C1 => n56, C2 => n505, A 
                           => n506, ZN => n495);
   U299 : AOI22_X1 port map( A1 => REGISTERS_11_13_port, A2 => n59, B1 => 
                           REGISTERS_10_13_port, B2 => n60, ZN => n506);
   U300 : OAI221_X1 port map( B1 => n61, B2 => n507, C1 => n63, C2 => n508, A 
                           => n509, ZN => n494);
   U301 : AOI22_X1 port map( A1 => REGISTERS_15_13_port, A2 => n66, B1 => 
                           REGISTERS_14_13_port, B2 => n67, ZN => n509);
   U302 : NAND2_X1 port map( A1 => n510, A2 => n511, ZN => N4361);
   U303 : NOR4_X1 port map( A1 => n512, A2 => n513, A3 => n514, A4 => n515, ZN 
                           => n511);
   U304 : OAI221_X1 port map( B1 => n8, B2 => n516, C1 => n10, C2 => n517, A =>
                           n518, ZN => n515);
   U305 : AOI22_X1 port map( A1 => REGISTERS_19_14_port, A2 => n13, B1 => 
                           REGISTERS_18_14_port, B2 => n14, ZN => n518);
   U306 : OAI221_X1 port map( B1 => n15, B2 => n519, C1 => n17, C2 => n520, A 
                           => n521, ZN => n514);
   U307 : AOI22_X1 port map( A1 => REGISTERS_23_14_port, A2 => n20, B1 => 
                           REGISTERS_22_14_port, B2 => n21, ZN => n521);
   U308 : OAI221_X1 port map( B1 => n22, B2 => n522, C1 => n24, C2 => n523, A 
                           => n524, ZN => n513);
   U309 : AOI22_X1 port map( A1 => REGISTERS_27_14_port, A2 => n27, B1 => 
                           REGISTERS_26_14_port, B2 => n28, ZN => n524);
   U310 : OAI221_X1 port map( B1 => n29, B2 => n525, C1 => n31, C2 => n526, A 
                           => n527, ZN => n512);
   U311 : AOI22_X1 port map( A1 => REGISTERS_29_14_port, A2 => n34, B1 => 
                           REGISTERS_28_14_port, B2 => n35, ZN => n527);
   U312 : NOR4_X1 port map( A1 => n528, A2 => n529, A3 => n530, A4 => n531, ZN 
                           => n510);
   U314 : AOI22_X1 port map( A1 => REGISTERS_3_14_port, A2 => n45, B1 => 
                           REGISTERS_2_14_port, B2 => n46, ZN => n534);
   U315 : OAI221_X1 port map( B1 => n47, B2 => n535, C1 => n49, C2 => n536, A 
                           => n537, ZN => n530);
   U316 : AOI22_X1 port map( A1 => REGISTERS_7_14_port, A2 => n52, B1 => 
                           REGISTERS_6_14_port, B2 => n53, ZN => n537);
   U317 : OAI221_X1 port map( B1 => n54, B2 => n538, C1 => n56, C2 => n539, A 
                           => n540, ZN => n529);
   U318 : AOI22_X1 port map( A1 => REGISTERS_11_14_port, A2 => n59, B1 => 
                           REGISTERS_10_14_port, B2 => n60, ZN => n540);
   U319 : OAI221_X1 port map( B1 => n61, B2 => n541, C1 => n63, C2 => n542, A 
                           => n543, ZN => n528);
   U320 : AOI22_X1 port map( A1 => REGISTERS_15_14_port, A2 => n66, B1 => 
                           REGISTERS_14_14_port, B2 => n67, ZN => n543);
   U321 : NAND2_X1 port map( A1 => n544, A2 => n545, ZN => N4360);
   U322 : NOR4_X1 port map( A1 => n546, A2 => n547, A3 => n548, A4 => n549, ZN 
                           => n545);
   U323 : OAI221_X1 port map( B1 => n8, B2 => n550, C1 => n10, C2 => n551, A =>
                           n552, ZN => n549);
   U324 : AOI22_X1 port map( A1 => REGISTERS_19_15_port, A2 => n13, B1 => 
                           REGISTERS_18_15_port, B2 => n14, ZN => n552);
   U325 : OAI221_X1 port map( B1 => n15, B2 => n553, C1 => n17, C2 => n554, A 
                           => n555, ZN => n548);
   U326 : AOI22_X1 port map( A1 => REGISTERS_23_15_port, A2 => n20, B1 => 
                           REGISTERS_22_15_port, B2 => n21, ZN => n555);
   U327 : OAI221_X1 port map( B1 => n22, B2 => n556, C1 => n24, C2 => n557, A 
                           => n558, ZN => n547);
   U328 : AOI22_X1 port map( A1 => REGISTERS_27_15_port, A2 => n27, B1 => 
                           REGISTERS_26_15_port, B2 => n28, ZN => n558);
   U329 : OAI221_X1 port map( B1 => n29, B2 => n559, C1 => n31, C2 => n560, A 
                           => n561, ZN => n546);
   U330 : AOI22_X1 port map( A1 => REGISTERS_29_15_port, A2 => n34, B1 => 
                           REGISTERS_28_15_port, B2 => n35, ZN => n561);
   U331 : NOR4_X1 port map( A1 => n562, A2 => n563, A3 => n564, A4 => n565, ZN 
                           => n544);
   U333 : AOI22_X1 port map( A1 => REGISTERS_3_15_port, A2 => n45, B1 => 
                           REGISTERS_2_15_port, B2 => n46, ZN => n568);
   U334 : OAI221_X1 port map( B1 => n47, B2 => n569, C1 => n49, C2 => n570, A 
                           => n571, ZN => n564);
   U335 : AOI22_X1 port map( A1 => REGISTERS_7_15_port, A2 => n52, B1 => 
                           REGISTERS_6_15_port, B2 => n53, ZN => n571);
   U336 : OAI221_X1 port map( B1 => n54, B2 => n572, C1 => n56, C2 => n573, A 
                           => n574, ZN => n563);
   U337 : AOI22_X1 port map( A1 => REGISTERS_11_15_port, A2 => n59, B1 => 
                           REGISTERS_10_15_port, B2 => n60, ZN => n574);
   U338 : OAI221_X1 port map( B1 => n61, B2 => n575, C1 => n63, C2 => n576, A 
                           => n577, ZN => n562);
   U339 : AOI22_X1 port map( A1 => REGISTERS_15_15_port, A2 => n66, B1 => 
                           REGISTERS_14_15_port, B2 => n67, ZN => n577);
   U340 : NAND2_X1 port map( A1 => n578, A2 => n579, ZN => N4359);
   U341 : NOR4_X1 port map( A1 => n580, A2 => n581, A3 => n582, A4 => n583, ZN 
                           => n579);
   U342 : OAI221_X1 port map( B1 => n8, B2 => n584, C1 => n10, C2 => n585, A =>
                           n586, ZN => n583);
   U343 : AOI22_X1 port map( A1 => REGISTERS_19_16_port, A2 => n13, B1 => 
                           REGISTERS_18_16_port, B2 => n14, ZN => n586);
   U344 : OAI221_X1 port map( B1 => n15, B2 => n587, C1 => n17, C2 => n588, A 
                           => n589, ZN => n582);
   U345 : AOI22_X1 port map( A1 => REGISTERS_23_16_port, A2 => n20, B1 => 
                           REGISTERS_22_16_port, B2 => n21, ZN => n589);
   U346 : OAI221_X1 port map( B1 => n22, B2 => n590, C1 => n24, C2 => n591, A 
                           => n592, ZN => n581);
   U347 : AOI22_X1 port map( A1 => REGISTERS_27_16_port, A2 => n27, B1 => 
                           REGISTERS_26_16_port, B2 => n28, ZN => n592);
   U348 : OAI221_X1 port map( B1 => n29, B2 => n593, C1 => n31, C2 => n594, A 
                           => n595, ZN => n580);
   U349 : AOI22_X1 port map( A1 => REGISTERS_29_16_port, A2 => n34, B1 => 
                           REGISTERS_28_16_port, B2 => n35, ZN => n595);
   U350 : NOR4_X1 port map( A1 => n596, A2 => n597, A3 => n598, A4 => n599, ZN 
                           => n578);
   U352 : AOI22_X1 port map( A1 => REGISTERS_3_16_port, A2 => n45, B1 => 
                           REGISTERS_2_16_port, B2 => n46, ZN => n602);
   U353 : OAI221_X1 port map( B1 => n47, B2 => n603, C1 => n49, C2 => n604, A 
                           => n605, ZN => n598);
   U354 : AOI22_X1 port map( A1 => REGISTERS_7_16_port, A2 => n52, B1 => 
                           REGISTERS_6_16_port, B2 => n53, ZN => n605);
   U355 : OAI221_X1 port map( B1 => n54, B2 => n606, C1 => n56, C2 => n607, A 
                           => n608, ZN => n597);
   U356 : AOI22_X1 port map( A1 => REGISTERS_11_16_port, A2 => n59, B1 => 
                           REGISTERS_10_16_port, B2 => n60, ZN => n608);
   U357 : OAI221_X1 port map( B1 => n61, B2 => n609, C1 => n63, C2 => n610, A 
                           => n611, ZN => n596);
   U358 : AOI22_X1 port map( A1 => REGISTERS_15_16_port, A2 => n66, B1 => 
                           REGISTERS_14_16_port, B2 => n67, ZN => n611);
   U359 : NAND2_X1 port map( A1 => n612, A2 => n613, ZN => N4358);
   U360 : NOR4_X1 port map( A1 => n614, A2 => n615, A3 => n616, A4 => n617, ZN 
                           => n613);
   U361 : OAI221_X1 port map( B1 => n8, B2 => n618, C1 => n10, C2 => n619, A =>
                           n620, ZN => n617);
   U362 : AOI22_X1 port map( A1 => REGISTERS_19_17_port, A2 => n13, B1 => 
                           REGISTERS_18_17_port, B2 => n14, ZN => n620);
   U363 : OAI221_X1 port map( B1 => n15, B2 => n621, C1 => n17, C2 => n622, A 
                           => n623, ZN => n616);
   U364 : AOI22_X1 port map( A1 => REGISTERS_23_17_port, A2 => n20, B1 => 
                           REGISTERS_22_17_port, B2 => n21, ZN => n623);
   U365 : OAI221_X1 port map( B1 => n22, B2 => n624, C1 => n24, C2 => n625, A 
                           => n626, ZN => n615);
   U366 : AOI22_X1 port map( A1 => REGISTERS_27_17_port, A2 => n27, B1 => 
                           REGISTERS_26_17_port, B2 => n28, ZN => n626);
   U367 : OAI221_X1 port map( B1 => n29, B2 => n627, C1 => n31, C2 => n628, A 
                           => n629, ZN => n614);
   U368 : AOI22_X1 port map( A1 => REGISTERS_29_17_port, A2 => n34, B1 => 
                           REGISTERS_28_17_port, B2 => n35, ZN => n629);
   U369 : NOR4_X1 port map( A1 => n630, A2 => n631, A3 => n632, A4 => n633, ZN 
                           => n612);
   U371 : AOI22_X1 port map( A1 => REGISTERS_3_17_port, A2 => n45, B1 => 
                           REGISTERS_2_17_port, B2 => n46, ZN => n636);
   U372 : OAI221_X1 port map( B1 => n47, B2 => n637, C1 => n49, C2 => n638, A 
                           => n639, ZN => n632);
   U373 : AOI22_X1 port map( A1 => REGISTERS_7_17_port, A2 => n52, B1 => 
                           REGISTERS_6_17_port, B2 => n53, ZN => n639);
   U374 : OAI221_X1 port map( B1 => n54, B2 => n640, C1 => n56, C2 => n641, A 
                           => n642, ZN => n631);
   U375 : AOI22_X1 port map( A1 => REGISTERS_11_17_port, A2 => n59, B1 => 
                           REGISTERS_10_17_port, B2 => n60, ZN => n642);
   U376 : OAI221_X1 port map( B1 => n61, B2 => n643, C1 => n63, C2 => n644, A 
                           => n645, ZN => n630);
   U377 : AOI22_X1 port map( A1 => REGISTERS_15_17_port, A2 => n66, B1 => 
                           REGISTERS_14_17_port, B2 => n67, ZN => n645);
   U378 : NAND2_X1 port map( A1 => n646, A2 => n647, ZN => N4357);
   U379 : NOR4_X1 port map( A1 => n648, A2 => n649, A3 => n650, A4 => n651, ZN 
                           => n647);
   U380 : OAI221_X1 port map( B1 => n8, B2 => n652, C1 => n10, C2 => n653, A =>
                           n654, ZN => n651);
   U381 : AOI22_X1 port map( A1 => REGISTERS_19_18_port, A2 => n13, B1 => 
                           REGISTERS_18_18_port, B2 => n14, ZN => n654);
   U382 : OAI221_X1 port map( B1 => n15, B2 => n655, C1 => n17, C2 => n656, A 
                           => n657, ZN => n650);
   U383 : AOI22_X1 port map( A1 => REGISTERS_23_18_port, A2 => n20, B1 => 
                           REGISTERS_22_18_port, B2 => n21, ZN => n657);
   U384 : OAI221_X1 port map( B1 => n22, B2 => n658, C1 => n24, C2 => n659, A 
                           => n660, ZN => n649);
   U385 : AOI22_X1 port map( A1 => REGISTERS_27_18_port, A2 => n27, B1 => 
                           REGISTERS_26_18_port, B2 => n28, ZN => n660);
   U386 : OAI221_X1 port map( B1 => n29, B2 => n661, C1 => n31, C2 => n662, A 
                           => n663, ZN => n648);
   U387 : AOI22_X1 port map( A1 => REGISTERS_29_18_port, A2 => n34, B1 => 
                           REGISTERS_28_18_port, B2 => n35, ZN => n663);
   U388 : NOR4_X1 port map( A1 => n664, A2 => n665, A3 => n666, A4 => n667, ZN 
                           => n646);
   U390 : AOI22_X1 port map( A1 => REGISTERS_3_18_port, A2 => n45, B1 => 
                           REGISTERS_2_18_port, B2 => n46, ZN => n670);
   U391 : OAI221_X1 port map( B1 => n47, B2 => n671, C1 => n49, C2 => n672, A 
                           => n673, ZN => n666);
   U392 : AOI22_X1 port map( A1 => REGISTERS_7_18_port, A2 => n52, B1 => 
                           REGISTERS_6_18_port, B2 => n53, ZN => n673);
   U393 : OAI221_X1 port map( B1 => n54, B2 => n674, C1 => n56, C2 => n675, A 
                           => n676, ZN => n665);
   U394 : AOI22_X1 port map( A1 => REGISTERS_11_18_port, A2 => n59, B1 => 
                           REGISTERS_10_18_port, B2 => n60, ZN => n676);
   U395 : OAI221_X1 port map( B1 => n61, B2 => n677, C1 => n63, C2 => n678, A 
                           => n679, ZN => n664);
   U396 : AOI22_X1 port map( A1 => REGISTERS_15_18_port, A2 => n66, B1 => 
                           REGISTERS_14_18_port, B2 => n67, ZN => n679);
   U397 : NAND2_X1 port map( A1 => n680, A2 => n681, ZN => N4356);
   U398 : NOR4_X1 port map( A1 => n682, A2 => n683, A3 => n684, A4 => n685, ZN 
                           => n681);
   U399 : OAI221_X1 port map( B1 => n8, B2 => n686, C1 => n10, C2 => n687, A =>
                           n688, ZN => n685);
   U400 : AOI22_X1 port map( A1 => REGISTERS_19_19_port, A2 => n13, B1 => 
                           REGISTERS_18_19_port, B2 => n14, ZN => n688);
   U401 : OAI221_X1 port map( B1 => n15, B2 => n689, C1 => n17, C2 => n690, A 
                           => n691, ZN => n684);
   U402 : AOI22_X1 port map( A1 => REGISTERS_23_19_port, A2 => n20, B1 => 
                           REGISTERS_22_19_port, B2 => n21, ZN => n691);
   U403 : OAI221_X1 port map( B1 => n22, B2 => n692, C1 => n24, C2 => n693, A 
                           => n694, ZN => n683);
   U404 : AOI22_X1 port map( A1 => REGISTERS_27_19_port, A2 => n27, B1 => 
                           REGISTERS_26_19_port, B2 => n28, ZN => n694);
   U405 : OAI221_X1 port map( B1 => n29, B2 => n695, C1 => n31, C2 => n696, A 
                           => n697, ZN => n682);
   U406 : AOI22_X1 port map( A1 => REGISTERS_29_19_port, A2 => n34, B1 => 
                           REGISTERS_28_19_port, B2 => n35, ZN => n697);
   U407 : NOR4_X1 port map( A1 => n698, A2 => n699, A3 => n700, A4 => n701, ZN 
                           => n680);
   U409 : AOI22_X1 port map( A1 => REGISTERS_3_19_port, A2 => n45, B1 => 
                           REGISTERS_2_19_port, B2 => n46, ZN => n704);
   U410 : OAI221_X1 port map( B1 => n47, B2 => n705, C1 => n49, C2 => n706, A 
                           => n707, ZN => n700);
   U411 : AOI22_X1 port map( A1 => REGISTERS_7_19_port, A2 => n52, B1 => 
                           REGISTERS_6_19_port, B2 => n53, ZN => n707);
   U412 : OAI221_X1 port map( B1 => n54, B2 => n708, C1 => n56, C2 => n709, A 
                           => n710, ZN => n699);
   U413 : AOI22_X1 port map( A1 => REGISTERS_11_19_port, A2 => n59, B1 => 
                           REGISTERS_10_19_port, B2 => n60, ZN => n710);
   U414 : OAI221_X1 port map( B1 => n61, B2 => n711, C1 => n63, C2 => n712, A 
                           => n713, ZN => n698);
   U415 : AOI22_X1 port map( A1 => REGISTERS_15_19_port, A2 => n66, B1 => 
                           REGISTERS_14_19_port, B2 => n67, ZN => n713);
   U416 : NAND2_X1 port map( A1 => n714, A2 => n715, ZN => N4355);
   U417 : NOR4_X1 port map( A1 => n716, A2 => n717, A3 => n718, A4 => n719, ZN 
                           => n715);
   U418 : OAI221_X1 port map( B1 => n8, B2 => n720, C1 => n10, C2 => n721, A =>
                           n722, ZN => n719);
   U419 : AOI22_X1 port map( A1 => REGISTERS_19_20_port, A2 => n13, B1 => 
                           REGISTERS_18_20_port, B2 => n14, ZN => n722);
   U420 : OAI221_X1 port map( B1 => n15, B2 => n723, C1 => n17, C2 => n724, A 
                           => n725, ZN => n718);
   U421 : AOI22_X1 port map( A1 => REGISTERS_23_20_port, A2 => n20, B1 => 
                           REGISTERS_22_20_port, B2 => n21, ZN => n725);
   U422 : OAI221_X1 port map( B1 => n22, B2 => n726, C1 => n24, C2 => n727, A 
                           => n728, ZN => n717);
   U423 : AOI22_X1 port map( A1 => REGISTERS_27_20_port, A2 => n27, B1 => 
                           REGISTERS_26_20_port, B2 => n28, ZN => n728);
   U424 : OAI221_X1 port map( B1 => n29, B2 => n729, C1 => n31, C2 => n730, A 
                           => n731, ZN => n716);
   U425 : AOI22_X1 port map( A1 => REGISTERS_29_20_port, A2 => n34, B1 => 
                           REGISTERS_28_20_port, B2 => n35, ZN => n731);
   U426 : NOR4_X1 port map( A1 => n732, A2 => n733, A3 => n734, A4 => n735, ZN 
                           => n714);
   U428 : AOI22_X1 port map( A1 => REGISTERS_3_20_port, A2 => n45, B1 => 
                           REGISTERS_2_20_port, B2 => n46, ZN => n738);
   U429 : OAI221_X1 port map( B1 => n47, B2 => n739, C1 => n49, C2 => n740, A 
                           => n741, ZN => n734);
   U430 : AOI22_X1 port map( A1 => REGISTERS_7_20_port, A2 => n52, B1 => 
                           REGISTERS_6_20_port, B2 => n53, ZN => n741);
   U431 : OAI221_X1 port map( B1 => n54, B2 => n742, C1 => n56, C2 => n743, A 
                           => n744, ZN => n733);
   U432 : AOI22_X1 port map( A1 => REGISTERS_11_20_port, A2 => n59, B1 => 
                           REGISTERS_10_20_port, B2 => n60, ZN => n744);
   U433 : OAI221_X1 port map( B1 => n61, B2 => n745, C1 => n63, C2 => n746, A 
                           => n747, ZN => n732);
   U434 : AOI22_X1 port map( A1 => REGISTERS_15_20_port, A2 => n66, B1 => 
                           REGISTERS_14_20_port, B2 => n67, ZN => n747);
   U435 : NAND2_X1 port map( A1 => n748, A2 => n749, ZN => N4354);
   U436 : NOR4_X1 port map( A1 => n750, A2 => n751, A3 => n752, A4 => n753, ZN 
                           => n749);
   U437 : OAI221_X1 port map( B1 => n8, B2 => n754, C1 => n10, C2 => n755, A =>
                           n756, ZN => n753);
   U438 : AOI22_X1 port map( A1 => REGISTERS_19_21_port, A2 => n13, B1 => 
                           REGISTERS_18_21_port, B2 => n14, ZN => n756);
   U439 : OAI221_X1 port map( B1 => n15, B2 => n757, C1 => n17, C2 => n758, A 
                           => n759, ZN => n752);
   U440 : AOI22_X1 port map( A1 => REGISTERS_23_21_port, A2 => n20, B1 => 
                           REGISTERS_22_21_port, B2 => n21, ZN => n759);
   U441 : OAI221_X1 port map( B1 => n22, B2 => n760, C1 => n24, C2 => n761, A 
                           => n762, ZN => n751);
   U442 : AOI22_X1 port map( A1 => REGISTERS_27_21_port, A2 => n27, B1 => 
                           REGISTERS_26_21_port, B2 => n28, ZN => n762);
   U443 : OAI221_X1 port map( B1 => n29, B2 => n763, C1 => n31, C2 => n764, A 
                           => n765, ZN => n750);
   U444 : AOI22_X1 port map( A1 => REGISTERS_29_21_port, A2 => n34, B1 => 
                           REGISTERS_28_21_port, B2 => n35, ZN => n765);
   U445 : NOR4_X1 port map( A1 => n766, A2 => n767, A3 => n768, A4 => n769, ZN 
                           => n748);
   U447 : AOI22_X1 port map( A1 => REGISTERS_3_21_port, A2 => n45, B1 => 
                           REGISTERS_2_21_port, B2 => n46, ZN => n772);
   U448 : OAI221_X1 port map( B1 => n47, B2 => n773, C1 => n49, C2 => n774, A 
                           => n775, ZN => n768);
   U449 : AOI22_X1 port map( A1 => REGISTERS_7_21_port, A2 => n52, B1 => 
                           REGISTERS_6_21_port, B2 => n53, ZN => n775);
   U450 : OAI221_X1 port map( B1 => n54, B2 => n776, C1 => n56, C2 => n777, A 
                           => n778, ZN => n767);
   U451 : AOI22_X1 port map( A1 => REGISTERS_11_21_port, A2 => n59, B1 => 
                           REGISTERS_10_21_port, B2 => n60, ZN => n778);
   U452 : OAI221_X1 port map( B1 => n61, B2 => n779, C1 => n63, C2 => n780, A 
                           => n781, ZN => n766);
   U453 : AOI22_X1 port map( A1 => REGISTERS_15_21_port, A2 => n66, B1 => 
                           REGISTERS_14_21_port, B2 => n67, ZN => n781);
   U454 : NAND2_X1 port map( A1 => n782, A2 => n783, ZN => N4353);
   U455 : NOR4_X1 port map( A1 => n784, A2 => n785, A3 => n786, A4 => n787, ZN 
                           => n783);
   U456 : OAI221_X1 port map( B1 => n8, B2 => n788, C1 => n10, C2 => n789, A =>
                           n790, ZN => n787);
   U457 : AOI22_X1 port map( A1 => REGISTERS_19_22_port, A2 => n13, B1 => 
                           REGISTERS_18_22_port, B2 => n14, ZN => n790);
   U458 : OAI221_X1 port map( B1 => n15, B2 => n791, C1 => n17, C2 => n792, A 
                           => n793, ZN => n786);
   U459 : AOI22_X1 port map( A1 => REGISTERS_23_22_port, A2 => n20, B1 => 
                           REGISTERS_22_22_port, B2 => n21, ZN => n793);
   U460 : OAI221_X1 port map( B1 => n22, B2 => n794, C1 => n24, C2 => n795, A 
                           => n796, ZN => n785);
   U461 : AOI22_X1 port map( A1 => REGISTERS_27_22_port, A2 => n27, B1 => 
                           REGISTERS_26_22_port, B2 => n28, ZN => n796);
   U462 : OAI221_X1 port map( B1 => n29, B2 => n797, C1 => n31, C2 => n798, A 
                           => n799, ZN => n784);
   U463 : AOI22_X1 port map( A1 => REGISTERS_29_22_port, A2 => n34, B1 => 
                           REGISTERS_28_22_port, B2 => n35, ZN => n799);
   U464 : NOR4_X1 port map( A1 => n800, A2 => n801, A3 => n802, A4 => n803, ZN 
                           => n782);
   U466 : AOI22_X1 port map( A1 => REGISTERS_3_22_port, A2 => n45, B1 => 
                           REGISTERS_2_22_port, B2 => n46, ZN => n806);
   U467 : OAI221_X1 port map( B1 => n47, B2 => n807, C1 => n49, C2 => n808, A 
                           => n809, ZN => n802);
   U468 : AOI22_X1 port map( A1 => REGISTERS_7_22_port, A2 => n52, B1 => 
                           REGISTERS_6_22_port, B2 => n53, ZN => n809);
   U469 : OAI221_X1 port map( B1 => n54, B2 => n810, C1 => n56, C2 => n811, A 
                           => n812, ZN => n801);
   U470 : AOI22_X1 port map( A1 => REGISTERS_11_22_port, A2 => n59, B1 => 
                           REGISTERS_10_22_port, B2 => n60, ZN => n812);
   U471 : OAI221_X1 port map( B1 => n61, B2 => n813, C1 => n63, C2 => n814, A 
                           => n815, ZN => n800);
   U472 : AOI22_X1 port map( A1 => REGISTERS_15_22_port, A2 => n66, B1 => 
                           REGISTERS_14_22_port, B2 => n67, ZN => n815);
   U473 : NAND2_X1 port map( A1 => n816, A2 => n817, ZN => N4352);
   U474 : NOR4_X1 port map( A1 => n818, A2 => n819, A3 => n820, A4 => n821, ZN 
                           => n817);
   U475 : OAI221_X1 port map( B1 => n8, B2 => n822, C1 => n10, C2 => n823, A =>
                           n824, ZN => n821);
   U476 : AOI22_X1 port map( A1 => REGISTERS_19_23_port, A2 => n13, B1 => 
                           REGISTERS_18_23_port, B2 => n14, ZN => n824);
   U477 : OAI221_X1 port map( B1 => n15, B2 => n825, C1 => n17, C2 => n826, A 
                           => n827, ZN => n820);
   U478 : AOI22_X1 port map( A1 => REGISTERS_23_23_port, A2 => n20, B1 => 
                           REGISTERS_22_23_port, B2 => n21, ZN => n827);
   U479 : OAI221_X1 port map( B1 => n22, B2 => n828, C1 => n24, C2 => n829, A 
                           => n830, ZN => n819);
   U480 : AOI22_X1 port map( A1 => REGISTERS_27_23_port, A2 => n27, B1 => 
                           REGISTERS_26_23_port, B2 => n28, ZN => n830);
   U481 : OAI221_X1 port map( B1 => n29, B2 => n831, C1 => n31, C2 => n832, A 
                           => n833, ZN => n818);
   U482 : AOI22_X1 port map( A1 => REGISTERS_29_23_port, A2 => n34, B1 => 
                           REGISTERS_28_23_port, B2 => n35, ZN => n833);
   U483 : NOR4_X1 port map( A1 => n834, A2 => n835, A3 => n836, A4 => n837, ZN 
                           => n816);
   U485 : AOI22_X1 port map( A1 => REGISTERS_3_23_port, A2 => n45, B1 => 
                           REGISTERS_2_23_port, B2 => n46, ZN => n840);
   U486 : OAI221_X1 port map( B1 => n47, B2 => n841, C1 => n49, C2 => n842, A 
                           => n843, ZN => n836);
   U487 : AOI22_X1 port map( A1 => REGISTERS_7_23_port, A2 => n52, B1 => 
                           REGISTERS_6_23_port, B2 => n53, ZN => n843);
   U488 : OAI221_X1 port map( B1 => n54, B2 => n844, C1 => n56, C2 => n845, A 
                           => n846, ZN => n835);
   U489 : AOI22_X1 port map( A1 => REGISTERS_11_23_port, A2 => n59, B1 => 
                           REGISTERS_10_23_port, B2 => n60, ZN => n846);
   U490 : OAI221_X1 port map( B1 => n61, B2 => n847, C1 => n63, C2 => n848, A 
                           => n849, ZN => n834);
   U491 : AOI22_X1 port map( A1 => REGISTERS_15_23_port, A2 => n66, B1 => 
                           REGISTERS_14_23_port, B2 => n67, ZN => n849);
   U492 : NAND2_X1 port map( A1 => n850, A2 => n851, ZN => N4351);
   U493 : NOR4_X1 port map( A1 => n852, A2 => n853, A3 => n854, A4 => n855, ZN 
                           => n851);
   U494 : OAI221_X1 port map( B1 => n8, B2 => n856, C1 => n10, C2 => n857, A =>
                           n858, ZN => n855);
   U495 : AOI22_X1 port map( A1 => REGISTERS_19_24_port, A2 => n13, B1 => 
                           REGISTERS_18_24_port, B2 => n14, ZN => n858);
   U496 : OAI221_X1 port map( B1 => n15, B2 => n859, C1 => n17, C2 => n860, A 
                           => n861, ZN => n854);
   U497 : AOI22_X1 port map( A1 => REGISTERS_23_24_port, A2 => n20, B1 => 
                           REGISTERS_22_24_port, B2 => n21, ZN => n861);
   U498 : OAI221_X1 port map( B1 => n22, B2 => n862, C1 => n24, C2 => n863, A 
                           => n864, ZN => n853);
   U499 : AOI22_X1 port map( A1 => REGISTERS_27_24_port, A2 => n27, B1 => 
                           REGISTERS_26_24_port, B2 => n28, ZN => n864);
   U500 : OAI221_X1 port map( B1 => n29, B2 => n865, C1 => n31, C2 => n866, A 
                           => n867, ZN => n852);
   U501 : AOI22_X1 port map( A1 => REGISTERS_29_24_port, A2 => n34, B1 => 
                           REGISTERS_28_24_port, B2 => n35, ZN => n867);
   U502 : NOR4_X1 port map( A1 => n868, A2 => n869, A3 => n870, A4 => n871, ZN 
                           => n850);
   U504 : AOI22_X1 port map( A1 => REGISTERS_3_24_port, A2 => n45, B1 => 
                           REGISTERS_2_24_port, B2 => n46, ZN => n874);
   U505 : OAI221_X1 port map( B1 => n47, B2 => n875, C1 => n49, C2 => n876, A 
                           => n877, ZN => n870);
   U506 : AOI22_X1 port map( A1 => REGISTERS_7_24_port, A2 => n52, B1 => 
                           REGISTERS_6_24_port, B2 => n53, ZN => n877);
   U507 : OAI221_X1 port map( B1 => n54, B2 => n878, C1 => n56, C2 => n879, A 
                           => n880, ZN => n869);
   U508 : AOI22_X1 port map( A1 => REGISTERS_11_24_port, A2 => n59, B1 => 
                           REGISTERS_10_24_port, B2 => n60, ZN => n880);
   U509 : OAI221_X1 port map( B1 => n61, B2 => n881, C1 => n63, C2 => n882, A 
                           => n883, ZN => n868);
   U510 : AOI22_X1 port map( A1 => REGISTERS_15_24_port, A2 => n66, B1 => 
                           REGISTERS_14_24_port, B2 => n67, ZN => n883);
   U511 : NAND2_X1 port map( A1 => n884, A2 => n885, ZN => N4350);
   U512 : NOR4_X1 port map( A1 => n886, A2 => n887, A3 => n888, A4 => n889, ZN 
                           => n885);
   U513 : OAI221_X1 port map( B1 => n8, B2 => n890, C1 => n10, C2 => n891, A =>
                           n892, ZN => n889);
   U514 : AOI22_X1 port map( A1 => REGISTERS_19_25_port, A2 => n13, B1 => 
                           REGISTERS_18_25_port, B2 => n14, ZN => n892);
   U515 : OAI221_X1 port map( B1 => n15, B2 => n893, C1 => n17, C2 => n894, A 
                           => n895, ZN => n888);
   U516 : AOI22_X1 port map( A1 => REGISTERS_23_25_port, A2 => n20, B1 => 
                           REGISTERS_22_25_port, B2 => n21, ZN => n895);
   U517 : OAI221_X1 port map( B1 => n22, B2 => n896, C1 => n24, C2 => n897, A 
                           => n898, ZN => n887);
   U518 : AOI22_X1 port map( A1 => REGISTERS_27_25_port, A2 => n27, B1 => 
                           REGISTERS_26_25_port, B2 => n28, ZN => n898);
   U519 : OAI221_X1 port map( B1 => n29, B2 => n899, C1 => n31, C2 => n900, A 
                           => n901, ZN => n886);
   U520 : AOI22_X1 port map( A1 => REGISTERS_29_25_port, A2 => n34, B1 => 
                           REGISTERS_28_25_port, B2 => n35, ZN => n901);
   U521 : NOR4_X1 port map( A1 => n902, A2 => n903, A3 => n904, A4 => n905, ZN 
                           => n884);
   U523 : AOI22_X1 port map( A1 => REGISTERS_3_25_port, A2 => n45, B1 => 
                           REGISTERS_2_25_port, B2 => n46, ZN => n908);
   U524 : OAI221_X1 port map( B1 => n47, B2 => n909, C1 => n49, C2 => n910, A 
                           => n911, ZN => n904);
   U525 : AOI22_X1 port map( A1 => REGISTERS_7_25_port, A2 => n52, B1 => 
                           REGISTERS_6_25_port, B2 => n53, ZN => n911);
   U526 : OAI221_X1 port map( B1 => n54, B2 => n912, C1 => n56, C2 => n913, A 
                           => n914, ZN => n903);
   U527 : AOI22_X1 port map( A1 => REGISTERS_11_25_port, A2 => n59, B1 => 
                           REGISTERS_10_25_port, B2 => n60, ZN => n914);
   U528 : OAI221_X1 port map( B1 => n61, B2 => n915, C1 => n63, C2 => n916, A 
                           => n917, ZN => n902);
   U529 : AOI22_X1 port map( A1 => REGISTERS_15_25_port, A2 => n66, B1 => 
                           REGISTERS_14_25_port, B2 => n67, ZN => n917);
   U530 : NAND2_X1 port map( A1 => n918, A2 => n919, ZN => N4349);
   U531 : NOR4_X1 port map( A1 => n920, A2 => n921, A3 => n922, A4 => n923, ZN 
                           => n919);
   U532 : OAI221_X1 port map( B1 => n8, B2 => n924, C1 => n10, C2 => n925, A =>
                           n926, ZN => n923);
   U533 : AOI22_X1 port map( A1 => REGISTERS_19_26_port, A2 => n13, B1 => 
                           REGISTERS_18_26_port, B2 => n14, ZN => n926);
   U534 : OAI221_X1 port map( B1 => n15, B2 => n927, C1 => n17, C2 => n928, A 
                           => n929, ZN => n922);
   U535 : AOI22_X1 port map( A1 => REGISTERS_23_26_port, A2 => n20, B1 => 
                           REGISTERS_22_26_port, B2 => n21, ZN => n929);
   U536 : OAI221_X1 port map( B1 => n22, B2 => n930, C1 => n24, C2 => n931, A 
                           => n932, ZN => n921);
   U537 : AOI22_X1 port map( A1 => REGISTERS_27_26_port, A2 => n27, B1 => 
                           REGISTERS_26_26_port, B2 => n28, ZN => n932);
   U538 : OAI221_X1 port map( B1 => n29, B2 => n933, C1 => n31, C2 => n934, A 
                           => n935, ZN => n920);
   U539 : AOI22_X1 port map( A1 => REGISTERS_29_26_port, A2 => n34, B1 => 
                           REGISTERS_28_26_port, B2 => n35, ZN => n935);
   U540 : NOR4_X1 port map( A1 => n936, A2 => n937, A3 => n938, A4 => n939, ZN 
                           => n918);
   U542 : AOI22_X1 port map( A1 => REGISTERS_3_26_port, A2 => n45, B1 => 
                           REGISTERS_2_26_port, B2 => n46, ZN => n942);
   U543 : OAI221_X1 port map( B1 => n47, B2 => n943, C1 => n49, C2 => n944, A 
                           => n945, ZN => n938);
   U544 : AOI22_X1 port map( A1 => REGISTERS_7_26_port, A2 => n52, B1 => 
                           REGISTERS_6_26_port, B2 => n53, ZN => n945);
   U545 : OAI221_X1 port map( B1 => n54, B2 => n946, C1 => n56, C2 => n947, A 
                           => n948, ZN => n937);
   U546 : AOI22_X1 port map( A1 => REGISTERS_11_26_port, A2 => n59, B1 => 
                           REGISTERS_10_26_port, B2 => n60, ZN => n948);
   U547 : OAI221_X1 port map( B1 => n61, B2 => n949, C1 => n63, C2 => n950, A 
                           => n951, ZN => n936);
   U548 : AOI22_X1 port map( A1 => REGISTERS_15_26_port, A2 => n66, B1 => 
                           REGISTERS_14_26_port, B2 => n67, ZN => n951);
   U549 : NAND2_X1 port map( A1 => n952, A2 => n953, ZN => N4348);
   U550 : NOR4_X1 port map( A1 => n954, A2 => n955, A3 => n956, A4 => n957, ZN 
                           => n953);
   U551 : OAI221_X1 port map( B1 => n8, B2 => n958, C1 => n10, C2 => n959, A =>
                           n960, ZN => n957);
   U552 : AOI22_X1 port map( A1 => REGISTERS_19_27_port, A2 => n13, B1 => 
                           REGISTERS_18_27_port, B2 => n14, ZN => n960);
   U553 : OAI221_X1 port map( B1 => n15, B2 => n961, C1 => n17, C2 => n962, A 
                           => n963, ZN => n956);
   U554 : AOI22_X1 port map( A1 => REGISTERS_23_27_port, A2 => n20, B1 => 
                           REGISTERS_22_27_port, B2 => n21, ZN => n963);
   U555 : OAI221_X1 port map( B1 => n22, B2 => n964, C1 => n24, C2 => n965, A 
                           => n966, ZN => n955);
   U556 : AOI22_X1 port map( A1 => REGISTERS_27_27_port, A2 => n27, B1 => 
                           REGISTERS_26_27_port, B2 => n28, ZN => n966);
   U557 : OAI221_X1 port map( B1 => n29, B2 => n967, C1 => n31, C2 => n968, A 
                           => n969, ZN => n954);
   U558 : AOI22_X1 port map( A1 => REGISTERS_29_27_port, A2 => n34, B1 => 
                           REGISTERS_28_27_port, B2 => n35, ZN => n969);
   U559 : NOR4_X1 port map( A1 => n970, A2 => n971, A3 => n972, A4 => n973, ZN 
                           => n952);
   U561 : AOI22_X1 port map( A1 => REGISTERS_3_27_port, A2 => n45, B1 => 
                           REGISTERS_2_27_port, B2 => n46, ZN => n976);
   U562 : OAI221_X1 port map( B1 => n47, B2 => n977, C1 => n49, C2 => n978, A 
                           => n979, ZN => n972);
   U563 : AOI22_X1 port map( A1 => REGISTERS_7_27_port, A2 => n52, B1 => 
                           REGISTERS_6_27_port, B2 => n53, ZN => n979);
   U564 : OAI221_X1 port map( B1 => n54, B2 => n980, C1 => n56, C2 => n981, A 
                           => n982, ZN => n971);
   U565 : AOI22_X1 port map( A1 => REGISTERS_11_27_port, A2 => n59, B1 => 
                           REGISTERS_10_27_port, B2 => n60, ZN => n982);
   U566 : OAI221_X1 port map( B1 => n61, B2 => n983, C1 => n63, C2 => n984, A 
                           => n985, ZN => n970);
   U567 : AOI22_X1 port map( A1 => REGISTERS_15_27_port, A2 => n66, B1 => 
                           REGISTERS_14_27_port, B2 => n67, ZN => n985);
   U568 : NAND2_X1 port map( A1 => n986, A2 => n987, ZN => N4347);
   U569 : NOR4_X1 port map( A1 => n988, A2 => n989, A3 => n990, A4 => n991, ZN 
                           => n987);
   U570 : OAI221_X1 port map( B1 => n8, B2 => n992, C1 => n10, C2 => n993, A =>
                           n994, ZN => n991);
   U571 : AOI22_X1 port map( A1 => REGISTERS_19_28_port, A2 => n13, B1 => 
                           REGISTERS_18_28_port, B2 => n14, ZN => n994);
   U572 : OAI221_X1 port map( B1 => n15, B2 => n995, C1 => n17, C2 => n996, A 
                           => n997, ZN => n990);
   U573 : AOI22_X1 port map( A1 => REGISTERS_23_28_port, A2 => n20, B1 => 
                           REGISTERS_22_28_port, B2 => n21, ZN => n997);
   U574 : OAI221_X1 port map( B1 => n22, B2 => n998, C1 => n24, C2 => n999, A 
                           => n1000, ZN => n989);
   U575 : AOI22_X1 port map( A1 => REGISTERS_27_28_port, A2 => n27, B1 => 
                           REGISTERS_26_28_port, B2 => n28, ZN => n1000);
   U576 : OAI221_X1 port map( B1 => n29, B2 => n1001, C1 => n31, C2 => n1002, A
                           => n1003, ZN => n988);
   U577 : AOI22_X1 port map( A1 => REGISTERS_29_28_port, A2 => n34, B1 => 
                           REGISTERS_28_28_port, B2 => n35, ZN => n1003);
   U578 : NOR4_X1 port map( A1 => n1004, A2 => n1005, A3 => n1006, A4 => n1007,
                           ZN => n986);
   U580 : AOI22_X1 port map( A1 => REGISTERS_3_28_port, A2 => n45, B1 => 
                           REGISTERS_2_28_port, B2 => n46, ZN => n1010);
   U581 : OAI221_X1 port map( B1 => n47, B2 => n1011, C1 => n49, C2 => n1012, A
                           => n1013, ZN => n1006);
   U582 : AOI22_X1 port map( A1 => REGISTERS_7_28_port, A2 => n52, B1 => 
                           REGISTERS_6_28_port, B2 => n53, ZN => n1013);
   U583 : OAI221_X1 port map( B1 => n54, B2 => n1014, C1 => n56, C2 => n1015, A
                           => n1016, ZN => n1005);
   U584 : AOI22_X1 port map( A1 => REGISTERS_11_28_port, A2 => n59, B1 => 
                           REGISTERS_10_28_port, B2 => n60, ZN => n1016);
   U585 : OAI221_X1 port map( B1 => n61, B2 => n1017, C1 => n63, C2 => n1018, A
                           => n1019, ZN => n1004);
   U586 : AOI22_X1 port map( A1 => REGISTERS_15_28_port, A2 => n66, B1 => 
                           REGISTERS_14_28_port, B2 => n67, ZN => n1019);
   U587 : NAND2_X1 port map( A1 => n1020, A2 => n1021, ZN => N4346);
   U588 : NOR4_X1 port map( A1 => n1022, A2 => n1023, A3 => n1024, A4 => n1025,
                           ZN => n1021);
   U589 : OAI221_X1 port map( B1 => n8, B2 => n1026, C1 => n10, C2 => n1027, A 
                           => n1028, ZN => n1025);
   U590 : AOI22_X1 port map( A1 => REGISTERS_19_29_port, A2 => n13, B1 => 
                           REGISTERS_18_29_port, B2 => n14, ZN => n1028);
   U591 : OAI221_X1 port map( B1 => n15, B2 => n1029, C1 => n17, C2 => n1030, A
                           => n1031, ZN => n1024);
   U592 : AOI22_X1 port map( A1 => REGISTERS_23_29_port, A2 => n20, B1 => 
                           REGISTERS_22_29_port, B2 => n21, ZN => n1031);
   U593 : OAI221_X1 port map( B1 => n22, B2 => n1032, C1 => n24, C2 => n1033, A
                           => n1034, ZN => n1023);
   U594 : AOI22_X1 port map( A1 => REGISTERS_27_29_port, A2 => n27, B1 => 
                           REGISTERS_26_29_port, B2 => n28, ZN => n1034);
   U595 : OAI221_X1 port map( B1 => n29, B2 => n1035, C1 => n31, C2 => n1036, A
                           => n1037, ZN => n1022);
   U596 : AOI22_X1 port map( A1 => REGISTERS_29_29_port, A2 => n34, B1 => 
                           REGISTERS_28_29_port, B2 => n35, ZN => n1037);
   U597 : NOR4_X1 port map( A1 => n1038, A2 => n1039, A3 => n1040, A4 => n1041,
                           ZN => n1020);
   U599 : AOI22_X1 port map( A1 => REGISTERS_3_29_port, A2 => n45, B1 => 
                           REGISTERS_2_29_port, B2 => n46, ZN => n1044);
   U600 : OAI221_X1 port map( B1 => n47, B2 => n1045, C1 => n49, C2 => n1046, A
                           => n1047, ZN => n1040);
   U601 : AOI22_X1 port map( A1 => REGISTERS_7_29_port, A2 => n52, B1 => 
                           REGISTERS_6_29_port, B2 => n53, ZN => n1047);
   U602 : OAI221_X1 port map( B1 => n54, B2 => n1048, C1 => n56, C2 => n1049, A
                           => n1050, ZN => n1039);
   U603 : AOI22_X1 port map( A1 => REGISTERS_11_29_port, A2 => n59, B1 => 
                           REGISTERS_10_29_port, B2 => n60, ZN => n1050);
   U604 : OAI221_X1 port map( B1 => n61, B2 => n1051, C1 => n63, C2 => n1052, A
                           => n1053, ZN => n1038);
   U605 : AOI22_X1 port map( A1 => REGISTERS_15_29_port, A2 => n66, B1 => 
                           REGISTERS_14_29_port, B2 => n67, ZN => n1053);
   U606 : NAND2_X1 port map( A1 => n1054, A2 => n1055, ZN => N4345);
   U607 : NOR4_X1 port map( A1 => n1056, A2 => n1057, A3 => n1058, A4 => n1059,
                           ZN => n1055);
   U608 : OAI221_X1 port map( B1 => n8, B2 => n1060, C1 => n10, C2 => n1061, A 
                           => n1062, ZN => n1059);
   U609 : AOI22_X1 port map( A1 => REGISTERS_19_30_port, A2 => n13, B1 => 
                           REGISTERS_18_30_port, B2 => n14, ZN => n1062);
   U610 : OAI221_X1 port map( B1 => n15, B2 => n1063, C1 => n17, C2 => n1064, A
                           => n1065, ZN => n1058);
   U611 : AOI22_X1 port map( A1 => REGISTERS_23_30_port, A2 => n20, B1 => 
                           REGISTERS_22_30_port, B2 => n21, ZN => n1065);
   U612 : OAI221_X1 port map( B1 => n22, B2 => n1066, C1 => n24, C2 => n1067, A
                           => n1068, ZN => n1057);
   U613 : AOI22_X1 port map( A1 => REGISTERS_27_30_port, A2 => n27, B1 => 
                           REGISTERS_26_30_port, B2 => n28, ZN => n1068);
   U614 : OAI221_X1 port map( B1 => n29, B2 => n1069, C1 => n31, C2 => n1070, A
                           => n1071, ZN => n1056);
   U615 : AOI22_X1 port map( A1 => REGISTERS_29_30_port, A2 => n34, B1 => 
                           REGISTERS_28_30_port, B2 => n35, ZN => n1071);
   U616 : NOR4_X1 port map( A1 => n1072, A2 => n1073, A3 => n1074, A4 => n1075,
                           ZN => n1054);
   U618 : AOI22_X1 port map( A1 => REGISTERS_3_30_port, A2 => n45, B1 => 
                           REGISTERS_2_30_port, B2 => n46, ZN => n1078);
   U619 : OAI221_X1 port map( B1 => n47, B2 => n1079, C1 => n49, C2 => n1080, A
                           => n1081, ZN => n1074);
   U620 : AOI22_X1 port map( A1 => REGISTERS_7_30_port, A2 => n52, B1 => 
                           REGISTERS_6_30_port, B2 => n53, ZN => n1081);
   U621 : OAI221_X1 port map( B1 => n54, B2 => n1082, C1 => n56, C2 => n1083, A
                           => n1084, ZN => n1073);
   U622 : AOI22_X1 port map( A1 => REGISTERS_11_30_port, A2 => n59, B1 => 
                           REGISTERS_10_30_port, B2 => n60, ZN => n1084);
   U623 : OAI221_X1 port map( B1 => n61, B2 => n1085, C1 => n63, C2 => n1086, A
                           => n1087, ZN => n1072);
   U624 : AOI22_X1 port map( A1 => REGISTERS_15_30_port, A2 => n66, B1 => 
                           REGISTERS_14_30_port, B2 => n67, ZN => n1087);
   U625 : NAND2_X1 port map( A1 => n1088, A2 => n1089, ZN => N4344);
   U626 : NOR4_X1 port map( A1 => n1090, A2 => n1091, A3 => n1092, A4 => n1093,
                           ZN => n1089);
   U627 : OAI221_X1 port map( B1 => n8, B2 => n1094, C1 => n10, C2 => n1095, A 
                           => n1096, ZN => n1093);
   U628 : AOI22_X1 port map( A1 => REGISTERS_19_31_port, A2 => n13, B1 => 
                           REGISTERS_18_31_port, B2 => n14, ZN => n1096);
   U633 : OAI221_X1 port map( B1 => n15, B2 => n1101, C1 => n17, C2 => n1102, A
                           => n1103, ZN => n1092);
   U634 : AOI22_X1 port map( A1 => REGISTERS_23_31_port, A2 => n20, B1 => 
                           REGISTERS_22_31_port, B2 => n21, ZN => n1103);
   U638 : AND2_X1 port map( A1 => n1106, A2 => n1107, ZN => n1097);
   U640 : AND2_X1 port map( A1 => n1106, A2 => ADD_RD2(0), ZN => n1099);
   U641 : AND2_X1 port map( A1 => ADD_RD2(4), A2 => n1108, ZN => n1106);
   U642 : OAI221_X1 port map( B1 => n22, B2 => n1109, C1 => n24, C2 => n1110, A
                           => n1111, ZN => n1091);
   U643 : AOI22_X1 port map( A1 => REGISTERS_27_31_port, A2 => n27, B1 => 
                           REGISTERS_26_31_port, B2 => n28, ZN => n1111);
   U648 : OAI221_X1 port map( B1 => n29, B2 => n1114, C1 => n31, C2 => n1115, A
                           => n1116, ZN => n1090);
   U649 : AOI22_X1 port map( A1 => REGISTERS_29_31_port, A2 => n34, B1 => 
                           REGISTERS_28_31_port, B2 => n35, ZN => n1116);
   U653 : AND2_X1 port map( A1 => n1117, A2 => n1107, ZN => n1112);
   U655 : AND2_X1 port map( A1 => ADD_RD2(0), A2 => n1117, ZN => n1113);
   U656 : AND2_X1 port map( A1 => ADD_RD2(4), A2 => ADD_RD2(3), ZN => n1117);
   U657 : NOR4_X1 port map( A1 => n1118, A2 => n1119, A3 => n1120, A4 => n1121,
                           ZN => n1088);
   U659 : AOI22_X1 port map( A1 => REGISTERS_3_31_port, A2 => n45, B1 => 
                           REGISTERS_2_31_port, B2 => n46, ZN => n1124);
   U664 : OAI221_X1 port map( B1 => n47, B2 => n1127, C1 => n49, C2 => n1128, A
                           => n1129, ZN => n1120);
   U665 : AOI22_X1 port map( A1 => REGISTERS_7_31_port, A2 => n52, B1 => 
                           REGISTERS_6_31_port, B2 => n53, ZN => n1129);
   U669 : AND2_X1 port map( A1 => n1130, A2 => n1107, ZN => n1125);
   U671 : AND2_X1 port map( A1 => n1130, A2 => ADD_RD2(0), ZN => n1126);
   U672 : NOR2_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), ZN => n1130);
   U673 : OAI221_X1 port map( B1 => n54, B2 => n1131, C1 => n56, C2 => n1132, A
                           => n1133, ZN => n1119);
   U674 : AOI22_X1 port map( A1 => REGISTERS_11_31_port, A2 => n59, B1 => 
                           REGISTERS_10_31_port, B2 => n60, ZN => n1133);
   U677 : NOR2_X1 port map( A1 => n1136, A2 => ADD_RD2(2), ZN => n1098);
   U680 : NOR2_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), ZN => n1100);
   U681 : OAI221_X1 port map( B1 => n61, B2 => n1137, C1 => n63, C2 => n1138, A
                           => n1139, ZN => n1118);
   U682 : AOI22_X1 port map( A1 => REGISTERS_15_31_port, A2 => n66, B1 => 
                           REGISTERS_14_31_port, B2 => n67, ZN => n1139);
   U685 : NOR2_X1 port map( A1 => n1140, A2 => n1136, ZN => n1104);
   U686 : INV_X1 port map( A => ADD_RD2(1), ZN => n1136);
   U688 : AND2_X1 port map( A1 => n1141, A2 => n1107, ZN => n1134);
   U689 : INV_X1 port map( A => ADD_RD2(0), ZN => n1107);
   U692 : INV_X1 port map( A => ADD_RD2(2), ZN => n1140);
   U693 : AND2_X1 port map( A1 => n1141, A2 => ADD_RD2(0), ZN => n1135);
   U694 : NOR2_X1 port map( A1 => n1108, A2 => ADD_RD2(4), ZN => n1141);
   U695 : INV_X1 port map( A => ADD_RD2(3), ZN => n1108);
   U696 : AND2_X1 port map( A1 => RD1, A2 => ENABLE, ZN => N4278);
   U697 : NAND2_X1 port map( A1 => n1142, A2 => n1143, ZN => N4246);
   U698 : NOR4_X1 port map( A1 => n1144, A2 => n1145, A3 => n1146, A4 => n1147,
                           ZN => n1143);
   U699 : OAI221_X1 port map( B1 => n9, B2 => n1148, C1 => n11, C2 => n1149, A 
                           => n1150, ZN => n1147);
   U700 : AOI22_X1 port map( A1 => n1151, A2 => REGISTERS_19_0_port, B1 => 
                           n1152, B2 => REGISTERS_18_0_port, ZN => n1150);
   U701 : INV_X1 port map( A => REGISTERS_16_0_port, ZN => n11);
   U702 : INV_X1 port map( A => REGISTERS_17_0_port, ZN => n9);
   U703 : OAI221_X1 port map( B1 => n16, B2 => n1153, C1 => n18, C2 => n1154, A
                           => n1155, ZN => n1146);
   U704 : AOI22_X1 port map( A1 => n1156, A2 => REGISTERS_23_0_port, B1 => 
                           n1157, B2 => REGISTERS_22_0_port, ZN => n1155);
   U705 : INV_X1 port map( A => REGISTERS_20_0_port, ZN => n18);
   U706 : INV_X1 port map( A => REGISTERS_21_0_port, ZN => n16);
   U707 : OAI221_X1 port map( B1 => n23, B2 => n1158, C1 => n25, C2 => n1159, A
                           => n1160, ZN => n1145);
   U708 : AOI22_X1 port map( A1 => n1161, A2 => REGISTERS_27_0_port, B1 => 
                           n1162, B2 => REGISTERS_26_0_port, ZN => n1160);
   U709 : INV_X1 port map( A => REGISTERS_24_0_port, ZN => n25);
   U710 : INV_X1 port map( A => REGISTERS_25_0_port, ZN => n23);
   U711 : OAI221_X1 port map( B1 => n30, B2 => n1163, C1 => n32, C2 => n1164, A
                           => n1165, ZN => n1144);
   U712 : AOI22_X1 port map( A1 => n1166, A2 => REGISTERS_29_0_port, B1 => 
                           n1167, B2 => REGISTERS_28_0_port, ZN => n1165);
   U713 : INV_X1 port map( A => REGISTERS_30_0_port, ZN => n32);
   U714 : INV_X1 port map( A => REGISTERS_31_0_port, ZN => n30);
   U715 : NOR4_X1 port map( A1 => n1168, A2 => n1169, A3 => n1170, A4 => n1171,
                           ZN => n1142);
   U717 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_3_0_port, B1 => n1176
                           , B2 => REGISTERS_2_0_port, ZN => n1174);
   U718 : INV_X1 port map( A => REGISTERS_1_0_port, ZN => n41);
   U719 : OAI221_X1 port map( B1 => n48, B2 => n1177, C1 => n50, C2 => n1178, A
                           => n1179, ZN => n1170);
   U720 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_7_0_port, B1 => n1181
                           , B2 => REGISTERS_6_0_port, ZN => n1179);
   U721 : INV_X1 port map( A => REGISTERS_4_0_port, ZN => n50);
   U722 : INV_X1 port map( A => REGISTERS_5_0_port, ZN => n48);
   U723 : OAI221_X1 port map( B1 => n55, B2 => n1182, C1 => n57, C2 => n1183, A
                           => n1184, ZN => n1169);
   U724 : AOI22_X1 port map( A1 => n1185, A2 => REGISTERS_11_0_port, B1 => 
                           n1186, B2 => REGISTERS_10_0_port, ZN => n1184);
   U725 : INV_X1 port map( A => REGISTERS_8_0_port, ZN => n57);
   U726 : INV_X1 port map( A => REGISTERS_9_0_port, ZN => n55);
   U727 : OAI221_X1 port map( B1 => n62, B2 => n1187, C1 => n64, C2 => n1188, A
                           => n1189, ZN => n1168);
   U728 : AOI22_X1 port map( A1 => n1190, A2 => REGISTERS_15_0_port, B1 => 
                           n1191, B2 => REGISTERS_14_0_port, ZN => n1189);
   U729 : INV_X1 port map( A => REGISTERS_12_0_port, ZN => n64);
   U730 : INV_X1 port map( A => REGISTERS_13_0_port, ZN => n62);
   U731 : NAND2_X1 port map( A1 => n1192, A2 => n1193, ZN => N4245);
   U732 : NOR4_X1 port map( A1 => n1194, A2 => n1195, A3 => n1196, A4 => n1197,
                           ZN => n1193);
   U733 : OAI221_X1 port map( B1 => n74, B2 => n1148, C1 => n75, C2 => n1149, A
                           => n1198, ZN => n1197);
   U734 : AOI22_X1 port map( A1 => n1151, A2 => REGISTERS_19_1_port, B1 => 
                           n1152, B2 => REGISTERS_18_1_port, ZN => n1198);
   U735 : INV_X1 port map( A => REGISTERS_16_1_port, ZN => n75);
   U736 : INV_X1 port map( A => REGISTERS_17_1_port, ZN => n74);
   U737 : OAI221_X1 port map( B1 => n77, B2 => n1153, C1 => n78, C2 => n1154, A
                           => n1199, ZN => n1196);
   U738 : AOI22_X1 port map( A1 => n1156, A2 => REGISTERS_23_1_port, B1 => 
                           n1157, B2 => REGISTERS_22_1_port, ZN => n1199);
   U739 : INV_X1 port map( A => REGISTERS_20_1_port, ZN => n78);
   U740 : INV_X1 port map( A => REGISTERS_21_1_port, ZN => n77);
   U741 : OAI221_X1 port map( B1 => n80, B2 => n1158, C1 => n81, C2 => n1159, A
                           => n1200, ZN => n1195);
   U742 : AOI22_X1 port map( A1 => n1161, A2 => REGISTERS_27_1_port, B1 => 
                           n1162, B2 => REGISTERS_26_1_port, ZN => n1200);
   U743 : INV_X1 port map( A => REGISTERS_24_1_port, ZN => n81);
   U744 : INV_X1 port map( A => REGISTERS_25_1_port, ZN => n80);
   U745 : OAI221_X1 port map( B1 => n83, B2 => n1163, C1 => n84, C2 => n1164, A
                           => n1201, ZN => n1194);
   U746 : AOI22_X1 port map( A1 => n1166, A2 => REGISTERS_29_1_port, B1 => 
                           n1167, B2 => REGISTERS_28_1_port, ZN => n1201);
   U747 : INV_X1 port map( A => REGISTERS_30_1_port, ZN => n84);
   U748 : INV_X1 port map( A => REGISTERS_31_1_port, ZN => n83);
   U749 : NOR4_X1 port map( A1 => n1202, A2 => n1203, A3 => n1204, A4 => n1205,
                           ZN => n1192);
   U751 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_3_1_port, B1 => n1176
                           , B2 => REGISTERS_2_1_port, ZN => n1206);
   U752 : INV_X1 port map( A => REGISTERS_1_1_port, ZN => n90);
   U753 : OAI221_X1 port map( B1 => n93, B2 => n1177, C1 => n94, C2 => n1178, A
                           => n1207, ZN => n1204);
   U754 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_7_1_port, B1 => n1181
                           , B2 => REGISTERS_6_1_port, ZN => n1207);
   U755 : INV_X1 port map( A => REGISTERS_4_1_port, ZN => n94);
   U756 : INV_X1 port map( A => REGISTERS_5_1_port, ZN => n93);
   U757 : OAI221_X1 port map( B1 => n96, B2 => n1182, C1 => n97, C2 => n1183, A
                           => n1208, ZN => n1203);
   U758 : AOI22_X1 port map( A1 => n1185, A2 => REGISTERS_11_1_port, B1 => 
                           n1186, B2 => REGISTERS_10_1_port, ZN => n1208);
   U759 : INV_X1 port map( A => REGISTERS_8_1_port, ZN => n97);
   U760 : INV_X1 port map( A => REGISTERS_9_1_port, ZN => n96);
   U761 : OAI221_X1 port map( B1 => n99, B2 => n1187, C1 => n100, C2 => n1188, 
                           A => n1209, ZN => n1202);
   U762 : AOI22_X1 port map( A1 => n1190, A2 => REGISTERS_15_1_port, B1 => 
                           n1191, B2 => REGISTERS_14_1_port, ZN => n1209);
   U763 : INV_X1 port map( A => REGISTERS_12_1_port, ZN => n100);
   U764 : INV_X1 port map( A => REGISTERS_13_1_port, ZN => n99);
   U765 : NAND2_X1 port map( A1 => n1210, A2 => n1211, ZN => N4244);
   U766 : NOR4_X1 port map( A1 => n1212, A2 => n1213, A3 => n1214, A4 => n1215,
                           ZN => n1211);
   U767 : OAI221_X1 port map( B1 => n108, B2 => n1148, C1 => n109, C2 => n1149,
                           A => n1216, ZN => n1215);
   U768 : AOI22_X1 port map( A1 => n1151, A2 => REGISTERS_19_2_port, B1 => 
                           n1152, B2 => REGISTERS_18_2_port, ZN => n1216);
   U769 : INV_X1 port map( A => REGISTERS_16_2_port, ZN => n109);
   U770 : INV_X1 port map( A => REGISTERS_17_2_port, ZN => n108);
   U771 : OAI221_X1 port map( B1 => n111, B2 => n1153, C1 => n112, C2 => n1154,
                           A => n1217, ZN => n1214);
   U772 : AOI22_X1 port map( A1 => n1156, A2 => REGISTERS_23_2_port, B1 => 
                           n1157, B2 => REGISTERS_22_2_port, ZN => n1217);
   U773 : INV_X1 port map( A => REGISTERS_20_2_port, ZN => n112);
   U774 : INV_X1 port map( A => REGISTERS_21_2_port, ZN => n111);
   U775 : OAI221_X1 port map( B1 => n114, B2 => n1158, C1 => n115, C2 => n1159,
                           A => n1218, ZN => n1213);
   U776 : AOI22_X1 port map( A1 => n1161, A2 => REGISTERS_27_2_port, B1 => 
                           n1162, B2 => REGISTERS_26_2_port, ZN => n1218);
   U777 : INV_X1 port map( A => REGISTERS_24_2_port, ZN => n115);
   U778 : INV_X1 port map( A => REGISTERS_25_2_port, ZN => n114);
   U779 : OAI221_X1 port map( B1 => n117, B2 => n1163, C1 => n118, C2 => n1164,
                           A => n1219, ZN => n1212);
   U780 : AOI22_X1 port map( A1 => n1166, A2 => REGISTERS_29_2_port, B1 => 
                           n1167, B2 => REGISTERS_28_2_port, ZN => n1219);
   U781 : INV_X1 port map( A => REGISTERS_30_2_port, ZN => n118);
   U782 : INV_X1 port map( A => REGISTERS_31_2_port, ZN => n117);
   U783 : NOR4_X1 port map( A1 => n1220, A2 => n1221, A3 => n1222, A4 => n1223,
                           ZN => n1210);
   U785 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_3_2_port, B1 => n1176
                           , B2 => REGISTERS_2_2_port, ZN => n1224);
   U786 : INV_X1 port map( A => REGISTERS_1_2_port, ZN => n124);
   U787 : OAI221_X1 port map( B1 => n127, B2 => n1177, C1 => n128, C2 => n1178,
                           A => n1225, ZN => n1222);
   U788 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_7_2_port, B1 => n1181
                           , B2 => REGISTERS_6_2_port, ZN => n1225);
   U789 : INV_X1 port map( A => REGISTERS_4_2_port, ZN => n128);
   U790 : INV_X1 port map( A => REGISTERS_5_2_port, ZN => n127);
   U791 : OAI221_X1 port map( B1 => n130, B2 => n1182, C1 => n131, C2 => n1183,
                           A => n1226, ZN => n1221);
   U792 : AOI22_X1 port map( A1 => n1185, A2 => REGISTERS_11_2_port, B1 => 
                           n1186, B2 => REGISTERS_10_2_port, ZN => n1226);
   U793 : INV_X1 port map( A => REGISTERS_8_2_port, ZN => n131);
   U794 : INV_X1 port map( A => REGISTERS_9_2_port, ZN => n130);
   U795 : OAI221_X1 port map( B1 => n133, B2 => n1187, C1 => n134, C2 => n1188,
                           A => n1227, ZN => n1220);
   U796 : AOI22_X1 port map( A1 => n1190, A2 => REGISTERS_15_2_port, B1 => 
                           n1191, B2 => REGISTERS_14_2_port, ZN => n1227);
   U797 : INV_X1 port map( A => REGISTERS_12_2_port, ZN => n134);
   U798 : INV_X1 port map( A => REGISTERS_13_2_port, ZN => n133);
   U799 : NAND2_X1 port map( A1 => n1228, A2 => n1229, ZN => N4243);
   U800 : NOR4_X1 port map( A1 => n1230, A2 => n1231, A3 => n1232, A4 => n1233,
                           ZN => n1229);
   U801 : OAI221_X1 port map( B1 => n142, B2 => n1148, C1 => n143, C2 => n1149,
                           A => n1234, ZN => n1233);
   U802 : AOI22_X1 port map( A1 => n1151, A2 => REGISTERS_19_3_port, B1 => 
                           n1152, B2 => REGISTERS_18_3_port, ZN => n1234);
   U803 : INV_X1 port map( A => REGISTERS_16_3_port, ZN => n143);
   U804 : INV_X1 port map( A => REGISTERS_17_3_port, ZN => n142);
   U805 : OAI221_X1 port map( B1 => n145, B2 => n1153, C1 => n146, C2 => n1154,
                           A => n1235, ZN => n1232);
   U806 : AOI22_X1 port map( A1 => n1156, A2 => REGISTERS_23_3_port, B1 => 
                           n1157, B2 => REGISTERS_22_3_port, ZN => n1235);
   U807 : INV_X1 port map( A => REGISTERS_20_3_port, ZN => n146);
   U808 : INV_X1 port map( A => REGISTERS_21_3_port, ZN => n145);
   U809 : OAI221_X1 port map( B1 => n148, B2 => n1158, C1 => n149, C2 => n1159,
                           A => n1236, ZN => n1231);
   U810 : AOI22_X1 port map( A1 => n1161, A2 => REGISTERS_27_3_port, B1 => 
                           n1162, B2 => REGISTERS_26_3_port, ZN => n1236);
   U811 : INV_X1 port map( A => REGISTERS_24_3_port, ZN => n149);
   U812 : INV_X1 port map( A => REGISTERS_25_3_port, ZN => n148);
   U813 : OAI221_X1 port map( B1 => n151, B2 => n1163, C1 => n152, C2 => n1164,
                           A => n1237, ZN => n1230);
   U814 : AOI22_X1 port map( A1 => n1166, A2 => REGISTERS_29_3_port, B1 => 
                           n1167, B2 => REGISTERS_28_3_port, ZN => n1237);
   U815 : INV_X1 port map( A => REGISTERS_30_3_port, ZN => n152);
   U816 : INV_X1 port map( A => REGISTERS_31_3_port, ZN => n151);
   U817 : NOR4_X1 port map( A1 => n1238, A2 => n1239, A3 => n1240, A4 => n1241,
                           ZN => n1228);
   U819 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_3_3_port, B1 => n1176
                           , B2 => REGISTERS_2_3_port, ZN => n1242);
   U820 : INV_X1 port map( A => REGISTERS_1_3_port, ZN => n158);
   U821 : OAI221_X1 port map( B1 => n161, B2 => n1177, C1 => n162, C2 => n1178,
                           A => n1243, ZN => n1240);
   U822 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_7_3_port, B1 => n1181
                           , B2 => REGISTERS_6_3_port, ZN => n1243);
   U823 : INV_X1 port map( A => REGISTERS_4_3_port, ZN => n162);
   U824 : INV_X1 port map( A => REGISTERS_5_3_port, ZN => n161);
   U825 : OAI221_X1 port map( B1 => n164, B2 => n1182, C1 => n165, C2 => n1183,
                           A => n1244, ZN => n1239);
   U826 : AOI22_X1 port map( A1 => n1185, A2 => REGISTERS_11_3_port, B1 => 
                           n1186, B2 => REGISTERS_10_3_port, ZN => n1244);
   U827 : INV_X1 port map( A => REGISTERS_8_3_port, ZN => n165);
   U828 : INV_X1 port map( A => REGISTERS_9_3_port, ZN => n164);
   U829 : OAI221_X1 port map( B1 => n167, B2 => n1187, C1 => n168, C2 => n1188,
                           A => n1245, ZN => n1238);
   U830 : AOI22_X1 port map( A1 => n1190, A2 => REGISTERS_15_3_port, B1 => 
                           n1191, B2 => REGISTERS_14_3_port, ZN => n1245);
   U831 : INV_X1 port map( A => REGISTERS_12_3_port, ZN => n168);
   U832 : INV_X1 port map( A => REGISTERS_13_3_port, ZN => n167);
   U833 : NAND2_X1 port map( A1 => n1246, A2 => n1247, ZN => N4242);
   U834 : NOR4_X1 port map( A1 => n1248, A2 => n1249, A3 => n1250, A4 => n1251,
                           ZN => n1247);
   U835 : OAI221_X1 port map( B1 => n176, B2 => n1148, C1 => n177, C2 => n1149,
                           A => n1252, ZN => n1251);
   U836 : AOI22_X1 port map( A1 => n1151, A2 => REGISTERS_19_4_port, B1 => 
                           n1152, B2 => REGISTERS_18_4_port, ZN => n1252);
   U837 : INV_X1 port map( A => REGISTERS_16_4_port, ZN => n177);
   U838 : INV_X1 port map( A => REGISTERS_17_4_port, ZN => n176);
   U839 : OAI221_X1 port map( B1 => n179, B2 => n1153, C1 => n180, C2 => n1154,
                           A => n1253, ZN => n1250);
   U840 : AOI22_X1 port map( A1 => n1156, A2 => REGISTERS_23_4_port, B1 => 
                           n1157, B2 => REGISTERS_22_4_port, ZN => n1253);
   U841 : INV_X1 port map( A => REGISTERS_20_4_port, ZN => n180);
   U842 : INV_X1 port map( A => REGISTERS_21_4_port, ZN => n179);
   U843 : OAI221_X1 port map( B1 => n182, B2 => n1158, C1 => n183, C2 => n1159,
                           A => n1254, ZN => n1249);
   U844 : AOI22_X1 port map( A1 => n1161, A2 => REGISTERS_27_4_port, B1 => 
                           n1162, B2 => REGISTERS_26_4_port, ZN => n1254);
   U845 : INV_X1 port map( A => REGISTERS_24_4_port, ZN => n183);
   U846 : INV_X1 port map( A => REGISTERS_25_4_port, ZN => n182);
   U847 : OAI221_X1 port map( B1 => n185, B2 => n1163, C1 => n186, C2 => n1164,
                           A => n1255, ZN => n1248);
   U848 : AOI22_X1 port map( A1 => n1166, A2 => REGISTERS_29_4_port, B1 => 
                           n1167, B2 => REGISTERS_28_4_port, ZN => n1255);
   U849 : INV_X1 port map( A => REGISTERS_30_4_port, ZN => n186);
   U850 : INV_X1 port map( A => REGISTERS_31_4_port, ZN => n185);
   U851 : NOR4_X1 port map( A1 => n1256, A2 => n1257, A3 => n1258, A4 => n1259,
                           ZN => n1246);
   U853 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_3_4_port, B1 => n1176
                           , B2 => REGISTERS_2_4_port, ZN => n1260);
   U854 : INV_X1 port map( A => REGISTERS_1_4_port, ZN => n192);
   U855 : OAI221_X1 port map( B1 => n195, B2 => n1177, C1 => n196, C2 => n1178,
                           A => n1261, ZN => n1258);
   U856 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_7_4_port, B1 => n1181
                           , B2 => REGISTERS_6_4_port, ZN => n1261);
   U857 : INV_X1 port map( A => REGISTERS_4_4_port, ZN => n196);
   U858 : INV_X1 port map( A => REGISTERS_5_4_port, ZN => n195);
   U859 : OAI221_X1 port map( B1 => n198, B2 => n1182, C1 => n199, C2 => n1183,
                           A => n1262, ZN => n1257);
   U860 : AOI22_X1 port map( A1 => n1185, A2 => REGISTERS_11_4_port, B1 => 
                           n1186, B2 => REGISTERS_10_4_port, ZN => n1262);
   U861 : INV_X1 port map( A => REGISTERS_8_4_port, ZN => n199);
   U862 : INV_X1 port map( A => REGISTERS_9_4_port, ZN => n198);
   U863 : OAI221_X1 port map( B1 => n201, B2 => n1187, C1 => n202, C2 => n1188,
                           A => n1263, ZN => n1256);
   U864 : AOI22_X1 port map( A1 => n1190, A2 => REGISTERS_15_4_port, B1 => 
                           n1191, B2 => REGISTERS_14_4_port, ZN => n1263);
   U865 : INV_X1 port map( A => REGISTERS_12_4_port, ZN => n202);
   U866 : INV_X1 port map( A => REGISTERS_13_4_port, ZN => n201);
   U867 : NAND2_X1 port map( A1 => n1264, A2 => n1265, ZN => N4241);
   U868 : NOR4_X1 port map( A1 => n1266, A2 => n1267, A3 => n1268, A4 => n1269,
                           ZN => n1265);
   U869 : OAI221_X1 port map( B1 => n210, B2 => n1148, C1 => n211, C2 => n1149,
                           A => n1270, ZN => n1269);
   U870 : AOI22_X1 port map( A1 => n1151, A2 => REGISTERS_19_5_port, B1 => 
                           n1152, B2 => REGISTERS_18_5_port, ZN => n1270);
   U871 : INV_X1 port map( A => REGISTERS_16_5_port, ZN => n211);
   U872 : INV_X1 port map( A => REGISTERS_17_5_port, ZN => n210);
   U873 : OAI221_X1 port map( B1 => n213, B2 => n1153, C1 => n214, C2 => n1154,
                           A => n1271, ZN => n1268);
   U874 : AOI22_X1 port map( A1 => n1156, A2 => REGISTERS_23_5_port, B1 => 
                           n1157, B2 => REGISTERS_22_5_port, ZN => n1271);
   U875 : INV_X1 port map( A => REGISTERS_20_5_port, ZN => n214);
   U876 : INV_X1 port map( A => REGISTERS_21_5_port, ZN => n213);
   U877 : OAI221_X1 port map( B1 => n216, B2 => n1158, C1 => n217, C2 => n1159,
                           A => n1272, ZN => n1267);
   U878 : AOI22_X1 port map( A1 => n1161, A2 => REGISTERS_27_5_port, B1 => 
                           n1162, B2 => REGISTERS_26_5_port, ZN => n1272);
   U879 : INV_X1 port map( A => REGISTERS_24_5_port, ZN => n217);
   U880 : INV_X1 port map( A => REGISTERS_25_5_port, ZN => n216);
   U881 : OAI221_X1 port map( B1 => n219, B2 => n1163, C1 => n220, C2 => n1164,
                           A => n1273, ZN => n1266);
   U882 : AOI22_X1 port map( A1 => n1166, A2 => REGISTERS_29_5_port, B1 => 
                           n1167, B2 => REGISTERS_28_5_port, ZN => n1273);
   U883 : INV_X1 port map( A => REGISTERS_30_5_port, ZN => n220);
   U884 : INV_X1 port map( A => REGISTERS_31_5_port, ZN => n219);
   U885 : NOR4_X1 port map( A1 => n1274, A2 => n1275, A3 => n1276, A4 => n1277,
                           ZN => n1264);
   U887 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_3_5_port, B1 => n1176
                           , B2 => REGISTERS_2_5_port, ZN => n1278);
   U888 : INV_X1 port map( A => REGISTERS_1_5_port, ZN => n226);
   U889 : OAI221_X1 port map( B1 => n229, B2 => n1177, C1 => n230, C2 => n1178,
                           A => n1279, ZN => n1276);
   U890 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_7_5_port, B1 => n1181
                           , B2 => REGISTERS_6_5_port, ZN => n1279);
   U891 : INV_X1 port map( A => REGISTERS_4_5_port, ZN => n230);
   U892 : INV_X1 port map( A => REGISTERS_5_5_port, ZN => n229);
   U893 : OAI221_X1 port map( B1 => n232, B2 => n1182, C1 => n233, C2 => n1183,
                           A => n1280, ZN => n1275);
   U894 : AOI22_X1 port map( A1 => n1185, A2 => REGISTERS_11_5_port, B1 => 
                           n1186, B2 => REGISTERS_10_5_port, ZN => n1280);
   U895 : INV_X1 port map( A => REGISTERS_8_5_port, ZN => n233);
   U896 : INV_X1 port map( A => REGISTERS_9_5_port, ZN => n232);
   U897 : OAI221_X1 port map( B1 => n235, B2 => n1187, C1 => n236, C2 => n1188,
                           A => n1281, ZN => n1274);
   U898 : AOI22_X1 port map( A1 => n1190, A2 => REGISTERS_15_5_port, B1 => 
                           n1191, B2 => REGISTERS_14_5_port, ZN => n1281);
   U899 : INV_X1 port map( A => REGISTERS_12_5_port, ZN => n236);
   U900 : INV_X1 port map( A => REGISTERS_13_5_port, ZN => n235);
   U901 : NAND2_X1 port map( A1 => n1282, A2 => n1283, ZN => N4240);
   U902 : NOR4_X1 port map( A1 => n1284, A2 => n1285, A3 => n1286, A4 => n1287,
                           ZN => n1283);
   U903 : OAI221_X1 port map( B1 => n244, B2 => n1148, C1 => n245, C2 => n1149,
                           A => n1288, ZN => n1287);
   U904 : AOI22_X1 port map( A1 => n1151, A2 => REGISTERS_19_6_port, B1 => 
                           n1152, B2 => REGISTERS_18_6_port, ZN => n1288);
   U905 : INV_X1 port map( A => REGISTERS_16_6_port, ZN => n245);
   U906 : INV_X1 port map( A => REGISTERS_17_6_port, ZN => n244);
   U907 : OAI221_X1 port map( B1 => n247, B2 => n1153, C1 => n248, C2 => n1154,
                           A => n1289, ZN => n1286);
   U908 : AOI22_X1 port map( A1 => n1156, A2 => REGISTERS_23_6_port, B1 => 
                           n1157, B2 => REGISTERS_22_6_port, ZN => n1289);
   U909 : INV_X1 port map( A => REGISTERS_20_6_port, ZN => n248);
   U910 : INV_X1 port map( A => REGISTERS_21_6_port, ZN => n247);
   U911 : OAI221_X1 port map( B1 => n250, B2 => n1158, C1 => n251, C2 => n1159,
                           A => n1290, ZN => n1285);
   U912 : AOI22_X1 port map( A1 => n1161, A2 => REGISTERS_27_6_port, B1 => 
                           n1162, B2 => REGISTERS_26_6_port, ZN => n1290);
   U913 : INV_X1 port map( A => REGISTERS_24_6_port, ZN => n251);
   U914 : INV_X1 port map( A => REGISTERS_25_6_port, ZN => n250);
   U915 : OAI221_X1 port map( B1 => n253, B2 => n1163, C1 => n254, C2 => n1164,
                           A => n1291, ZN => n1284);
   U916 : AOI22_X1 port map( A1 => n1166, A2 => REGISTERS_29_6_port, B1 => 
                           n1167, B2 => REGISTERS_28_6_port, ZN => n1291);
   U917 : INV_X1 port map( A => REGISTERS_30_6_port, ZN => n254);
   U918 : INV_X1 port map( A => REGISTERS_31_6_port, ZN => n253);
   U919 : NOR4_X1 port map( A1 => n1292, A2 => n1293, A3 => n1294, A4 => n1295,
                           ZN => n1282);
   U921 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_3_6_port, B1 => n1176
                           , B2 => REGISTERS_2_6_port, ZN => n1296);
   U922 : INV_X1 port map( A => REGISTERS_1_6_port, ZN => n260);
   U923 : OAI221_X1 port map( B1 => n263, B2 => n1177, C1 => n264, C2 => n1178,
                           A => n1297, ZN => n1294);
   U924 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_7_6_port, B1 => n1181
                           , B2 => REGISTERS_6_6_port, ZN => n1297);
   U925 : INV_X1 port map( A => REGISTERS_4_6_port, ZN => n264);
   U926 : INV_X1 port map( A => REGISTERS_5_6_port, ZN => n263);
   U927 : OAI221_X1 port map( B1 => n266, B2 => n1182, C1 => n267, C2 => n1183,
                           A => n1298, ZN => n1293);
   U928 : AOI22_X1 port map( A1 => n1185, A2 => REGISTERS_11_6_port, B1 => 
                           n1186, B2 => REGISTERS_10_6_port, ZN => n1298);
   U929 : INV_X1 port map( A => REGISTERS_8_6_port, ZN => n267);
   U930 : INV_X1 port map( A => REGISTERS_9_6_port, ZN => n266);
   U931 : OAI221_X1 port map( B1 => n269, B2 => n1187, C1 => n270, C2 => n1188,
                           A => n1299, ZN => n1292);
   U932 : AOI22_X1 port map( A1 => n1190, A2 => REGISTERS_15_6_port, B1 => 
                           n1191, B2 => REGISTERS_14_6_port, ZN => n1299);
   U933 : INV_X1 port map( A => REGISTERS_12_6_port, ZN => n270);
   U934 : INV_X1 port map( A => REGISTERS_13_6_port, ZN => n269);
   U935 : NAND2_X1 port map( A1 => n1300, A2 => n1301, ZN => N4239);
   U936 : NOR4_X1 port map( A1 => n1302, A2 => n1303, A3 => n1304, A4 => n1305,
                           ZN => n1301);
   U937 : OAI221_X1 port map( B1 => n278, B2 => n1148, C1 => n279, C2 => n1149,
                           A => n1306, ZN => n1305);
   U938 : AOI22_X1 port map( A1 => n1151, A2 => REGISTERS_19_7_port, B1 => 
                           n1152, B2 => REGISTERS_18_7_port, ZN => n1306);
   U939 : INV_X1 port map( A => REGISTERS_16_7_port, ZN => n279);
   U940 : INV_X1 port map( A => REGISTERS_17_7_port, ZN => n278);
   U941 : OAI221_X1 port map( B1 => n281, B2 => n1153, C1 => n282, C2 => n1154,
                           A => n1307, ZN => n1304);
   U942 : AOI22_X1 port map( A1 => n1156, A2 => REGISTERS_23_7_port, B1 => 
                           n1157, B2 => REGISTERS_22_7_port, ZN => n1307);
   U943 : INV_X1 port map( A => REGISTERS_20_7_port, ZN => n282);
   U944 : INV_X1 port map( A => REGISTERS_21_7_port, ZN => n281);
   U945 : OAI221_X1 port map( B1 => n284, B2 => n1158, C1 => n285, C2 => n1159,
                           A => n1308, ZN => n1303);
   U946 : AOI22_X1 port map( A1 => n1161, A2 => REGISTERS_27_7_port, B1 => 
                           n1162, B2 => REGISTERS_26_7_port, ZN => n1308);
   U947 : INV_X1 port map( A => REGISTERS_24_7_port, ZN => n285);
   U948 : INV_X1 port map( A => REGISTERS_25_7_port, ZN => n284);
   U949 : OAI221_X1 port map( B1 => n287, B2 => n1163, C1 => n288, C2 => n1164,
                           A => n1309, ZN => n1302);
   U950 : AOI22_X1 port map( A1 => n1166, A2 => REGISTERS_29_7_port, B1 => 
                           n1167, B2 => REGISTERS_28_7_port, ZN => n1309);
   U951 : INV_X1 port map( A => REGISTERS_30_7_port, ZN => n288);
   U952 : INV_X1 port map( A => REGISTERS_31_7_port, ZN => n287);
   U953 : NOR4_X1 port map( A1 => n1310, A2 => n1311, A3 => n1312, A4 => n1313,
                           ZN => n1300);
   U955 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_3_7_port, B1 => n1176
                           , B2 => REGISTERS_2_7_port, ZN => n1314);
   U956 : INV_X1 port map( A => REGISTERS_1_7_port, ZN => n294);
   U957 : OAI221_X1 port map( B1 => n297, B2 => n1177, C1 => n298, C2 => n1178,
                           A => n1315, ZN => n1312);
   U958 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_7_7_port, B1 => n1181
                           , B2 => REGISTERS_6_7_port, ZN => n1315);
   U959 : INV_X1 port map( A => REGISTERS_4_7_port, ZN => n298);
   U960 : INV_X1 port map( A => REGISTERS_5_7_port, ZN => n297);
   U961 : OAI221_X1 port map( B1 => n300, B2 => n1182, C1 => n301, C2 => n1183,
                           A => n1316, ZN => n1311);
   U962 : AOI22_X1 port map( A1 => n1185, A2 => REGISTERS_11_7_port, B1 => 
                           n1186, B2 => REGISTERS_10_7_port, ZN => n1316);
   U963 : INV_X1 port map( A => REGISTERS_8_7_port, ZN => n301);
   U964 : INV_X1 port map( A => REGISTERS_9_7_port, ZN => n300);
   U965 : OAI221_X1 port map( B1 => n303, B2 => n1187, C1 => n304, C2 => n1188,
                           A => n1317, ZN => n1310);
   U966 : AOI22_X1 port map( A1 => n1190, A2 => REGISTERS_15_7_port, B1 => 
                           n1191, B2 => REGISTERS_14_7_port, ZN => n1317);
   U967 : INV_X1 port map( A => REGISTERS_12_7_port, ZN => n304);
   U968 : INV_X1 port map( A => REGISTERS_13_7_port, ZN => n303);
   U969 : NAND2_X1 port map( A1 => n1318, A2 => n1319, ZN => N4238);
   U970 : NOR4_X1 port map( A1 => n1320, A2 => n1321, A3 => n1322, A4 => n1323,
                           ZN => n1319);
   U971 : OAI221_X1 port map( B1 => n312, B2 => n1148, C1 => n313, C2 => n1149,
                           A => n1324, ZN => n1323);
   U972 : AOI22_X1 port map( A1 => n1151, A2 => REGISTERS_19_8_port, B1 => 
                           n1152, B2 => REGISTERS_18_8_port, ZN => n1324);
   U973 : INV_X1 port map( A => REGISTERS_16_8_port, ZN => n313);
   U974 : INV_X1 port map( A => REGISTERS_17_8_port, ZN => n312);
   U975 : OAI221_X1 port map( B1 => n315, B2 => n1153, C1 => n316, C2 => n1154,
                           A => n1325, ZN => n1322);
   U976 : AOI22_X1 port map( A1 => n1156, A2 => REGISTERS_23_8_port, B1 => 
                           n1157, B2 => REGISTERS_22_8_port, ZN => n1325);
   U977 : INV_X1 port map( A => REGISTERS_20_8_port, ZN => n316);
   U978 : INV_X1 port map( A => REGISTERS_21_8_port, ZN => n315);
   U979 : OAI221_X1 port map( B1 => n318, B2 => n1158, C1 => n319, C2 => n1159,
                           A => n1326, ZN => n1321);
   U980 : AOI22_X1 port map( A1 => n1161, A2 => REGISTERS_27_8_port, B1 => 
                           n1162, B2 => REGISTERS_26_8_port, ZN => n1326);
   U981 : INV_X1 port map( A => REGISTERS_24_8_port, ZN => n319);
   U982 : INV_X1 port map( A => REGISTERS_25_8_port, ZN => n318);
   U983 : OAI221_X1 port map( B1 => n321, B2 => n1163, C1 => n322, C2 => n1164,
                           A => n1327, ZN => n1320);
   U984 : AOI22_X1 port map( A1 => n1166, A2 => REGISTERS_29_8_port, B1 => 
                           n1167, B2 => REGISTERS_28_8_port, ZN => n1327);
   U985 : INV_X1 port map( A => REGISTERS_30_8_port, ZN => n322);
   U986 : INV_X1 port map( A => REGISTERS_31_8_port, ZN => n321);
   U987 : NOR4_X1 port map( A1 => n1328, A2 => n1329, A3 => n1330, A4 => n1331,
                           ZN => n1318);
   U989 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_3_8_port, B1 => n1176
                           , B2 => REGISTERS_2_8_port, ZN => n1332);
   U990 : INV_X1 port map( A => REGISTERS_1_8_port, ZN => n328);
   U991 : OAI221_X1 port map( B1 => n331, B2 => n1177, C1 => n332, C2 => n1178,
                           A => n1333, ZN => n1330);
   U992 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_7_8_port, B1 => n1181
                           , B2 => REGISTERS_6_8_port, ZN => n1333);
   U993 : INV_X1 port map( A => REGISTERS_4_8_port, ZN => n332);
   U994 : INV_X1 port map( A => REGISTERS_5_8_port, ZN => n331);
   U995 : OAI221_X1 port map( B1 => n334, B2 => n1182, C1 => n335, C2 => n1183,
                           A => n1334, ZN => n1329);
   U996 : AOI22_X1 port map( A1 => n1185, A2 => REGISTERS_11_8_port, B1 => 
                           n1186, B2 => REGISTERS_10_8_port, ZN => n1334);
   U997 : INV_X1 port map( A => REGISTERS_8_8_port, ZN => n335);
   U998 : INV_X1 port map( A => REGISTERS_9_8_port, ZN => n334);
   U999 : OAI221_X1 port map( B1 => n337, B2 => n1187, C1 => n338, C2 => n1188,
                           A => n1335, ZN => n1328);
   U1000 : AOI22_X1 port map( A1 => n1190, A2 => REGISTERS_15_8_port, B1 => 
                           n1191, B2 => REGISTERS_14_8_port, ZN => n1335);
   U1001 : INV_X1 port map( A => REGISTERS_12_8_port, ZN => n338);
   U1002 : INV_X1 port map( A => REGISTERS_13_8_port, ZN => n337);
   U1003 : NAND2_X1 port map( A1 => n1336, A2 => n1337, ZN => N4237);
   U1004 : NOR4_X1 port map( A1 => n1338, A2 => n1339, A3 => n1340, A4 => n1341
                           , ZN => n1337);
   U1005 : OAI221_X1 port map( B1 => n346, B2 => n1148, C1 => n347, C2 => n1149
                           , A => n1342, ZN => n1341);
   U1006 : AOI22_X1 port map( A1 => n1151, A2 => REGISTERS_19_9_port, B1 => 
                           n1152, B2 => REGISTERS_18_9_port, ZN => n1342);
   U1007 : INV_X1 port map( A => REGISTERS_16_9_port, ZN => n347);
   U1008 : INV_X1 port map( A => REGISTERS_17_9_port, ZN => n346);
   U1009 : OAI221_X1 port map( B1 => n349, B2 => n1153, C1 => n350, C2 => n1154
                           , A => n1343, ZN => n1340);
   U1010 : AOI22_X1 port map( A1 => n1156, A2 => REGISTERS_23_9_port, B1 => 
                           n1157, B2 => REGISTERS_22_9_port, ZN => n1343);
   U1011 : INV_X1 port map( A => REGISTERS_20_9_port, ZN => n350);
   U1012 : INV_X1 port map( A => REGISTERS_21_9_port, ZN => n349);
   U1013 : OAI221_X1 port map( B1 => n352, B2 => n1158, C1 => n353, C2 => n1159
                           , A => n1344, ZN => n1339);
   U1014 : AOI22_X1 port map( A1 => n1161, A2 => REGISTERS_27_9_port, B1 => 
                           n1162, B2 => REGISTERS_26_9_port, ZN => n1344);
   U1015 : INV_X1 port map( A => REGISTERS_24_9_port, ZN => n353);
   U1016 : INV_X1 port map( A => REGISTERS_25_9_port, ZN => n352);
   U1017 : OAI221_X1 port map( B1 => n355, B2 => n1163, C1 => n356, C2 => n1164
                           , A => n1345, ZN => n1338);
   U1018 : AOI22_X1 port map( A1 => n1166, A2 => REGISTERS_29_9_port, B1 => 
                           n1167, B2 => REGISTERS_28_9_port, ZN => n1345);
   U1019 : INV_X1 port map( A => REGISTERS_30_9_port, ZN => n356);
   U1020 : INV_X1 port map( A => REGISTERS_31_9_port, ZN => n355);
   U1021 : NOR4_X1 port map( A1 => n1346, A2 => n1347, A3 => n1348, A4 => n1349
                           , ZN => n1336);
   U1023 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_3_9_port, B1 => 
                           n1176, B2 => REGISTERS_2_9_port, ZN => n1350);
   U1024 : INV_X1 port map( A => REGISTERS_1_9_port, ZN => n362);
   U1025 : OAI221_X1 port map( B1 => n365, B2 => n1177, C1 => n366, C2 => n1178
                           , A => n1351, ZN => n1348);
   U1026 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_7_9_port, B1 => 
                           n1181, B2 => REGISTERS_6_9_port, ZN => n1351);
   U1027 : INV_X1 port map( A => REGISTERS_4_9_port, ZN => n366);
   U1028 : INV_X1 port map( A => REGISTERS_5_9_port, ZN => n365);
   U1029 : OAI221_X1 port map( B1 => n368, B2 => n1182, C1 => n369, C2 => n1183
                           , A => n1352, ZN => n1347);
   U1030 : AOI22_X1 port map( A1 => n1185, A2 => REGISTERS_11_9_port, B1 => 
                           n1186, B2 => REGISTERS_10_9_port, ZN => n1352);
   U1031 : INV_X1 port map( A => REGISTERS_8_9_port, ZN => n369);
   U1032 : INV_X1 port map( A => REGISTERS_9_9_port, ZN => n368);
   U1033 : OAI221_X1 port map( B1 => n371, B2 => n1187, C1 => n372, C2 => n1188
                           , A => n1353, ZN => n1346);
   U1034 : AOI22_X1 port map( A1 => n1190, A2 => REGISTERS_15_9_port, B1 => 
                           n1191, B2 => REGISTERS_14_9_port, ZN => n1353);
   U1035 : INV_X1 port map( A => REGISTERS_12_9_port, ZN => n372);
   U1036 : INV_X1 port map( A => REGISTERS_13_9_port, ZN => n371);
   U1037 : NAND2_X1 port map( A1 => n1354, A2 => n1355, ZN => N4236);
   U1038 : NOR4_X1 port map( A1 => n1356, A2 => n1357, A3 => n1358, A4 => n1359
                           , ZN => n1355);
   U1039 : OAI221_X1 port map( B1 => n380, B2 => n1148, C1 => n381, C2 => n1149
                           , A => n1360, ZN => n1359);
   U1040 : AOI22_X1 port map( A1 => n1151, A2 => REGISTERS_19_10_port, B1 => 
                           n1152, B2 => REGISTERS_18_10_port, ZN => n1360);
   U1041 : INV_X1 port map( A => REGISTERS_16_10_port, ZN => n381);
   U1042 : INV_X1 port map( A => REGISTERS_17_10_port, ZN => n380);
   U1043 : OAI221_X1 port map( B1 => n383, B2 => n1153, C1 => n384, C2 => n1154
                           , A => n1361, ZN => n1358);
   U1044 : AOI22_X1 port map( A1 => n1156, A2 => REGISTERS_23_10_port, B1 => 
                           n1157, B2 => REGISTERS_22_10_port, ZN => n1361);
   U1045 : INV_X1 port map( A => REGISTERS_20_10_port, ZN => n384);
   U1046 : INV_X1 port map( A => REGISTERS_21_10_port, ZN => n383);
   U1047 : OAI221_X1 port map( B1 => n386, B2 => n1158, C1 => n387, C2 => n1159
                           , A => n1362, ZN => n1357);
   U1048 : AOI22_X1 port map( A1 => n1161, A2 => REGISTERS_27_10_port, B1 => 
                           n1162, B2 => REGISTERS_26_10_port, ZN => n1362);
   U1049 : INV_X1 port map( A => REGISTERS_24_10_port, ZN => n387);
   U1050 : INV_X1 port map( A => REGISTERS_25_10_port, ZN => n386);
   U1051 : OAI221_X1 port map( B1 => n389, B2 => n1163, C1 => n390, C2 => n1164
                           , A => n1363, ZN => n1356);
   U1052 : AOI22_X1 port map( A1 => n1166, A2 => REGISTERS_29_10_port, B1 => 
                           n1167, B2 => REGISTERS_28_10_port, ZN => n1363);
   U1053 : INV_X1 port map( A => REGISTERS_30_10_port, ZN => n390);
   U1054 : INV_X1 port map( A => REGISTERS_31_10_port, ZN => n389);
   U1055 : NOR4_X1 port map( A1 => n1364, A2 => n1365, A3 => n1366, A4 => n1367
                           , ZN => n1354);
   U1057 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_3_10_port, B1 => 
                           n1176, B2 => REGISTERS_2_10_port, ZN => n1368);
   U1058 : INV_X1 port map( A => REGISTERS_1_10_port, ZN => n396);
   U1059 : OAI221_X1 port map( B1 => n399, B2 => n1177, C1 => n400, C2 => n1178
                           , A => n1369, ZN => n1366);
   U1060 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_7_10_port, B1 => 
                           n1181, B2 => REGISTERS_6_10_port, ZN => n1369);
   U1061 : INV_X1 port map( A => REGISTERS_4_10_port, ZN => n400);
   U1062 : INV_X1 port map( A => REGISTERS_5_10_port, ZN => n399);
   U1063 : OAI221_X1 port map( B1 => n402, B2 => n1182, C1 => n403, C2 => n1183
                           , A => n1370, ZN => n1365);
   U1064 : AOI22_X1 port map( A1 => n1185, A2 => REGISTERS_11_10_port, B1 => 
                           n1186, B2 => REGISTERS_10_10_port, ZN => n1370);
   U1065 : INV_X1 port map( A => REGISTERS_8_10_port, ZN => n403);
   U1066 : INV_X1 port map( A => REGISTERS_9_10_port, ZN => n402);
   U1067 : OAI221_X1 port map( B1 => n405, B2 => n1187, C1 => n406, C2 => n1188
                           , A => n1371, ZN => n1364);
   U1068 : AOI22_X1 port map( A1 => n1190, A2 => REGISTERS_15_10_port, B1 => 
                           n1191, B2 => REGISTERS_14_10_port, ZN => n1371);
   U1069 : INV_X1 port map( A => REGISTERS_12_10_port, ZN => n406);
   U1070 : INV_X1 port map( A => REGISTERS_13_10_port, ZN => n405);
   U1071 : NAND2_X1 port map( A1 => n1372, A2 => n1373, ZN => N4235);
   U1072 : NOR4_X1 port map( A1 => n1374, A2 => n1375, A3 => n1376, A4 => n1377
                           , ZN => n1373);
   U1073 : OAI221_X1 port map( B1 => n414, B2 => n1148, C1 => n415, C2 => n1149
                           , A => n1378, ZN => n1377);
   U1074 : AOI22_X1 port map( A1 => n1151, A2 => REGISTERS_19_11_port, B1 => 
                           n1152, B2 => REGISTERS_18_11_port, ZN => n1378);
   U1075 : INV_X1 port map( A => REGISTERS_16_11_port, ZN => n415);
   U1076 : INV_X1 port map( A => REGISTERS_17_11_port, ZN => n414);
   U1077 : OAI221_X1 port map( B1 => n417, B2 => n1153, C1 => n418, C2 => n1154
                           , A => n1379, ZN => n1376);
   U1078 : AOI22_X1 port map( A1 => n1156, A2 => REGISTERS_23_11_port, B1 => 
                           n1157, B2 => REGISTERS_22_11_port, ZN => n1379);
   U1079 : INV_X1 port map( A => REGISTERS_20_11_port, ZN => n418);
   U1080 : INV_X1 port map( A => REGISTERS_21_11_port, ZN => n417);
   U1081 : OAI221_X1 port map( B1 => n420, B2 => n1158, C1 => n421, C2 => n1159
                           , A => n1380, ZN => n1375);
   U1082 : AOI22_X1 port map( A1 => n1161, A2 => REGISTERS_27_11_port, B1 => 
                           n1162, B2 => REGISTERS_26_11_port, ZN => n1380);
   U1083 : INV_X1 port map( A => REGISTERS_24_11_port, ZN => n421);
   U1084 : INV_X1 port map( A => REGISTERS_25_11_port, ZN => n420);
   U1085 : OAI221_X1 port map( B1 => n423, B2 => n1163, C1 => n424, C2 => n1164
                           , A => n1381, ZN => n1374);
   U1086 : AOI22_X1 port map( A1 => n1166, A2 => REGISTERS_29_11_port, B1 => 
                           n1167, B2 => REGISTERS_28_11_port, ZN => n1381);
   U1087 : INV_X1 port map( A => REGISTERS_30_11_port, ZN => n424);
   U1088 : INV_X1 port map( A => REGISTERS_31_11_port, ZN => n423);
   U1089 : NOR4_X1 port map( A1 => n1382, A2 => n1383, A3 => n1384, A4 => n1385
                           , ZN => n1372);
   U1091 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_3_11_port, B1 => 
                           n1176, B2 => REGISTERS_2_11_port, ZN => n1386);
   U1092 : INV_X1 port map( A => REGISTERS_1_11_port, ZN => n430);
   U1093 : OAI221_X1 port map( B1 => n433, B2 => n1177, C1 => n434, C2 => n1178
                           , A => n1387, ZN => n1384);
   U1094 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_7_11_port, B1 => 
                           n1181, B2 => REGISTERS_6_11_port, ZN => n1387);
   U1095 : INV_X1 port map( A => REGISTERS_4_11_port, ZN => n434);
   U1096 : INV_X1 port map( A => REGISTERS_5_11_port, ZN => n433);
   U1097 : OAI221_X1 port map( B1 => n436, B2 => n1182, C1 => n437, C2 => n1183
                           , A => n1388, ZN => n1383);
   U1098 : AOI22_X1 port map( A1 => n1185, A2 => REGISTERS_11_11_port, B1 => 
                           n1186, B2 => REGISTERS_10_11_port, ZN => n1388);
   U1099 : INV_X1 port map( A => REGISTERS_8_11_port, ZN => n437);
   U1100 : INV_X1 port map( A => REGISTERS_9_11_port, ZN => n436);
   U1101 : OAI221_X1 port map( B1 => n439, B2 => n1187, C1 => n440, C2 => n1188
                           , A => n1389, ZN => n1382);
   U1102 : AOI22_X1 port map( A1 => n1190, A2 => REGISTERS_15_11_port, B1 => 
                           n1191, B2 => REGISTERS_14_11_port, ZN => n1389);
   U1103 : INV_X1 port map( A => REGISTERS_12_11_port, ZN => n440);
   U1104 : INV_X1 port map( A => REGISTERS_13_11_port, ZN => n439);
   U1105 : NAND2_X1 port map( A1 => n1390, A2 => n1391, ZN => N4234);
   U1106 : NOR4_X1 port map( A1 => n1392, A2 => n1393, A3 => n1394, A4 => n1395
                           , ZN => n1391);
   U1107 : OAI221_X1 port map( B1 => n448, B2 => n1148, C1 => n449, C2 => n1149
                           , A => n1396, ZN => n1395);
   U1108 : AOI22_X1 port map( A1 => n1151, A2 => REGISTERS_19_12_port, B1 => 
                           n1152, B2 => REGISTERS_18_12_port, ZN => n1396);
   U1109 : INV_X1 port map( A => REGISTERS_16_12_port, ZN => n449);
   U1110 : INV_X1 port map( A => REGISTERS_17_12_port, ZN => n448);
   U1111 : OAI221_X1 port map( B1 => n451, B2 => n1153, C1 => n452, C2 => n1154
                           , A => n1397, ZN => n1394);
   U1112 : AOI22_X1 port map( A1 => n1156, A2 => REGISTERS_23_12_port, B1 => 
                           n1157, B2 => REGISTERS_22_12_port, ZN => n1397);
   U1113 : INV_X1 port map( A => REGISTERS_20_12_port, ZN => n452);
   U1114 : INV_X1 port map( A => REGISTERS_21_12_port, ZN => n451);
   U1115 : OAI221_X1 port map( B1 => n454, B2 => n1158, C1 => n455, C2 => n1159
                           , A => n1398, ZN => n1393);
   U1116 : AOI22_X1 port map( A1 => n1161, A2 => REGISTERS_27_12_port, B1 => 
                           n1162, B2 => REGISTERS_26_12_port, ZN => n1398);
   U1117 : INV_X1 port map( A => REGISTERS_24_12_port, ZN => n455);
   U1118 : INV_X1 port map( A => REGISTERS_25_12_port, ZN => n454);
   U1119 : OAI221_X1 port map( B1 => n457, B2 => n1163, C1 => n458, C2 => n1164
                           , A => n1399, ZN => n1392);
   U1120 : AOI22_X1 port map( A1 => n1166, A2 => REGISTERS_29_12_port, B1 => 
                           n1167, B2 => REGISTERS_28_12_port, ZN => n1399);
   U1121 : INV_X1 port map( A => REGISTERS_30_12_port, ZN => n458);
   U1122 : INV_X1 port map( A => REGISTERS_31_12_port, ZN => n457);
   U1123 : NOR4_X1 port map( A1 => n1400, A2 => n1401, A3 => n1402, A4 => n1403
                           , ZN => n1390);
   U1125 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_3_12_port, B1 => 
                           n1176, B2 => REGISTERS_2_12_port, ZN => n1404);
   U1126 : INV_X1 port map( A => REGISTERS_1_12_port, ZN => n464);
   U1127 : OAI221_X1 port map( B1 => n467, B2 => n1177, C1 => n468, C2 => n1178
                           , A => n1405, ZN => n1402);
   U1128 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_7_12_port, B1 => 
                           n1181, B2 => REGISTERS_6_12_port, ZN => n1405);
   U1129 : INV_X1 port map( A => REGISTERS_4_12_port, ZN => n468);
   U1130 : INV_X1 port map( A => REGISTERS_5_12_port, ZN => n467);
   U1131 : OAI221_X1 port map( B1 => n470, B2 => n1182, C1 => n471, C2 => n1183
                           , A => n1406, ZN => n1401);
   U1132 : AOI22_X1 port map( A1 => n1185, A2 => REGISTERS_11_12_port, B1 => 
                           n1186, B2 => REGISTERS_10_12_port, ZN => n1406);
   U1133 : INV_X1 port map( A => REGISTERS_8_12_port, ZN => n471);
   U1134 : INV_X1 port map( A => REGISTERS_9_12_port, ZN => n470);
   U1135 : OAI221_X1 port map( B1 => n473, B2 => n1187, C1 => n474, C2 => n1188
                           , A => n1407, ZN => n1400);
   U1136 : AOI22_X1 port map( A1 => n1190, A2 => REGISTERS_15_12_port, B1 => 
                           n1191, B2 => REGISTERS_14_12_port, ZN => n1407);
   U1137 : INV_X1 port map( A => REGISTERS_12_12_port, ZN => n474);
   U1138 : INV_X1 port map( A => REGISTERS_13_12_port, ZN => n473);
   U1139 : NAND2_X1 port map( A1 => n1408, A2 => n1409, ZN => N4233);
   U1140 : NOR4_X1 port map( A1 => n1410, A2 => n1411, A3 => n1412, A4 => n1413
                           , ZN => n1409);
   U1141 : OAI221_X1 port map( B1 => n482, B2 => n1148, C1 => n483, C2 => n1149
                           , A => n1414, ZN => n1413);
   U1142 : AOI22_X1 port map( A1 => n1151, A2 => REGISTERS_19_13_port, B1 => 
                           n1152, B2 => REGISTERS_18_13_port, ZN => n1414);
   U1143 : INV_X1 port map( A => REGISTERS_16_13_port, ZN => n483);
   U1144 : INV_X1 port map( A => REGISTERS_17_13_port, ZN => n482);
   U1145 : OAI221_X1 port map( B1 => n485, B2 => n1153, C1 => n486, C2 => n1154
                           , A => n1415, ZN => n1412);
   U1146 : AOI22_X1 port map( A1 => n1156, A2 => REGISTERS_23_13_port, B1 => 
                           n1157, B2 => REGISTERS_22_13_port, ZN => n1415);
   U1147 : INV_X1 port map( A => REGISTERS_20_13_port, ZN => n486);
   U1148 : INV_X1 port map( A => REGISTERS_21_13_port, ZN => n485);
   U1149 : OAI221_X1 port map( B1 => n488, B2 => n1158, C1 => n489, C2 => n1159
                           , A => n1416, ZN => n1411);
   U1150 : AOI22_X1 port map( A1 => n1161, A2 => REGISTERS_27_13_port, B1 => 
                           n1162, B2 => REGISTERS_26_13_port, ZN => n1416);
   U1151 : INV_X1 port map( A => REGISTERS_24_13_port, ZN => n489);
   U1152 : INV_X1 port map( A => REGISTERS_25_13_port, ZN => n488);
   U1153 : OAI221_X1 port map( B1 => n491, B2 => n1163, C1 => n492, C2 => n1164
                           , A => n1417, ZN => n1410);
   U1154 : AOI22_X1 port map( A1 => n1166, A2 => REGISTERS_29_13_port, B1 => 
                           n1167, B2 => REGISTERS_28_13_port, ZN => n1417);
   U1155 : INV_X1 port map( A => REGISTERS_30_13_port, ZN => n492);
   U1156 : INV_X1 port map( A => REGISTERS_31_13_port, ZN => n491);
   U1157 : NOR4_X1 port map( A1 => n1418, A2 => n1419, A3 => n1420, A4 => n1421
                           , ZN => n1408);
   U1159 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_3_13_port, B1 => 
                           n1176, B2 => REGISTERS_2_13_port, ZN => n1422);
   U1160 : INV_X1 port map( A => REGISTERS_1_13_port, ZN => n498);
   U1161 : OAI221_X1 port map( B1 => n501, B2 => n1177, C1 => n502, C2 => n1178
                           , A => n1423, ZN => n1420);
   U1162 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_7_13_port, B1 => 
                           n1181, B2 => REGISTERS_6_13_port, ZN => n1423);
   U1163 : INV_X1 port map( A => REGISTERS_4_13_port, ZN => n502);
   U1164 : INV_X1 port map( A => REGISTERS_5_13_port, ZN => n501);
   U1165 : OAI221_X1 port map( B1 => n504, B2 => n1182, C1 => n505, C2 => n1183
                           , A => n1424, ZN => n1419);
   U1166 : AOI22_X1 port map( A1 => n1185, A2 => REGISTERS_11_13_port, B1 => 
                           n1186, B2 => REGISTERS_10_13_port, ZN => n1424);
   U1167 : INV_X1 port map( A => REGISTERS_8_13_port, ZN => n505);
   U1168 : INV_X1 port map( A => REGISTERS_9_13_port, ZN => n504);
   U1169 : OAI221_X1 port map( B1 => n507, B2 => n1187, C1 => n508, C2 => n1188
                           , A => n1425, ZN => n1418);
   U1170 : AOI22_X1 port map( A1 => n1190, A2 => REGISTERS_15_13_port, B1 => 
                           n1191, B2 => REGISTERS_14_13_port, ZN => n1425);
   U1171 : INV_X1 port map( A => REGISTERS_12_13_port, ZN => n508);
   U1172 : INV_X1 port map( A => REGISTERS_13_13_port, ZN => n507);
   U1173 : NAND2_X1 port map( A1 => n1426, A2 => n1427, ZN => N4232);
   U1174 : NOR4_X1 port map( A1 => n1428, A2 => n1429, A3 => n1430, A4 => n1431
                           , ZN => n1427);
   U1175 : OAI221_X1 port map( B1 => n516, B2 => n1148, C1 => n517, C2 => n1149
                           , A => n1432, ZN => n1431);
   U1176 : AOI22_X1 port map( A1 => n1151, A2 => REGISTERS_19_14_port, B1 => 
                           n1152, B2 => REGISTERS_18_14_port, ZN => n1432);
   U1177 : INV_X1 port map( A => REGISTERS_16_14_port, ZN => n517);
   U1178 : INV_X1 port map( A => REGISTERS_17_14_port, ZN => n516);
   U1179 : OAI221_X1 port map( B1 => n519, B2 => n1153, C1 => n520, C2 => n1154
                           , A => n1433, ZN => n1430);
   U1180 : AOI22_X1 port map( A1 => n1156, A2 => REGISTERS_23_14_port, B1 => 
                           n1157, B2 => REGISTERS_22_14_port, ZN => n1433);
   U1181 : INV_X1 port map( A => REGISTERS_20_14_port, ZN => n520);
   U1182 : INV_X1 port map( A => REGISTERS_21_14_port, ZN => n519);
   U1183 : OAI221_X1 port map( B1 => n522, B2 => n1158, C1 => n523, C2 => n1159
                           , A => n1434, ZN => n1429);
   U1184 : AOI22_X1 port map( A1 => n1161, A2 => REGISTERS_27_14_port, B1 => 
                           n1162, B2 => REGISTERS_26_14_port, ZN => n1434);
   U1185 : INV_X1 port map( A => REGISTERS_24_14_port, ZN => n523);
   U1186 : INV_X1 port map( A => REGISTERS_25_14_port, ZN => n522);
   U1187 : OAI221_X1 port map( B1 => n525, B2 => n1163, C1 => n526, C2 => n1164
                           , A => n1435, ZN => n1428);
   U1188 : AOI22_X1 port map( A1 => n1166, A2 => REGISTERS_29_14_port, B1 => 
                           n1167, B2 => REGISTERS_28_14_port, ZN => n1435);
   U1189 : INV_X1 port map( A => REGISTERS_30_14_port, ZN => n526);
   U1190 : INV_X1 port map( A => REGISTERS_31_14_port, ZN => n525);
   U1191 : NOR4_X1 port map( A1 => n1436, A2 => n1437, A3 => n1438, A4 => n1439
                           , ZN => n1426);
   U1193 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_3_14_port, B1 => 
                           n1176, B2 => REGISTERS_2_14_port, ZN => n1440);
   U1194 : INV_X1 port map( A => REGISTERS_1_14_port, ZN => n532);
   U1195 : OAI221_X1 port map( B1 => n535, B2 => n1177, C1 => n536, C2 => n1178
                           , A => n1441, ZN => n1438);
   U1196 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_7_14_port, B1 => 
                           n1181, B2 => REGISTERS_6_14_port, ZN => n1441);
   U1197 : INV_X1 port map( A => REGISTERS_4_14_port, ZN => n536);
   U1198 : INV_X1 port map( A => REGISTERS_5_14_port, ZN => n535);
   U1199 : OAI221_X1 port map( B1 => n538, B2 => n1182, C1 => n539, C2 => n1183
                           , A => n1442, ZN => n1437);
   U1200 : AOI22_X1 port map( A1 => n1185, A2 => REGISTERS_11_14_port, B1 => 
                           n1186, B2 => REGISTERS_10_14_port, ZN => n1442);
   U1201 : INV_X1 port map( A => REGISTERS_8_14_port, ZN => n539);
   U1202 : INV_X1 port map( A => REGISTERS_9_14_port, ZN => n538);
   U1203 : OAI221_X1 port map( B1 => n541, B2 => n1187, C1 => n542, C2 => n1188
                           , A => n1443, ZN => n1436);
   U1204 : AOI22_X1 port map( A1 => n1190, A2 => REGISTERS_15_14_port, B1 => 
                           n1191, B2 => REGISTERS_14_14_port, ZN => n1443);
   U1205 : INV_X1 port map( A => REGISTERS_12_14_port, ZN => n542);
   U1206 : INV_X1 port map( A => REGISTERS_13_14_port, ZN => n541);
   U1207 : NAND2_X1 port map( A1 => n1444, A2 => n1445, ZN => N4231);
   U1208 : NOR4_X1 port map( A1 => n1446, A2 => n1447, A3 => n1448, A4 => n1449
                           , ZN => n1445);
   U1209 : OAI221_X1 port map( B1 => n550, B2 => n1148, C1 => n551, C2 => n1149
                           , A => n1450, ZN => n1449);
   U1210 : AOI22_X1 port map( A1 => n1151, A2 => REGISTERS_19_15_port, B1 => 
                           n1152, B2 => REGISTERS_18_15_port, ZN => n1450);
   U1211 : INV_X1 port map( A => REGISTERS_16_15_port, ZN => n551);
   U1212 : INV_X1 port map( A => REGISTERS_17_15_port, ZN => n550);
   U1213 : OAI221_X1 port map( B1 => n553, B2 => n1153, C1 => n554, C2 => n1154
                           , A => n1451, ZN => n1448);
   U1214 : AOI22_X1 port map( A1 => n1156, A2 => REGISTERS_23_15_port, B1 => 
                           n1157, B2 => REGISTERS_22_15_port, ZN => n1451);
   U1215 : INV_X1 port map( A => REGISTERS_20_15_port, ZN => n554);
   U1216 : INV_X1 port map( A => REGISTERS_21_15_port, ZN => n553);
   U1217 : OAI221_X1 port map( B1 => n556, B2 => n1158, C1 => n557, C2 => n1159
                           , A => n1452, ZN => n1447);
   U1218 : AOI22_X1 port map( A1 => n1161, A2 => REGISTERS_27_15_port, B1 => 
                           n1162, B2 => REGISTERS_26_15_port, ZN => n1452);
   U1219 : INV_X1 port map( A => REGISTERS_24_15_port, ZN => n557);
   U1220 : INV_X1 port map( A => REGISTERS_25_15_port, ZN => n556);
   U1221 : OAI221_X1 port map( B1 => n559, B2 => n1163, C1 => n560, C2 => n1164
                           , A => n1453, ZN => n1446);
   U1222 : AOI22_X1 port map( A1 => n1166, A2 => REGISTERS_29_15_port, B1 => 
                           n1167, B2 => REGISTERS_28_15_port, ZN => n1453);
   U1223 : INV_X1 port map( A => REGISTERS_30_15_port, ZN => n560);
   U1224 : INV_X1 port map( A => REGISTERS_31_15_port, ZN => n559);
   U1225 : NOR4_X1 port map( A1 => n1454, A2 => n1455, A3 => n1456, A4 => n1457
                           , ZN => n1444);
   U1227 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_3_15_port, B1 => 
                           n1176, B2 => REGISTERS_2_15_port, ZN => n1458);
   U1228 : INV_X1 port map( A => REGISTERS_1_15_port, ZN => n566);
   U1229 : OAI221_X1 port map( B1 => n569, B2 => n1177, C1 => n570, C2 => n1178
                           , A => n1459, ZN => n1456);
   U1230 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_7_15_port, B1 => 
                           n1181, B2 => REGISTERS_6_15_port, ZN => n1459);
   U1231 : INV_X1 port map( A => REGISTERS_4_15_port, ZN => n570);
   U1232 : INV_X1 port map( A => REGISTERS_5_15_port, ZN => n569);
   U1233 : OAI221_X1 port map( B1 => n572, B2 => n1182, C1 => n573, C2 => n1183
                           , A => n1460, ZN => n1455);
   U1234 : AOI22_X1 port map( A1 => n1185, A2 => REGISTERS_11_15_port, B1 => 
                           n1186, B2 => REGISTERS_10_15_port, ZN => n1460);
   U1235 : INV_X1 port map( A => REGISTERS_8_15_port, ZN => n573);
   U1236 : INV_X1 port map( A => REGISTERS_9_15_port, ZN => n572);
   U1237 : OAI221_X1 port map( B1 => n575, B2 => n1187, C1 => n576, C2 => n1188
                           , A => n1461, ZN => n1454);
   U1238 : AOI22_X1 port map( A1 => n1190, A2 => REGISTERS_15_15_port, B1 => 
                           n1191, B2 => REGISTERS_14_15_port, ZN => n1461);
   U1239 : INV_X1 port map( A => REGISTERS_12_15_port, ZN => n576);
   U1240 : INV_X1 port map( A => REGISTERS_13_15_port, ZN => n575);
   U1241 : NAND2_X1 port map( A1 => n1462, A2 => n1463, ZN => N4230);
   U1242 : NOR4_X1 port map( A1 => n1464, A2 => n1465, A3 => n1466, A4 => n1467
                           , ZN => n1463);
   U1243 : OAI221_X1 port map( B1 => n584, B2 => n1148, C1 => n585, C2 => n1149
                           , A => n1468, ZN => n1467);
   U1244 : AOI22_X1 port map( A1 => n1151, A2 => REGISTERS_19_16_port, B1 => 
                           n1152, B2 => REGISTERS_18_16_port, ZN => n1468);
   U1245 : INV_X1 port map( A => REGISTERS_16_16_port, ZN => n585);
   U1246 : INV_X1 port map( A => REGISTERS_17_16_port, ZN => n584);
   U1247 : OAI221_X1 port map( B1 => n587, B2 => n1153, C1 => n588, C2 => n1154
                           , A => n1469, ZN => n1466);
   U1248 : AOI22_X1 port map( A1 => n1156, A2 => REGISTERS_23_16_port, B1 => 
                           n1157, B2 => REGISTERS_22_16_port, ZN => n1469);
   U1249 : INV_X1 port map( A => REGISTERS_20_16_port, ZN => n588);
   U1250 : INV_X1 port map( A => REGISTERS_21_16_port, ZN => n587);
   U1251 : OAI221_X1 port map( B1 => n590, B2 => n1158, C1 => n591, C2 => n1159
                           , A => n1470, ZN => n1465);
   U1252 : AOI22_X1 port map( A1 => n1161, A2 => REGISTERS_27_16_port, B1 => 
                           n1162, B2 => REGISTERS_26_16_port, ZN => n1470);
   U1253 : INV_X1 port map( A => REGISTERS_24_16_port, ZN => n591);
   U1254 : INV_X1 port map( A => REGISTERS_25_16_port, ZN => n590);
   U1255 : OAI221_X1 port map( B1 => n593, B2 => n1163, C1 => n594, C2 => n1164
                           , A => n1471, ZN => n1464);
   U1256 : AOI22_X1 port map( A1 => n1166, A2 => REGISTERS_29_16_port, B1 => 
                           n1167, B2 => REGISTERS_28_16_port, ZN => n1471);
   U1257 : INV_X1 port map( A => REGISTERS_30_16_port, ZN => n594);
   U1258 : INV_X1 port map( A => REGISTERS_31_16_port, ZN => n593);
   U1259 : NOR4_X1 port map( A1 => n1472, A2 => n1473, A3 => n1474, A4 => n1475
                           , ZN => n1462);
   U1261 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_3_16_port, B1 => 
                           n1176, B2 => REGISTERS_2_16_port, ZN => n1476);
   U1262 : INV_X1 port map( A => REGISTERS_1_16_port, ZN => n600);
   U1263 : OAI221_X1 port map( B1 => n603, B2 => n1177, C1 => n604, C2 => n1178
                           , A => n1477, ZN => n1474);
   U1264 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_7_16_port, B1 => 
                           n1181, B2 => REGISTERS_6_16_port, ZN => n1477);
   U1265 : INV_X1 port map( A => REGISTERS_4_16_port, ZN => n604);
   U1266 : INV_X1 port map( A => REGISTERS_5_16_port, ZN => n603);
   U1267 : OAI221_X1 port map( B1 => n606, B2 => n1182, C1 => n607, C2 => n1183
                           , A => n1478, ZN => n1473);
   U1268 : AOI22_X1 port map( A1 => n1185, A2 => REGISTERS_11_16_port, B1 => 
                           n1186, B2 => REGISTERS_10_16_port, ZN => n1478);
   U1269 : INV_X1 port map( A => REGISTERS_8_16_port, ZN => n607);
   U1270 : INV_X1 port map( A => REGISTERS_9_16_port, ZN => n606);
   U1271 : OAI221_X1 port map( B1 => n609, B2 => n1187, C1 => n610, C2 => n1188
                           , A => n1479, ZN => n1472);
   U1272 : AOI22_X1 port map( A1 => n1190, A2 => REGISTERS_15_16_port, B1 => 
                           n1191, B2 => REGISTERS_14_16_port, ZN => n1479);
   U1273 : INV_X1 port map( A => REGISTERS_12_16_port, ZN => n610);
   U1274 : INV_X1 port map( A => REGISTERS_13_16_port, ZN => n609);
   U1275 : NAND2_X1 port map( A1 => n1480, A2 => n1481, ZN => N4229);
   U1276 : NOR4_X1 port map( A1 => n1482, A2 => n1483, A3 => n1484, A4 => n1485
                           , ZN => n1481);
   U1277 : OAI221_X1 port map( B1 => n618, B2 => n1148, C1 => n619, C2 => n1149
                           , A => n1486, ZN => n1485);
   U1278 : AOI22_X1 port map( A1 => n1151, A2 => REGISTERS_19_17_port, B1 => 
                           n1152, B2 => REGISTERS_18_17_port, ZN => n1486);
   U1279 : INV_X1 port map( A => REGISTERS_16_17_port, ZN => n619);
   U1280 : INV_X1 port map( A => REGISTERS_17_17_port, ZN => n618);
   U1281 : OAI221_X1 port map( B1 => n621, B2 => n1153, C1 => n622, C2 => n1154
                           , A => n1487, ZN => n1484);
   U1282 : AOI22_X1 port map( A1 => n1156, A2 => REGISTERS_23_17_port, B1 => 
                           n1157, B2 => REGISTERS_22_17_port, ZN => n1487);
   U1283 : INV_X1 port map( A => REGISTERS_20_17_port, ZN => n622);
   U1284 : INV_X1 port map( A => REGISTERS_21_17_port, ZN => n621);
   U1285 : OAI221_X1 port map( B1 => n624, B2 => n1158, C1 => n625, C2 => n1159
                           , A => n1488, ZN => n1483);
   U1286 : AOI22_X1 port map( A1 => n1161, A2 => REGISTERS_27_17_port, B1 => 
                           n1162, B2 => REGISTERS_26_17_port, ZN => n1488);
   U1287 : INV_X1 port map( A => REGISTERS_24_17_port, ZN => n625);
   U1288 : INV_X1 port map( A => REGISTERS_25_17_port, ZN => n624);
   U1289 : OAI221_X1 port map( B1 => n627, B2 => n1163, C1 => n628, C2 => n1164
                           , A => n1489, ZN => n1482);
   U1290 : AOI22_X1 port map( A1 => n1166, A2 => REGISTERS_29_17_port, B1 => 
                           n1167, B2 => REGISTERS_28_17_port, ZN => n1489);
   U1291 : INV_X1 port map( A => REGISTERS_30_17_port, ZN => n628);
   U1292 : INV_X1 port map( A => REGISTERS_31_17_port, ZN => n627);
   U1293 : NOR4_X1 port map( A1 => n1490, A2 => n1491, A3 => n1492, A4 => n1493
                           , ZN => n1480);
   U1295 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_3_17_port, B1 => 
                           n1176, B2 => REGISTERS_2_17_port, ZN => n1494);
   U1296 : INV_X1 port map( A => REGISTERS_1_17_port, ZN => n634);
   U1297 : OAI221_X1 port map( B1 => n637, B2 => n1177, C1 => n638, C2 => n1178
                           , A => n1495, ZN => n1492);
   U1298 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_7_17_port, B1 => 
                           n1181, B2 => REGISTERS_6_17_port, ZN => n1495);
   U1299 : INV_X1 port map( A => REGISTERS_4_17_port, ZN => n638);
   U1300 : INV_X1 port map( A => REGISTERS_5_17_port, ZN => n637);
   U1301 : OAI221_X1 port map( B1 => n640, B2 => n1182, C1 => n641, C2 => n1183
                           , A => n1496, ZN => n1491);
   U1302 : AOI22_X1 port map( A1 => n1185, A2 => REGISTERS_11_17_port, B1 => 
                           n1186, B2 => REGISTERS_10_17_port, ZN => n1496);
   U1303 : INV_X1 port map( A => REGISTERS_8_17_port, ZN => n641);
   U1304 : INV_X1 port map( A => REGISTERS_9_17_port, ZN => n640);
   U1305 : OAI221_X1 port map( B1 => n643, B2 => n1187, C1 => n644, C2 => n1188
                           , A => n1497, ZN => n1490);
   U1306 : AOI22_X1 port map( A1 => n1190, A2 => REGISTERS_15_17_port, B1 => 
                           n1191, B2 => REGISTERS_14_17_port, ZN => n1497);
   U1307 : INV_X1 port map( A => REGISTERS_12_17_port, ZN => n644);
   U1308 : INV_X1 port map( A => REGISTERS_13_17_port, ZN => n643);
   U1309 : NAND2_X1 port map( A1 => n1498, A2 => n1499, ZN => N4228);
   U1310 : NOR4_X1 port map( A1 => n1500, A2 => n1501, A3 => n1502, A4 => n1503
                           , ZN => n1499);
   U1311 : OAI221_X1 port map( B1 => n652, B2 => n1148, C1 => n653, C2 => n1149
                           , A => n1504, ZN => n1503);
   U1312 : AOI22_X1 port map( A1 => n1151, A2 => REGISTERS_19_18_port, B1 => 
                           n1152, B2 => REGISTERS_18_18_port, ZN => n1504);
   U1313 : INV_X1 port map( A => REGISTERS_16_18_port, ZN => n653);
   U1314 : INV_X1 port map( A => REGISTERS_17_18_port, ZN => n652);
   U1315 : OAI221_X1 port map( B1 => n655, B2 => n1153, C1 => n656, C2 => n1154
                           , A => n1505, ZN => n1502);
   U1316 : AOI22_X1 port map( A1 => n1156, A2 => REGISTERS_23_18_port, B1 => 
                           n1157, B2 => REGISTERS_22_18_port, ZN => n1505);
   U1317 : INV_X1 port map( A => REGISTERS_20_18_port, ZN => n656);
   U1318 : INV_X1 port map( A => REGISTERS_21_18_port, ZN => n655);
   U1319 : OAI221_X1 port map( B1 => n658, B2 => n1158, C1 => n659, C2 => n1159
                           , A => n1506, ZN => n1501);
   U1320 : AOI22_X1 port map( A1 => n1161, A2 => REGISTERS_27_18_port, B1 => 
                           n1162, B2 => REGISTERS_26_18_port, ZN => n1506);
   U1321 : INV_X1 port map( A => REGISTERS_24_18_port, ZN => n659);
   U1322 : INV_X1 port map( A => REGISTERS_25_18_port, ZN => n658);
   U1323 : OAI221_X1 port map( B1 => n661, B2 => n1163, C1 => n662, C2 => n1164
                           , A => n1507, ZN => n1500);
   U1324 : AOI22_X1 port map( A1 => n1166, A2 => REGISTERS_29_18_port, B1 => 
                           n1167, B2 => REGISTERS_28_18_port, ZN => n1507);
   U1325 : INV_X1 port map( A => REGISTERS_30_18_port, ZN => n662);
   U1326 : INV_X1 port map( A => REGISTERS_31_18_port, ZN => n661);
   U1327 : NOR4_X1 port map( A1 => n1508, A2 => n1509, A3 => n1510, A4 => n1511
                           , ZN => n1498);
   U1329 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_3_18_port, B1 => 
                           n1176, B2 => REGISTERS_2_18_port, ZN => n1512);
   U1330 : INV_X1 port map( A => REGISTERS_1_18_port, ZN => n668);
   U1331 : OAI221_X1 port map( B1 => n671, B2 => n1177, C1 => n672, C2 => n1178
                           , A => n1513, ZN => n1510);
   U1332 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_7_18_port, B1 => 
                           n1181, B2 => REGISTERS_6_18_port, ZN => n1513);
   U1333 : INV_X1 port map( A => REGISTERS_4_18_port, ZN => n672);
   U1334 : INV_X1 port map( A => REGISTERS_5_18_port, ZN => n671);
   U1335 : OAI221_X1 port map( B1 => n674, B2 => n1182, C1 => n675, C2 => n1183
                           , A => n1514, ZN => n1509);
   U1336 : AOI22_X1 port map( A1 => n1185, A2 => REGISTERS_11_18_port, B1 => 
                           n1186, B2 => REGISTERS_10_18_port, ZN => n1514);
   U1337 : INV_X1 port map( A => REGISTERS_8_18_port, ZN => n675);
   U1338 : INV_X1 port map( A => REGISTERS_9_18_port, ZN => n674);
   U1339 : OAI221_X1 port map( B1 => n677, B2 => n1187, C1 => n678, C2 => n1188
                           , A => n1515, ZN => n1508);
   U1340 : AOI22_X1 port map( A1 => n1190, A2 => REGISTERS_15_18_port, B1 => 
                           n1191, B2 => REGISTERS_14_18_port, ZN => n1515);
   U1341 : INV_X1 port map( A => REGISTERS_12_18_port, ZN => n678);
   U1342 : INV_X1 port map( A => REGISTERS_13_18_port, ZN => n677);
   U1343 : NAND2_X1 port map( A1 => n1516, A2 => n1517, ZN => N4227);
   U1344 : NOR4_X1 port map( A1 => n1518, A2 => n1519, A3 => n1520, A4 => n1521
                           , ZN => n1517);
   U1345 : OAI221_X1 port map( B1 => n686, B2 => n1148, C1 => n687, C2 => n1149
                           , A => n1522, ZN => n1521);
   U1346 : AOI22_X1 port map( A1 => n1151, A2 => REGISTERS_19_19_port, B1 => 
                           n1152, B2 => REGISTERS_18_19_port, ZN => n1522);
   U1347 : INV_X1 port map( A => REGISTERS_16_19_port, ZN => n687);
   U1348 : INV_X1 port map( A => REGISTERS_17_19_port, ZN => n686);
   U1349 : OAI221_X1 port map( B1 => n689, B2 => n1153, C1 => n690, C2 => n1154
                           , A => n1523, ZN => n1520);
   U1350 : AOI22_X1 port map( A1 => n1156, A2 => REGISTERS_23_19_port, B1 => 
                           n1157, B2 => REGISTERS_22_19_port, ZN => n1523);
   U1351 : INV_X1 port map( A => REGISTERS_20_19_port, ZN => n690);
   U1352 : INV_X1 port map( A => REGISTERS_21_19_port, ZN => n689);
   U1353 : OAI221_X1 port map( B1 => n692, B2 => n1158, C1 => n693, C2 => n1159
                           , A => n1524, ZN => n1519);
   U1354 : AOI22_X1 port map( A1 => n1161, A2 => REGISTERS_27_19_port, B1 => 
                           n1162, B2 => REGISTERS_26_19_port, ZN => n1524);
   U1355 : INV_X1 port map( A => REGISTERS_24_19_port, ZN => n693);
   U1356 : INV_X1 port map( A => REGISTERS_25_19_port, ZN => n692);
   U1357 : OAI221_X1 port map( B1 => n695, B2 => n1163, C1 => n696, C2 => n1164
                           , A => n1525, ZN => n1518);
   U1358 : AOI22_X1 port map( A1 => n1166, A2 => REGISTERS_29_19_port, B1 => 
                           n1167, B2 => REGISTERS_28_19_port, ZN => n1525);
   U1359 : INV_X1 port map( A => REGISTERS_30_19_port, ZN => n696);
   U1360 : INV_X1 port map( A => REGISTERS_31_19_port, ZN => n695);
   U1361 : NOR4_X1 port map( A1 => n1526, A2 => n1527, A3 => n1528, A4 => n1529
                           , ZN => n1516);
   U1363 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_3_19_port, B1 => 
                           n1176, B2 => REGISTERS_2_19_port, ZN => n1530);
   U1364 : INV_X1 port map( A => REGISTERS_1_19_port, ZN => n702);
   U1365 : OAI221_X1 port map( B1 => n705, B2 => n1177, C1 => n706, C2 => n1178
                           , A => n1531, ZN => n1528);
   U1366 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_7_19_port, B1 => 
                           n1181, B2 => REGISTERS_6_19_port, ZN => n1531);
   U1367 : INV_X1 port map( A => REGISTERS_4_19_port, ZN => n706);
   U1368 : INV_X1 port map( A => REGISTERS_5_19_port, ZN => n705);
   U1369 : OAI221_X1 port map( B1 => n708, B2 => n1182, C1 => n709, C2 => n1183
                           , A => n1532, ZN => n1527);
   U1370 : AOI22_X1 port map( A1 => n1185, A2 => REGISTERS_11_19_port, B1 => 
                           n1186, B2 => REGISTERS_10_19_port, ZN => n1532);
   U1371 : INV_X1 port map( A => REGISTERS_8_19_port, ZN => n709);
   U1372 : INV_X1 port map( A => REGISTERS_9_19_port, ZN => n708);
   U1373 : OAI221_X1 port map( B1 => n711, B2 => n1187, C1 => n712, C2 => n1188
                           , A => n1533, ZN => n1526);
   U1374 : AOI22_X1 port map( A1 => n1190, A2 => REGISTERS_15_19_port, B1 => 
                           n1191, B2 => REGISTERS_14_19_port, ZN => n1533);
   U1375 : INV_X1 port map( A => REGISTERS_12_19_port, ZN => n712);
   U1376 : INV_X1 port map( A => REGISTERS_13_19_port, ZN => n711);
   U1377 : NAND2_X1 port map( A1 => n1534, A2 => n1535, ZN => N4226);
   U1378 : NOR4_X1 port map( A1 => n1536, A2 => n1537, A3 => n1538, A4 => n1539
                           , ZN => n1535);
   U1379 : OAI221_X1 port map( B1 => n720, B2 => n1148, C1 => n721, C2 => n1149
                           , A => n1540, ZN => n1539);
   U1380 : AOI22_X1 port map( A1 => n1151, A2 => REGISTERS_19_20_port, B1 => 
                           n1152, B2 => REGISTERS_18_20_port, ZN => n1540);
   U1381 : INV_X1 port map( A => REGISTERS_16_20_port, ZN => n721);
   U1382 : INV_X1 port map( A => REGISTERS_17_20_port, ZN => n720);
   U1383 : OAI221_X1 port map( B1 => n723, B2 => n1153, C1 => n724, C2 => n1154
                           , A => n1541, ZN => n1538);
   U1384 : AOI22_X1 port map( A1 => n1156, A2 => REGISTERS_23_20_port, B1 => 
                           n1157, B2 => REGISTERS_22_20_port, ZN => n1541);
   U1385 : INV_X1 port map( A => REGISTERS_20_20_port, ZN => n724);
   U1386 : INV_X1 port map( A => REGISTERS_21_20_port, ZN => n723);
   U1387 : OAI221_X1 port map( B1 => n726, B2 => n1158, C1 => n727, C2 => n1159
                           , A => n1542, ZN => n1537);
   U1388 : AOI22_X1 port map( A1 => n1161, A2 => REGISTERS_27_20_port, B1 => 
                           n1162, B2 => REGISTERS_26_20_port, ZN => n1542);
   U1389 : INV_X1 port map( A => REGISTERS_24_20_port, ZN => n727);
   U1390 : INV_X1 port map( A => REGISTERS_25_20_port, ZN => n726);
   U1391 : OAI221_X1 port map( B1 => n729, B2 => n1163, C1 => n730, C2 => n1164
                           , A => n1543, ZN => n1536);
   U1392 : AOI22_X1 port map( A1 => n1166, A2 => REGISTERS_29_20_port, B1 => 
                           n1167, B2 => REGISTERS_28_20_port, ZN => n1543);
   U1393 : INV_X1 port map( A => REGISTERS_30_20_port, ZN => n730);
   U1394 : INV_X1 port map( A => REGISTERS_31_20_port, ZN => n729);
   U1395 : NOR4_X1 port map( A1 => n1544, A2 => n1545, A3 => n1546, A4 => n1547
                           , ZN => n1534);
   U1397 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_3_20_port, B1 => 
                           n1176, B2 => REGISTERS_2_20_port, ZN => n1548);
   U1398 : INV_X1 port map( A => REGISTERS_1_20_port, ZN => n736);
   U1399 : OAI221_X1 port map( B1 => n739, B2 => n1177, C1 => n740, C2 => n1178
                           , A => n1549, ZN => n1546);
   U1400 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_7_20_port, B1 => 
                           n1181, B2 => REGISTERS_6_20_port, ZN => n1549);
   U1401 : INV_X1 port map( A => REGISTERS_4_20_port, ZN => n740);
   U1402 : INV_X1 port map( A => REGISTERS_5_20_port, ZN => n739);
   U1403 : OAI221_X1 port map( B1 => n742, B2 => n1182, C1 => n743, C2 => n1183
                           , A => n1550, ZN => n1545);
   U1404 : AOI22_X1 port map( A1 => n1185, A2 => REGISTERS_11_20_port, B1 => 
                           n1186, B2 => REGISTERS_10_20_port, ZN => n1550);
   U1405 : INV_X1 port map( A => REGISTERS_8_20_port, ZN => n743);
   U1406 : INV_X1 port map( A => REGISTERS_9_20_port, ZN => n742);
   U1407 : OAI221_X1 port map( B1 => n745, B2 => n1187, C1 => n746, C2 => n1188
                           , A => n1551, ZN => n1544);
   U1408 : AOI22_X1 port map( A1 => n1190, A2 => REGISTERS_15_20_port, B1 => 
                           n1191, B2 => REGISTERS_14_20_port, ZN => n1551);
   U1409 : INV_X1 port map( A => REGISTERS_12_20_port, ZN => n746);
   U1410 : INV_X1 port map( A => REGISTERS_13_20_port, ZN => n745);
   U1411 : NAND2_X1 port map( A1 => n1552, A2 => n1553, ZN => N4225);
   U1412 : NOR4_X1 port map( A1 => n1554, A2 => n1555, A3 => n1556, A4 => n1557
                           , ZN => n1553);
   U1413 : OAI221_X1 port map( B1 => n754, B2 => n1148, C1 => n755, C2 => n1149
                           , A => n1558, ZN => n1557);
   U1414 : AOI22_X1 port map( A1 => n1151, A2 => REGISTERS_19_21_port, B1 => 
                           n1152, B2 => REGISTERS_18_21_port, ZN => n1558);
   U1415 : INV_X1 port map( A => REGISTERS_16_21_port, ZN => n755);
   U1416 : INV_X1 port map( A => REGISTERS_17_21_port, ZN => n754);
   U1417 : OAI221_X1 port map( B1 => n757, B2 => n1153, C1 => n758, C2 => n1154
                           , A => n1559, ZN => n1556);
   U1418 : AOI22_X1 port map( A1 => n1156, A2 => REGISTERS_23_21_port, B1 => 
                           n1157, B2 => REGISTERS_22_21_port, ZN => n1559);
   U1419 : INV_X1 port map( A => REGISTERS_20_21_port, ZN => n758);
   U1420 : INV_X1 port map( A => REGISTERS_21_21_port, ZN => n757);
   U1421 : OAI221_X1 port map( B1 => n760, B2 => n1158, C1 => n761, C2 => n1159
                           , A => n1560, ZN => n1555);
   U1422 : AOI22_X1 port map( A1 => n1161, A2 => REGISTERS_27_21_port, B1 => 
                           n1162, B2 => REGISTERS_26_21_port, ZN => n1560);
   U1423 : INV_X1 port map( A => REGISTERS_24_21_port, ZN => n761);
   U1424 : INV_X1 port map( A => REGISTERS_25_21_port, ZN => n760);
   U1425 : OAI221_X1 port map( B1 => n763, B2 => n1163, C1 => n764, C2 => n1164
                           , A => n1561, ZN => n1554);
   U1426 : AOI22_X1 port map( A1 => n1166, A2 => REGISTERS_29_21_port, B1 => 
                           n1167, B2 => REGISTERS_28_21_port, ZN => n1561);
   U1427 : INV_X1 port map( A => REGISTERS_30_21_port, ZN => n764);
   U1428 : INV_X1 port map( A => REGISTERS_31_21_port, ZN => n763);
   U1429 : NOR4_X1 port map( A1 => n1562, A2 => n1563, A3 => n1564, A4 => n1565
                           , ZN => n1552);
   U1431 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_3_21_port, B1 => 
                           n1176, B2 => REGISTERS_2_21_port, ZN => n1566);
   U1432 : INV_X1 port map( A => REGISTERS_1_21_port, ZN => n770);
   U1433 : OAI221_X1 port map( B1 => n773, B2 => n1177, C1 => n774, C2 => n1178
                           , A => n1567, ZN => n1564);
   U1434 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_7_21_port, B1 => 
                           n1181, B2 => REGISTERS_6_21_port, ZN => n1567);
   U1435 : INV_X1 port map( A => REGISTERS_4_21_port, ZN => n774);
   U1436 : INV_X1 port map( A => REGISTERS_5_21_port, ZN => n773);
   U1437 : OAI221_X1 port map( B1 => n776, B2 => n1182, C1 => n777, C2 => n1183
                           , A => n1568, ZN => n1563);
   U1438 : AOI22_X1 port map( A1 => n1185, A2 => REGISTERS_11_21_port, B1 => 
                           n1186, B2 => REGISTERS_10_21_port, ZN => n1568);
   U1439 : INV_X1 port map( A => REGISTERS_8_21_port, ZN => n777);
   U1440 : INV_X1 port map( A => REGISTERS_9_21_port, ZN => n776);
   U1441 : OAI221_X1 port map( B1 => n779, B2 => n1187, C1 => n780, C2 => n1188
                           , A => n1569, ZN => n1562);
   U1442 : AOI22_X1 port map( A1 => n1190, A2 => REGISTERS_15_21_port, B1 => 
                           n1191, B2 => REGISTERS_14_21_port, ZN => n1569);
   U1443 : INV_X1 port map( A => REGISTERS_12_21_port, ZN => n780);
   U1444 : INV_X1 port map( A => REGISTERS_13_21_port, ZN => n779);
   U1445 : NAND2_X1 port map( A1 => n1570, A2 => n1571, ZN => N4224);
   U1446 : NOR4_X1 port map( A1 => n1572, A2 => n1573, A3 => n1574, A4 => n1575
                           , ZN => n1571);
   U1447 : OAI221_X1 port map( B1 => n788, B2 => n1148, C1 => n789, C2 => n1149
                           , A => n1576, ZN => n1575);
   U1448 : AOI22_X1 port map( A1 => n1151, A2 => REGISTERS_19_22_port, B1 => 
                           n1152, B2 => REGISTERS_18_22_port, ZN => n1576);
   U1449 : INV_X1 port map( A => REGISTERS_16_22_port, ZN => n789);
   U1450 : INV_X1 port map( A => REGISTERS_17_22_port, ZN => n788);
   U1451 : OAI221_X1 port map( B1 => n791, B2 => n1153, C1 => n792, C2 => n1154
                           , A => n1577, ZN => n1574);
   U1452 : AOI22_X1 port map( A1 => n1156, A2 => REGISTERS_23_22_port, B1 => 
                           n1157, B2 => REGISTERS_22_22_port, ZN => n1577);
   U1453 : INV_X1 port map( A => REGISTERS_20_22_port, ZN => n792);
   U1454 : INV_X1 port map( A => REGISTERS_21_22_port, ZN => n791);
   U1455 : OAI221_X1 port map( B1 => n794, B2 => n1158, C1 => n795, C2 => n1159
                           , A => n1578, ZN => n1573);
   U1456 : AOI22_X1 port map( A1 => n1161, A2 => REGISTERS_27_22_port, B1 => 
                           n1162, B2 => REGISTERS_26_22_port, ZN => n1578);
   U1457 : INV_X1 port map( A => REGISTERS_24_22_port, ZN => n795);
   U1458 : INV_X1 port map( A => REGISTERS_25_22_port, ZN => n794);
   U1459 : OAI221_X1 port map( B1 => n797, B2 => n1163, C1 => n798, C2 => n1164
                           , A => n1579, ZN => n1572);
   U1460 : AOI22_X1 port map( A1 => n1166, A2 => REGISTERS_29_22_port, B1 => 
                           n1167, B2 => REGISTERS_28_22_port, ZN => n1579);
   U1461 : INV_X1 port map( A => REGISTERS_30_22_port, ZN => n798);
   U1462 : INV_X1 port map( A => REGISTERS_31_22_port, ZN => n797);
   U1463 : NOR4_X1 port map( A1 => n1580, A2 => n1581, A3 => n1582, A4 => n1583
                           , ZN => n1570);
   U1465 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_3_22_port, B1 => 
                           n1176, B2 => REGISTERS_2_22_port, ZN => n1584);
   U1466 : INV_X1 port map( A => REGISTERS_1_22_port, ZN => n804);
   U1467 : OAI221_X1 port map( B1 => n807, B2 => n1177, C1 => n808, C2 => n1178
                           , A => n1585, ZN => n1582);
   U1468 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_7_22_port, B1 => 
                           n1181, B2 => REGISTERS_6_22_port, ZN => n1585);
   U1469 : INV_X1 port map( A => REGISTERS_4_22_port, ZN => n808);
   U1470 : INV_X1 port map( A => REGISTERS_5_22_port, ZN => n807);
   U1471 : OAI221_X1 port map( B1 => n810, B2 => n1182, C1 => n811, C2 => n1183
                           , A => n1586, ZN => n1581);
   U1472 : AOI22_X1 port map( A1 => n1185, A2 => REGISTERS_11_22_port, B1 => 
                           n1186, B2 => REGISTERS_10_22_port, ZN => n1586);
   U1473 : INV_X1 port map( A => REGISTERS_8_22_port, ZN => n811);
   U1474 : INV_X1 port map( A => REGISTERS_9_22_port, ZN => n810);
   U1475 : OAI221_X1 port map( B1 => n813, B2 => n1187, C1 => n814, C2 => n1188
                           , A => n1587, ZN => n1580);
   U1476 : AOI22_X1 port map( A1 => n1190, A2 => REGISTERS_15_22_port, B1 => 
                           n1191, B2 => REGISTERS_14_22_port, ZN => n1587);
   U1477 : INV_X1 port map( A => REGISTERS_12_22_port, ZN => n814);
   U1478 : INV_X1 port map( A => REGISTERS_13_22_port, ZN => n813);
   U1479 : NAND2_X1 port map( A1 => n1588, A2 => n1589, ZN => N4223);
   U1480 : NOR4_X1 port map( A1 => n1590, A2 => n1591, A3 => n1592, A4 => n1593
                           , ZN => n1589);
   U1481 : OAI221_X1 port map( B1 => n822, B2 => n1148, C1 => n823, C2 => n1149
                           , A => n1594, ZN => n1593);
   U1482 : AOI22_X1 port map( A1 => n1151, A2 => REGISTERS_19_23_port, B1 => 
                           n1152, B2 => REGISTERS_18_23_port, ZN => n1594);
   U1483 : INV_X1 port map( A => REGISTERS_16_23_port, ZN => n823);
   U1484 : INV_X1 port map( A => REGISTERS_17_23_port, ZN => n822);
   U1485 : OAI221_X1 port map( B1 => n825, B2 => n1153, C1 => n826, C2 => n1154
                           , A => n1595, ZN => n1592);
   U1486 : AOI22_X1 port map( A1 => n1156, A2 => REGISTERS_23_23_port, B1 => 
                           n1157, B2 => REGISTERS_22_23_port, ZN => n1595);
   U1487 : INV_X1 port map( A => REGISTERS_20_23_port, ZN => n826);
   U1488 : INV_X1 port map( A => REGISTERS_21_23_port, ZN => n825);
   U1489 : OAI221_X1 port map( B1 => n828, B2 => n1158, C1 => n829, C2 => n1159
                           , A => n1596, ZN => n1591);
   U1490 : AOI22_X1 port map( A1 => n1161, A2 => REGISTERS_27_23_port, B1 => 
                           n1162, B2 => REGISTERS_26_23_port, ZN => n1596);
   U1491 : INV_X1 port map( A => REGISTERS_24_23_port, ZN => n829);
   U1492 : INV_X1 port map( A => REGISTERS_25_23_port, ZN => n828);
   U1493 : OAI221_X1 port map( B1 => n831, B2 => n1163, C1 => n832, C2 => n1164
                           , A => n1597, ZN => n1590);
   U1494 : AOI22_X1 port map( A1 => n1166, A2 => REGISTERS_29_23_port, B1 => 
                           n1167, B2 => REGISTERS_28_23_port, ZN => n1597);
   U1495 : INV_X1 port map( A => REGISTERS_30_23_port, ZN => n832);
   U1496 : INV_X1 port map( A => REGISTERS_31_23_port, ZN => n831);
   U1497 : NOR4_X1 port map( A1 => n1598, A2 => n1599, A3 => n1600, A4 => n1601
                           , ZN => n1588);
   U1499 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_3_23_port, B1 => 
                           n1176, B2 => REGISTERS_2_23_port, ZN => n1602);
   U1500 : INV_X1 port map( A => REGISTERS_1_23_port, ZN => n838);
   U1501 : OAI221_X1 port map( B1 => n841, B2 => n1177, C1 => n842, C2 => n1178
                           , A => n1603, ZN => n1600);
   U1502 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_7_23_port, B1 => 
                           n1181, B2 => REGISTERS_6_23_port, ZN => n1603);
   U1503 : INV_X1 port map( A => REGISTERS_4_23_port, ZN => n842);
   U1504 : INV_X1 port map( A => REGISTERS_5_23_port, ZN => n841);
   U1505 : OAI221_X1 port map( B1 => n844, B2 => n1182, C1 => n845, C2 => n1183
                           , A => n1604, ZN => n1599);
   U1506 : AOI22_X1 port map( A1 => n1185, A2 => REGISTERS_11_23_port, B1 => 
                           n1186, B2 => REGISTERS_10_23_port, ZN => n1604);
   U1507 : INV_X1 port map( A => REGISTERS_8_23_port, ZN => n845);
   U1508 : INV_X1 port map( A => REGISTERS_9_23_port, ZN => n844);
   U1509 : OAI221_X1 port map( B1 => n847, B2 => n1187, C1 => n848, C2 => n1188
                           , A => n1605, ZN => n1598);
   U1510 : AOI22_X1 port map( A1 => n1190, A2 => REGISTERS_15_23_port, B1 => 
                           n1191, B2 => REGISTERS_14_23_port, ZN => n1605);
   U1511 : INV_X1 port map( A => REGISTERS_12_23_port, ZN => n848);
   U1512 : INV_X1 port map( A => REGISTERS_13_23_port, ZN => n847);
   U1513 : NAND2_X1 port map( A1 => n1606, A2 => n1607, ZN => N4222);
   U1514 : NOR4_X1 port map( A1 => n1608, A2 => n1609, A3 => n1610, A4 => n1611
                           , ZN => n1607);
   U1515 : OAI221_X1 port map( B1 => n856, B2 => n1148, C1 => n857, C2 => n1149
                           , A => n1612, ZN => n1611);
   U1516 : AOI22_X1 port map( A1 => n1151, A2 => REGISTERS_19_24_port, B1 => 
                           n1152, B2 => REGISTERS_18_24_port, ZN => n1612);
   U1517 : INV_X1 port map( A => REGISTERS_16_24_port, ZN => n857);
   U1518 : INV_X1 port map( A => REGISTERS_17_24_port, ZN => n856);
   U1519 : OAI221_X1 port map( B1 => n859, B2 => n1153, C1 => n860, C2 => n1154
                           , A => n1613, ZN => n1610);
   U1520 : AOI22_X1 port map( A1 => n1156, A2 => REGISTERS_23_24_port, B1 => 
                           n1157, B2 => REGISTERS_22_24_port, ZN => n1613);
   U1521 : INV_X1 port map( A => REGISTERS_20_24_port, ZN => n860);
   U1522 : INV_X1 port map( A => REGISTERS_21_24_port, ZN => n859);
   U1523 : OAI221_X1 port map( B1 => n862, B2 => n1158, C1 => n863, C2 => n1159
                           , A => n1614, ZN => n1609);
   U1524 : AOI22_X1 port map( A1 => n1161, A2 => REGISTERS_27_24_port, B1 => 
                           n1162, B2 => REGISTERS_26_24_port, ZN => n1614);
   U1525 : INV_X1 port map( A => REGISTERS_24_24_port, ZN => n863);
   U1526 : INV_X1 port map( A => REGISTERS_25_24_port, ZN => n862);
   U1527 : OAI221_X1 port map( B1 => n865, B2 => n1163, C1 => n866, C2 => n1164
                           , A => n1615, ZN => n1608);
   U1528 : AOI22_X1 port map( A1 => n1166, A2 => REGISTERS_29_24_port, B1 => 
                           n1167, B2 => REGISTERS_28_24_port, ZN => n1615);
   U1529 : INV_X1 port map( A => REGISTERS_30_24_port, ZN => n866);
   U1530 : INV_X1 port map( A => REGISTERS_31_24_port, ZN => n865);
   U1531 : NOR4_X1 port map( A1 => n1616, A2 => n1617, A3 => n1618, A4 => n1619
                           , ZN => n1606);
   U1533 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_3_24_port, B1 => 
                           n1176, B2 => REGISTERS_2_24_port, ZN => n1620);
   U1534 : INV_X1 port map( A => REGISTERS_1_24_port, ZN => n872);
   U1535 : OAI221_X1 port map( B1 => n875, B2 => n1177, C1 => n876, C2 => n1178
                           , A => n1621, ZN => n1618);
   U1536 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_7_24_port, B1 => 
                           n1181, B2 => REGISTERS_6_24_port, ZN => n1621);
   U1537 : INV_X1 port map( A => REGISTERS_4_24_port, ZN => n876);
   U1538 : INV_X1 port map( A => REGISTERS_5_24_port, ZN => n875);
   U1539 : OAI221_X1 port map( B1 => n878, B2 => n1182, C1 => n879, C2 => n1183
                           , A => n1622, ZN => n1617);
   U1540 : AOI22_X1 port map( A1 => n1185, A2 => REGISTERS_11_24_port, B1 => 
                           n1186, B2 => REGISTERS_10_24_port, ZN => n1622);
   U1541 : INV_X1 port map( A => REGISTERS_8_24_port, ZN => n879);
   U1542 : INV_X1 port map( A => REGISTERS_9_24_port, ZN => n878);
   U1543 : OAI221_X1 port map( B1 => n881, B2 => n1187, C1 => n882, C2 => n1188
                           , A => n1623, ZN => n1616);
   U1544 : AOI22_X1 port map( A1 => n1190, A2 => REGISTERS_15_24_port, B1 => 
                           n1191, B2 => REGISTERS_14_24_port, ZN => n1623);
   U1545 : INV_X1 port map( A => REGISTERS_12_24_port, ZN => n882);
   U1546 : INV_X1 port map( A => REGISTERS_13_24_port, ZN => n881);
   U1547 : NAND2_X1 port map( A1 => n1624, A2 => n1625, ZN => N4221);
   U1548 : NOR4_X1 port map( A1 => n1626, A2 => n1627, A3 => n1628, A4 => n1629
                           , ZN => n1625);
   U1549 : OAI221_X1 port map( B1 => n890, B2 => n1148, C1 => n891, C2 => n1149
                           , A => n1630, ZN => n1629);
   U1550 : AOI22_X1 port map( A1 => n1151, A2 => REGISTERS_19_25_port, B1 => 
                           n1152, B2 => REGISTERS_18_25_port, ZN => n1630);
   U1551 : INV_X1 port map( A => REGISTERS_16_25_port, ZN => n891);
   U1552 : INV_X1 port map( A => REGISTERS_17_25_port, ZN => n890);
   U1553 : OAI221_X1 port map( B1 => n893, B2 => n1153, C1 => n894, C2 => n1154
                           , A => n1631, ZN => n1628);
   U1554 : AOI22_X1 port map( A1 => n1156, A2 => REGISTERS_23_25_port, B1 => 
                           n1157, B2 => REGISTERS_22_25_port, ZN => n1631);
   U1555 : INV_X1 port map( A => REGISTERS_20_25_port, ZN => n894);
   U1556 : INV_X1 port map( A => REGISTERS_21_25_port, ZN => n893);
   U1557 : OAI221_X1 port map( B1 => n896, B2 => n1158, C1 => n897, C2 => n1159
                           , A => n1632, ZN => n1627);
   U1558 : AOI22_X1 port map( A1 => n1161, A2 => REGISTERS_27_25_port, B1 => 
                           n1162, B2 => REGISTERS_26_25_port, ZN => n1632);
   U1559 : INV_X1 port map( A => REGISTERS_24_25_port, ZN => n897);
   U1560 : INV_X1 port map( A => REGISTERS_25_25_port, ZN => n896);
   U1561 : OAI221_X1 port map( B1 => n899, B2 => n1163, C1 => n900, C2 => n1164
                           , A => n1633, ZN => n1626);
   U1562 : AOI22_X1 port map( A1 => n1166, A2 => REGISTERS_29_25_port, B1 => 
                           n1167, B2 => REGISTERS_28_25_port, ZN => n1633);
   U1563 : INV_X1 port map( A => REGISTERS_30_25_port, ZN => n900);
   U1564 : INV_X1 port map( A => REGISTERS_31_25_port, ZN => n899);
   U1565 : NOR4_X1 port map( A1 => n1634, A2 => n1635, A3 => n1636, A4 => n1637
                           , ZN => n1624);
   U1567 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_3_25_port, B1 => 
                           n1176, B2 => REGISTERS_2_25_port, ZN => n1638);
   U1568 : INV_X1 port map( A => REGISTERS_1_25_port, ZN => n906);
   U1569 : OAI221_X1 port map( B1 => n909, B2 => n1177, C1 => n910, C2 => n1178
                           , A => n1639, ZN => n1636);
   U1570 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_7_25_port, B1 => 
                           n1181, B2 => REGISTERS_6_25_port, ZN => n1639);
   U1571 : INV_X1 port map( A => REGISTERS_4_25_port, ZN => n910);
   U1572 : INV_X1 port map( A => REGISTERS_5_25_port, ZN => n909);
   U1573 : OAI221_X1 port map( B1 => n912, B2 => n1182, C1 => n913, C2 => n1183
                           , A => n1640, ZN => n1635);
   U1574 : AOI22_X1 port map( A1 => n1185, A2 => REGISTERS_11_25_port, B1 => 
                           n1186, B2 => REGISTERS_10_25_port, ZN => n1640);
   U1575 : INV_X1 port map( A => REGISTERS_8_25_port, ZN => n913);
   U1576 : INV_X1 port map( A => REGISTERS_9_25_port, ZN => n912);
   U1577 : OAI221_X1 port map( B1 => n915, B2 => n1187, C1 => n916, C2 => n1188
                           , A => n1641, ZN => n1634);
   U1578 : AOI22_X1 port map( A1 => n1190, A2 => REGISTERS_15_25_port, B1 => 
                           n1191, B2 => REGISTERS_14_25_port, ZN => n1641);
   U1579 : INV_X1 port map( A => REGISTERS_12_25_port, ZN => n916);
   U1580 : INV_X1 port map( A => REGISTERS_13_25_port, ZN => n915);
   U1581 : NAND2_X1 port map( A1 => n1642, A2 => n1643, ZN => N4220);
   U1582 : NOR4_X1 port map( A1 => n1644, A2 => n1645, A3 => n1646, A4 => n1647
                           , ZN => n1643);
   U1583 : OAI221_X1 port map( B1 => n924, B2 => n1148, C1 => n925, C2 => n1149
                           , A => n1648, ZN => n1647);
   U1584 : AOI22_X1 port map( A1 => n1151, A2 => REGISTERS_19_26_port, B1 => 
                           n1152, B2 => REGISTERS_18_26_port, ZN => n1648);
   U1585 : INV_X1 port map( A => REGISTERS_16_26_port, ZN => n925);
   U1586 : INV_X1 port map( A => REGISTERS_17_26_port, ZN => n924);
   U1587 : OAI221_X1 port map( B1 => n927, B2 => n1153, C1 => n928, C2 => n1154
                           , A => n1649, ZN => n1646);
   U1588 : AOI22_X1 port map( A1 => n1156, A2 => REGISTERS_23_26_port, B1 => 
                           n1157, B2 => REGISTERS_22_26_port, ZN => n1649);
   U1589 : INV_X1 port map( A => REGISTERS_20_26_port, ZN => n928);
   U1590 : INV_X1 port map( A => REGISTERS_21_26_port, ZN => n927);
   U1591 : OAI221_X1 port map( B1 => n930, B2 => n1158, C1 => n931, C2 => n1159
                           , A => n1650, ZN => n1645);
   U1592 : AOI22_X1 port map( A1 => n1161, A2 => REGISTERS_27_26_port, B1 => 
                           n1162, B2 => REGISTERS_26_26_port, ZN => n1650);
   U1593 : INV_X1 port map( A => REGISTERS_24_26_port, ZN => n931);
   U1594 : INV_X1 port map( A => REGISTERS_25_26_port, ZN => n930);
   U1595 : OAI221_X1 port map( B1 => n933, B2 => n1163, C1 => n934, C2 => n1164
                           , A => n1651, ZN => n1644);
   U1596 : AOI22_X1 port map( A1 => n1166, A2 => REGISTERS_29_26_port, B1 => 
                           n1167, B2 => REGISTERS_28_26_port, ZN => n1651);
   U1597 : INV_X1 port map( A => REGISTERS_30_26_port, ZN => n934);
   U1598 : INV_X1 port map( A => REGISTERS_31_26_port, ZN => n933);
   U1599 : NOR4_X1 port map( A1 => n1652, A2 => n1653, A3 => n1654, A4 => n1655
                           , ZN => n1642);
   U1601 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_3_26_port, B1 => 
                           n1176, B2 => REGISTERS_2_26_port, ZN => n1656);
   U1602 : INV_X1 port map( A => REGISTERS_1_26_port, ZN => n940);
   U1603 : OAI221_X1 port map( B1 => n943, B2 => n1177, C1 => n944, C2 => n1178
                           , A => n1657, ZN => n1654);
   U1604 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_7_26_port, B1 => 
                           n1181, B2 => REGISTERS_6_26_port, ZN => n1657);
   U1605 : INV_X1 port map( A => REGISTERS_4_26_port, ZN => n944);
   U1606 : INV_X1 port map( A => REGISTERS_5_26_port, ZN => n943);
   U1607 : OAI221_X1 port map( B1 => n946, B2 => n1182, C1 => n947, C2 => n1183
                           , A => n1658, ZN => n1653);
   U1608 : AOI22_X1 port map( A1 => n1185, A2 => REGISTERS_11_26_port, B1 => 
                           n1186, B2 => REGISTERS_10_26_port, ZN => n1658);
   U1609 : INV_X1 port map( A => REGISTERS_8_26_port, ZN => n947);
   U1610 : INV_X1 port map( A => REGISTERS_9_26_port, ZN => n946);
   U1611 : OAI221_X1 port map( B1 => n949, B2 => n1187, C1 => n950, C2 => n1188
                           , A => n1659, ZN => n1652);
   U1612 : AOI22_X1 port map( A1 => n1190, A2 => REGISTERS_15_26_port, B1 => 
                           n1191, B2 => REGISTERS_14_26_port, ZN => n1659);
   U1613 : INV_X1 port map( A => REGISTERS_12_26_port, ZN => n950);
   U1614 : INV_X1 port map( A => REGISTERS_13_26_port, ZN => n949);
   U1615 : NAND2_X1 port map( A1 => n1660, A2 => n1661, ZN => N4219);
   U1616 : NOR4_X1 port map( A1 => n1662, A2 => n1663, A3 => n1664, A4 => n1665
                           , ZN => n1661);
   U1617 : OAI221_X1 port map( B1 => n958, B2 => n1148, C1 => n959, C2 => n1149
                           , A => n1666, ZN => n1665);
   U1618 : AOI22_X1 port map( A1 => n1151, A2 => REGISTERS_19_27_port, B1 => 
                           n1152, B2 => REGISTERS_18_27_port, ZN => n1666);
   U1619 : INV_X1 port map( A => REGISTERS_16_27_port, ZN => n959);
   U1620 : INV_X1 port map( A => REGISTERS_17_27_port, ZN => n958);
   U1621 : OAI221_X1 port map( B1 => n961, B2 => n1153, C1 => n962, C2 => n1154
                           , A => n1667, ZN => n1664);
   U1622 : AOI22_X1 port map( A1 => n1156, A2 => REGISTERS_23_27_port, B1 => 
                           n1157, B2 => REGISTERS_22_27_port, ZN => n1667);
   U1623 : INV_X1 port map( A => REGISTERS_20_27_port, ZN => n962);
   U1624 : INV_X1 port map( A => REGISTERS_21_27_port, ZN => n961);
   U1625 : OAI221_X1 port map( B1 => n964, B2 => n1158, C1 => n965, C2 => n1159
                           , A => n1668, ZN => n1663);
   U1626 : AOI22_X1 port map( A1 => n1161, A2 => REGISTERS_27_27_port, B1 => 
                           n1162, B2 => REGISTERS_26_27_port, ZN => n1668);
   U1627 : INV_X1 port map( A => REGISTERS_24_27_port, ZN => n965);
   U1628 : INV_X1 port map( A => REGISTERS_25_27_port, ZN => n964);
   U1629 : OAI221_X1 port map( B1 => n967, B2 => n1163, C1 => n968, C2 => n1164
                           , A => n1669, ZN => n1662);
   U1630 : AOI22_X1 port map( A1 => n1166, A2 => REGISTERS_29_27_port, B1 => 
                           n1167, B2 => REGISTERS_28_27_port, ZN => n1669);
   U1631 : INV_X1 port map( A => REGISTERS_30_27_port, ZN => n968);
   U1632 : INV_X1 port map( A => REGISTERS_31_27_port, ZN => n967);
   U1633 : NOR4_X1 port map( A1 => n1670, A2 => n1671, A3 => n1672, A4 => n1673
                           , ZN => n1660);
   U1635 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_3_27_port, B1 => 
                           n1176, B2 => REGISTERS_2_27_port, ZN => n1674);
   U1636 : INV_X1 port map( A => REGISTERS_1_27_port, ZN => n974);
   U1637 : OAI221_X1 port map( B1 => n977, B2 => n1177, C1 => n978, C2 => n1178
                           , A => n1675, ZN => n1672);
   U1638 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_7_27_port, B1 => 
                           n1181, B2 => REGISTERS_6_27_port, ZN => n1675);
   U1639 : INV_X1 port map( A => REGISTERS_4_27_port, ZN => n978);
   U1640 : INV_X1 port map( A => REGISTERS_5_27_port, ZN => n977);
   U1641 : OAI221_X1 port map( B1 => n980, B2 => n1182, C1 => n981, C2 => n1183
                           , A => n1676, ZN => n1671);
   U1642 : AOI22_X1 port map( A1 => n1185, A2 => REGISTERS_11_27_port, B1 => 
                           n1186, B2 => REGISTERS_10_27_port, ZN => n1676);
   U1643 : INV_X1 port map( A => REGISTERS_8_27_port, ZN => n981);
   U1644 : INV_X1 port map( A => REGISTERS_9_27_port, ZN => n980);
   U1645 : OAI221_X1 port map( B1 => n983, B2 => n1187, C1 => n984, C2 => n1188
                           , A => n1677, ZN => n1670);
   U1646 : AOI22_X1 port map( A1 => n1190, A2 => REGISTERS_15_27_port, B1 => 
                           n1191, B2 => REGISTERS_14_27_port, ZN => n1677);
   U1647 : INV_X1 port map( A => REGISTERS_12_27_port, ZN => n984);
   U1648 : INV_X1 port map( A => REGISTERS_13_27_port, ZN => n983);
   U1649 : NAND2_X1 port map( A1 => n1678, A2 => n1679, ZN => N4218);
   U1650 : NOR4_X1 port map( A1 => n1680, A2 => n1681, A3 => n1682, A4 => n1683
                           , ZN => n1679);
   U1651 : OAI221_X1 port map( B1 => n992, B2 => n1148, C1 => n993, C2 => n1149
                           , A => n1684, ZN => n1683);
   U1652 : AOI22_X1 port map( A1 => n1151, A2 => REGISTERS_19_28_port, B1 => 
                           n1152, B2 => REGISTERS_18_28_port, ZN => n1684);
   U1653 : INV_X1 port map( A => REGISTERS_16_28_port, ZN => n993);
   U1654 : INV_X1 port map( A => REGISTERS_17_28_port, ZN => n992);
   U1655 : OAI221_X1 port map( B1 => n995, B2 => n1153, C1 => n996, C2 => n1154
                           , A => n1685, ZN => n1682);
   U1656 : AOI22_X1 port map( A1 => n1156, A2 => REGISTERS_23_28_port, B1 => 
                           n1157, B2 => REGISTERS_22_28_port, ZN => n1685);
   U1657 : INV_X1 port map( A => REGISTERS_20_28_port, ZN => n996);
   U1658 : INV_X1 port map( A => REGISTERS_21_28_port, ZN => n995);
   U1659 : OAI221_X1 port map( B1 => n998, B2 => n1158, C1 => n999, C2 => n1159
                           , A => n1686, ZN => n1681);
   U1660 : AOI22_X1 port map( A1 => n1161, A2 => REGISTERS_27_28_port, B1 => 
                           n1162, B2 => REGISTERS_26_28_port, ZN => n1686);
   U1661 : INV_X1 port map( A => REGISTERS_24_28_port, ZN => n999);
   U1662 : INV_X1 port map( A => REGISTERS_25_28_port, ZN => n998);
   U1663 : OAI221_X1 port map( B1 => n1001, B2 => n1163, C1 => n1002, C2 => 
                           n1164, A => n1687, ZN => n1680);
   U1664 : AOI22_X1 port map( A1 => n1166, A2 => REGISTERS_29_28_port, B1 => 
                           n1167, B2 => REGISTERS_28_28_port, ZN => n1687);
   U1665 : INV_X1 port map( A => REGISTERS_30_28_port, ZN => n1002);
   U1666 : INV_X1 port map( A => REGISTERS_31_28_port, ZN => n1001);
   U1667 : NOR4_X1 port map( A1 => n1688, A2 => n1689, A3 => n1690, A4 => n1691
                           , ZN => n1678);
   U1669 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_3_28_port, B1 => 
                           n1176, B2 => REGISTERS_2_28_port, ZN => n1692);
   U1670 : INV_X1 port map( A => REGISTERS_1_28_port, ZN => n1008);
   U1671 : OAI221_X1 port map( B1 => n1011, B2 => n1177, C1 => n1012, C2 => 
                           n1178, A => n1693, ZN => n1690);
   U1672 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_7_28_port, B1 => 
                           n1181, B2 => REGISTERS_6_28_port, ZN => n1693);
   U1673 : INV_X1 port map( A => REGISTERS_4_28_port, ZN => n1012);
   U1674 : INV_X1 port map( A => REGISTERS_5_28_port, ZN => n1011);
   U1675 : OAI221_X1 port map( B1 => n1014, B2 => n1182, C1 => n1015, C2 => 
                           n1183, A => n1694, ZN => n1689);
   U1676 : AOI22_X1 port map( A1 => n1185, A2 => REGISTERS_11_28_port, B1 => 
                           n1186, B2 => REGISTERS_10_28_port, ZN => n1694);
   U1677 : INV_X1 port map( A => REGISTERS_8_28_port, ZN => n1015);
   U1678 : INV_X1 port map( A => REGISTERS_9_28_port, ZN => n1014);
   U1679 : OAI221_X1 port map( B1 => n1017, B2 => n1187, C1 => n1018, C2 => 
                           n1188, A => n1695, ZN => n1688);
   U1680 : AOI22_X1 port map( A1 => n1190, A2 => REGISTERS_15_28_port, B1 => 
                           n1191, B2 => REGISTERS_14_28_port, ZN => n1695);
   U1681 : INV_X1 port map( A => REGISTERS_12_28_port, ZN => n1018);
   U1682 : INV_X1 port map( A => REGISTERS_13_28_port, ZN => n1017);
   U1683 : NAND2_X1 port map( A1 => n1696, A2 => n1697, ZN => N4217);
   U1684 : NOR4_X1 port map( A1 => n1698, A2 => n1699, A3 => n1700, A4 => n1701
                           , ZN => n1697);
   U1685 : OAI221_X1 port map( B1 => n1026, B2 => n1148, C1 => n1027, C2 => 
                           n1149, A => n1702, ZN => n1701);
   U1686 : AOI22_X1 port map( A1 => n1151, A2 => REGISTERS_19_29_port, B1 => 
                           n1152, B2 => REGISTERS_18_29_port, ZN => n1702);
   U1687 : INV_X1 port map( A => REGISTERS_16_29_port, ZN => n1027);
   U1688 : INV_X1 port map( A => REGISTERS_17_29_port, ZN => n1026);
   U1689 : OAI221_X1 port map( B1 => n1029, B2 => n1153, C1 => n1030, C2 => 
                           n1154, A => n1703, ZN => n1700);
   U1690 : AOI22_X1 port map( A1 => n1156, A2 => REGISTERS_23_29_port, B1 => 
                           n1157, B2 => REGISTERS_22_29_port, ZN => n1703);
   U1691 : INV_X1 port map( A => REGISTERS_20_29_port, ZN => n1030);
   U1692 : INV_X1 port map( A => REGISTERS_21_29_port, ZN => n1029);
   U1693 : OAI221_X1 port map( B1 => n1032, B2 => n1158, C1 => n1033, C2 => 
                           n1159, A => n1704, ZN => n1699);
   U1694 : AOI22_X1 port map( A1 => n1161, A2 => REGISTERS_27_29_port, B1 => 
                           n1162, B2 => REGISTERS_26_29_port, ZN => n1704);
   U1695 : INV_X1 port map( A => REGISTERS_24_29_port, ZN => n1033);
   U1696 : INV_X1 port map( A => REGISTERS_25_29_port, ZN => n1032);
   U1697 : OAI221_X1 port map( B1 => n1035, B2 => n1163, C1 => n1036, C2 => 
                           n1164, A => n1705, ZN => n1698);
   U1698 : AOI22_X1 port map( A1 => n1166, A2 => REGISTERS_29_29_port, B1 => 
                           n1167, B2 => REGISTERS_28_29_port, ZN => n1705);
   U1699 : INV_X1 port map( A => REGISTERS_30_29_port, ZN => n1036);
   U1700 : INV_X1 port map( A => REGISTERS_31_29_port, ZN => n1035);
   U1701 : NOR4_X1 port map( A1 => n1706, A2 => n1707, A3 => n1708, A4 => n1709
                           , ZN => n1696);
   U1703 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_3_29_port, B1 => 
                           n1176, B2 => REGISTERS_2_29_port, ZN => n1710);
   U1704 : INV_X1 port map( A => REGISTERS_1_29_port, ZN => n1042);
   U1705 : OAI221_X1 port map( B1 => n1045, B2 => n1177, C1 => n1046, C2 => 
                           n1178, A => n1711, ZN => n1708);
   U1706 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_7_29_port, B1 => 
                           n1181, B2 => REGISTERS_6_29_port, ZN => n1711);
   U1707 : INV_X1 port map( A => REGISTERS_4_29_port, ZN => n1046);
   U1708 : INV_X1 port map( A => REGISTERS_5_29_port, ZN => n1045);
   U1709 : OAI221_X1 port map( B1 => n1048, B2 => n1182, C1 => n1049, C2 => 
                           n1183, A => n1712, ZN => n1707);
   U1710 : AOI22_X1 port map( A1 => n1185, A2 => REGISTERS_11_29_port, B1 => 
                           n1186, B2 => REGISTERS_10_29_port, ZN => n1712);
   U1711 : INV_X1 port map( A => REGISTERS_8_29_port, ZN => n1049);
   U1712 : INV_X1 port map( A => REGISTERS_9_29_port, ZN => n1048);
   U1713 : OAI221_X1 port map( B1 => n1051, B2 => n1187, C1 => n1052, C2 => 
                           n1188, A => n1713, ZN => n1706);
   U1714 : AOI22_X1 port map( A1 => n1190, A2 => REGISTERS_15_29_port, B1 => 
                           n1191, B2 => REGISTERS_14_29_port, ZN => n1713);
   U1715 : INV_X1 port map( A => REGISTERS_12_29_port, ZN => n1052);
   U1716 : INV_X1 port map( A => REGISTERS_13_29_port, ZN => n1051);
   U1717 : NAND2_X1 port map( A1 => n1714, A2 => n1715, ZN => N4216);
   U1718 : NOR4_X1 port map( A1 => n1716, A2 => n1717, A3 => n1718, A4 => n1719
                           , ZN => n1715);
   U1719 : OAI221_X1 port map( B1 => n1060, B2 => n1148, C1 => n1061, C2 => 
                           n1149, A => n1720, ZN => n1719);
   U1720 : AOI22_X1 port map( A1 => n1151, A2 => REGISTERS_19_30_port, B1 => 
                           n1152, B2 => REGISTERS_18_30_port, ZN => n1720);
   U1721 : INV_X1 port map( A => REGISTERS_16_30_port, ZN => n1061);
   U1722 : INV_X1 port map( A => REGISTERS_17_30_port, ZN => n1060);
   U1723 : OAI221_X1 port map( B1 => n1063, B2 => n1153, C1 => n1064, C2 => 
                           n1154, A => n1721, ZN => n1718);
   U1724 : AOI22_X1 port map( A1 => n1156, A2 => REGISTERS_23_30_port, B1 => 
                           n1157, B2 => REGISTERS_22_30_port, ZN => n1721);
   U1725 : INV_X1 port map( A => REGISTERS_20_30_port, ZN => n1064);
   U1726 : INV_X1 port map( A => REGISTERS_21_30_port, ZN => n1063);
   U1727 : OAI221_X1 port map( B1 => n1066, B2 => n1158, C1 => n1067, C2 => 
                           n1159, A => n1722, ZN => n1717);
   U1728 : AOI22_X1 port map( A1 => n1161, A2 => REGISTERS_27_30_port, B1 => 
                           n1162, B2 => REGISTERS_26_30_port, ZN => n1722);
   U1729 : INV_X1 port map( A => REGISTERS_24_30_port, ZN => n1067);
   U1730 : INV_X1 port map( A => REGISTERS_25_30_port, ZN => n1066);
   U1731 : OAI221_X1 port map( B1 => n1069, B2 => n1163, C1 => n1070, C2 => 
                           n1164, A => n1723, ZN => n1716);
   U1732 : AOI22_X1 port map( A1 => n1166, A2 => REGISTERS_29_30_port, B1 => 
                           n1167, B2 => REGISTERS_28_30_port, ZN => n1723);
   U1733 : INV_X1 port map( A => REGISTERS_30_30_port, ZN => n1070);
   U1734 : INV_X1 port map( A => REGISTERS_31_30_port, ZN => n1069);
   U1735 : NOR4_X1 port map( A1 => n1724, A2 => n1725, A3 => n1726, A4 => n1727
                           , ZN => n1714);
   U1737 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_3_30_port, B1 => 
                           n1176, B2 => REGISTERS_2_30_port, ZN => n1728);
   U1738 : INV_X1 port map( A => REGISTERS_1_30_port, ZN => n1076);
   U1739 : OAI221_X1 port map( B1 => n1079, B2 => n1177, C1 => n1080, C2 => 
                           n1178, A => n1729, ZN => n1726);
   U1740 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_7_30_port, B1 => 
                           n1181, B2 => REGISTERS_6_30_port, ZN => n1729);
   U1741 : INV_X1 port map( A => REGISTERS_4_30_port, ZN => n1080);
   U1742 : INV_X1 port map( A => REGISTERS_5_30_port, ZN => n1079);
   U1743 : OAI221_X1 port map( B1 => n1082, B2 => n1182, C1 => n1083, C2 => 
                           n1183, A => n1730, ZN => n1725);
   U1744 : AOI22_X1 port map( A1 => n1185, A2 => REGISTERS_11_30_port, B1 => 
                           n1186, B2 => REGISTERS_10_30_port, ZN => n1730);
   U1745 : INV_X1 port map( A => REGISTERS_8_30_port, ZN => n1083);
   U1746 : INV_X1 port map( A => REGISTERS_9_30_port, ZN => n1082);
   U1747 : OAI221_X1 port map( B1 => n1085, B2 => n1187, C1 => n1086, C2 => 
                           n1188, A => n1731, ZN => n1724);
   U1748 : AOI22_X1 port map( A1 => n1190, A2 => REGISTERS_15_30_port, B1 => 
                           n1191, B2 => REGISTERS_14_30_port, ZN => n1731);
   U1749 : INV_X1 port map( A => REGISTERS_12_30_port, ZN => n1086);
   U1750 : INV_X1 port map( A => REGISTERS_13_30_port, ZN => n1085);
   U1751 : NAND2_X1 port map( A1 => n1732, A2 => n1733, ZN => N4215);
   U1752 : NOR4_X1 port map( A1 => n1734, A2 => n1735, A3 => n1736, A4 => n1737
                           , ZN => n1733);
   U1753 : OAI221_X1 port map( B1 => n1094, B2 => n1148, C1 => n1095, C2 => 
                           n1149, A => n1738, ZN => n1737);
   U1754 : AOI22_X1 port map( A1 => n1151, A2 => REGISTERS_19_31_port, B1 => 
                           n1152, B2 => REGISTERS_18_31_port, ZN => n1738);
   U1758 : INV_X1 port map( A => REGISTERS_16_31_port, ZN => n1095);
   U1760 : INV_X1 port map( A => REGISTERS_17_31_port, ZN => n1094);
   U1761 : OAI221_X1 port map( B1 => n1101, B2 => n1153, C1 => n1102, C2 => 
                           n1154, A => n1743, ZN => n1736);
   U1762 : AOI22_X1 port map( A1 => n1156, A2 => REGISTERS_23_31_port, B1 => 
                           n1157, B2 => REGISTERS_22_31_port, ZN => n1743);
   U1766 : AND2_X1 port map( A1 => n1746, A2 => n1747, ZN => n1739);
   U1767 : INV_X1 port map( A => REGISTERS_20_31_port, ZN => n1102);
   U1769 : AND2_X1 port map( A1 => n1746, A2 => ADD_RD1(0), ZN => n1741);
   U1770 : AND2_X1 port map( A1 => ADD_RD1(4), A2 => n1748, ZN => n1746);
   U1771 : INV_X1 port map( A => REGISTERS_21_31_port, ZN => n1101);
   U1772 : OAI221_X1 port map( B1 => n1109, B2 => n1158, C1 => n1110, C2 => 
                           n1159, A => n1749, ZN => n1735);
   U1773 : AOI22_X1 port map( A1 => n1161, A2 => REGISTERS_27_31_port, B1 => 
                           n1162, B2 => REGISTERS_26_31_port, ZN => n1749);
   U1777 : INV_X1 port map( A => REGISTERS_24_31_port, ZN => n1110);
   U1779 : INV_X1 port map( A => REGISTERS_25_31_port, ZN => n1109);
   U1780 : OAI221_X1 port map( B1 => n1114, B2 => n1163, C1 => n1115, C2 => 
                           n1164, A => n1752, ZN => n1734);
   U1781 : AOI22_X1 port map( A1 => n1166, A2 => REGISTERS_29_31_port, B1 => 
                           n1167, B2 => REGISTERS_28_31_port, ZN => n1752);
   U1785 : AND2_X1 port map( A1 => n1753, A2 => n1747, ZN => n1750);
   U1786 : INV_X1 port map( A => REGISTERS_30_31_port, ZN => n1115);
   U1788 : AND2_X1 port map( A1 => ADD_RD1(0), A2 => n1753, ZN => n1751);
   U1789 : AND2_X1 port map( A1 => ADD_RD1(4), A2 => ADD_RD1(3), ZN => n1753);
   U1790 : INV_X1 port map( A => REGISTERS_31_31_port, ZN => n1114);
   U1791 : NOR4_X1 port map( A1 => n1754, A2 => n1755, A3 => n1756, A4 => n1757
                           , ZN => n1732);
   U1793 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_3_31_port, B1 => 
                           n1176, B2 => REGISTERS_2_31_port, ZN => n1758);
   U1798 : INV_X1 port map( A => REGISTERS_1_31_port, ZN => n1122);
   U1799 : OAI221_X1 port map( B1 => n1127, B2 => n1177, C1 => n1128, C2 => 
                           n1178, A => n1761, ZN => n1756);
   U1800 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_7_31_port, B1 => 
                           n1181, B2 => REGISTERS_6_31_port, ZN => n1761);
   U1804 : AND2_X1 port map( A1 => n1762, A2 => n1747, ZN => n1759);
   U1805 : INV_X1 port map( A => REGISTERS_4_31_port, ZN => n1128);
   U1807 : AND2_X1 port map( A1 => n1762, A2 => ADD_RD1(0), ZN => n1760);
   U1808 : NOR2_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), ZN => n1762);
   U1809 : INV_X1 port map( A => REGISTERS_5_31_port, ZN => n1127);
   U1810 : OAI221_X1 port map( B1 => n1131, B2 => n1182, C1 => n1132, C2 => 
                           n1183, A => n1763, ZN => n1755);
   U1811 : AOI22_X1 port map( A1 => n1185, A2 => REGISTERS_11_31_port, B1 => 
                           n1186, B2 => REGISTERS_10_31_port, ZN => n1763);
   U1814 : NOR2_X1 port map( A1 => n1766, A2 => ADD_RD1(2), ZN => n1740);
   U1816 : INV_X1 port map( A => REGISTERS_8_31_port, ZN => n1132);
   U1818 : NOR2_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), ZN => n1742);
   U1819 : INV_X1 port map( A => REGISTERS_9_31_port, ZN => n1131);
   U1820 : OAI221_X1 port map( B1 => n1137, B2 => n1187, C1 => n1138, C2 => 
                           n1188, A => n1767, ZN => n1754);
   U1821 : AOI22_X1 port map( A1 => n1190, A2 => REGISTERS_15_31_port, B1 => 
                           n1191, B2 => REGISTERS_14_31_port, ZN => n1767);
   U1824 : NOR2_X1 port map( A1 => n1768, A2 => n1766, ZN => n1744);
   U1825 : INV_X1 port map( A => ADD_RD1(1), ZN => n1766);
   U1827 : AND2_X1 port map( A1 => n1769, A2 => n1747, ZN => n1764);
   U1828 : INV_X1 port map( A => ADD_RD1(0), ZN => n1747);
   U1829 : INV_X1 port map( A => REGISTERS_12_31_port, ZN => n1138);
   U1832 : INV_X1 port map( A => ADD_RD1(2), ZN => n1768);
   U1833 : AND2_X1 port map( A1 => n1769, A2 => ADD_RD1(0), ZN => n1765);
   U1834 : NOR2_X1 port map( A1 => n1748, A2 => ADD_RD1(4), ZN => n1769);
   U1835 : INV_X1 port map( A => ADD_RD1(3), ZN => n1748);
   U1836 : INV_X1 port map( A => REGISTERS_13_31_port, ZN => n1137);
   U1837 : NAND2_X1 port map( A1 => n1770, A2 => n193, ZN => N4083);
   U1838 : NAND3_X1 port map( A1 => n1771, A2 => n1, A3 => n1773, ZN => n1770);
   U1839 : NAND2_X1 port map( A1 => n1774, A2 => n193, ZN => N4019);
   U1840 : NAND3_X1 port map( A1 => n1773, A2 => n1772, A3 => n1775, ZN => 
                           n1774);
   U1841 : NAND2_X1 port map( A1 => n1776, A2 => n193, ZN => N3955);
   U1842 : NAND3_X1 port map( A1 => n1773, A2 => n1772, A3 => n1777, ZN => 
                           n1776);
   U1843 : NAND2_X1 port map( A1 => n1778, A2 => n193, ZN => N3891);
   U1844 : NAND3_X1 port map( A1 => n1773, A2 => n1772, A3 => n1779, ZN => 
                           n1778);
   U1845 : NAND2_X1 port map( A1 => n1780, A2 => n193, ZN => N3827);
   U1846 : NAND3_X1 port map( A1 => n1773, A2 => n1772, A3 => n1781, ZN => 
                           n1780);
   U1847 : NAND2_X1 port map( A1 => n1782, A2 => n193, ZN => N3763);
   U1848 : NAND3_X1 port map( A1 => n1773, A2 => n1772, A3 => n1783, ZN => 
                           n1782);
   U1849 : NAND2_X1 port map( A1 => n1784, A2 => n193, ZN => N3699);
   U1850 : NAND3_X1 port map( A1 => n1773, A2 => n1772, A3 => n1785, ZN => 
                           n1784);
   U1851 : NOR2_X1 port map( A1 => ADD_WR(3), A2 => ADD_WR(4), ZN => n1773);
   U1852 : NAND2_X1 port map( A1 => n1786, A2 => n193, ZN => N3635);
   U1853 : NAND3_X1 port map( A1 => n1787, A2 => n1772, A3 => n1788, ZN => 
                           n1786);
   U1854 : NAND2_X1 port map( A1 => n1789, A2 => n193, ZN => N3571);
   U1855 : NAND3_X1 port map( A1 => n1771, A2 => n1772, A3 => n1787, ZN => 
                           n1789);
   U1856 : NAND2_X1 port map( A1 => n1790, A2 => n193, ZN => N3507);
   U1857 : NAND3_X1 port map( A1 => n1775, A2 => n1772, A3 => n1787, ZN => 
                           n1790);
   U1858 : NAND2_X1 port map( A1 => n1791, A2 => n193, ZN => N3443);
   U1859 : NAND3_X1 port map( A1 => n1777, A2 => n1772, A3 => n1787, ZN => 
                           n1791);
   U1860 : NAND2_X1 port map( A1 => n1792, A2 => n193, ZN => N3379);
   U1861 : NAND3_X1 port map( A1 => n1779, A2 => n1772, A3 => n1787, ZN => 
                           n1792);
   U1862 : NAND2_X1 port map( A1 => n1793, A2 => n227, ZN => N3315);
   U1863 : NAND3_X1 port map( A1 => n1781, A2 => n1772, A3 => n1787, ZN => 
                           n1793);
   U1864 : NAND2_X1 port map( A1 => n1794, A2 => n227, ZN => N3251);
   U1865 : NAND3_X1 port map( A1 => n1783, A2 => n1772, A3 => n1787, ZN => 
                           n1794);
   U1866 : NAND2_X1 port map( A1 => n1795, A2 => n227, ZN => N3187);
   U1867 : NAND3_X1 port map( A1 => n1785, A2 => n1772, A3 => n1787, ZN => 
                           n1795);
   U1868 : NOR2_X1 port map( A1 => n1796, A2 => ADD_WR(4), ZN => n1787);
   U1869 : NAND2_X1 port map( A1 => n1797, A2 => n227, ZN => N3123);
   U1870 : NAND3_X1 port map( A1 => n1788, A2 => n1772, A3 => n1798, ZN => 
                           n1797);
   U1871 : NAND2_X1 port map( A1 => n1799, A2 => n227, ZN => N3059);
   U1872 : NAND3_X1 port map( A1 => n1771, A2 => n1772, A3 => n1798, ZN => 
                           n1799);
   U1873 : NAND2_X1 port map( A1 => n1800, A2 => n227, ZN => N2995);
   U1874 : NAND3_X1 port map( A1 => n1775, A2 => n1772, A3 => n1798, ZN => 
                           n1800);
   U1875 : NAND2_X1 port map( A1 => n1801, A2 => n227, ZN => N2931);
   U1876 : NAND3_X1 port map( A1 => n1777, A2 => n1772, A3 => n1798, ZN => 
                           n1801);
   U1877 : NAND2_X1 port map( A1 => n1802, A2 => n227, ZN => N2867);
   U1878 : NAND3_X1 port map( A1 => n1779, A2 => n1772, A3 => n1798, ZN => 
                           n1802);
   U1879 : NAND2_X1 port map( A1 => n1803, A2 => n227, ZN => N2803);
   U1880 : NAND3_X1 port map( A1 => n1781, A2 => n1772, A3 => n1798, ZN => 
                           n1803);
   U1881 : NAND2_X1 port map( A1 => n1804, A2 => n227, ZN => N2739);
   U1882 : NAND3_X1 port map( A1 => n1783, A2 => n1772, A3 => n1798, ZN => 
                           n1804);
   U1883 : NAND2_X1 port map( A1 => n1805, A2 => n227, ZN => N2675);
   U1884 : NAND3_X1 port map( A1 => n1785, A2 => n1772, A3 => n1798, ZN => 
                           n1805);
   U1885 : AND2_X1 port map( A1 => ADD_WR(4), A2 => n1796, ZN => n1798);
   U1886 : INV_X1 port map( A => ADD_WR(3), ZN => n1796);
   U1887 : NAND2_X1 port map( A1 => n1806, A2 => n227, ZN => N2611);
   U1888 : NAND3_X1 port map( A1 => n1788, A2 => n1772, A3 => n1807, ZN => 
                           n1806);
   U1889 : NOR3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(2), A3 => ADD_WR(0),
                           ZN => n1788);
   U1890 : NAND2_X1 port map( A1 => n1808, A2 => n261, ZN => N2547);
   U1891 : NAND3_X1 port map( A1 => n1771, A2 => n1772, A3 => n1807, ZN => 
                           n1808);
   U1892 : NOR3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(2), A3 => n1809, ZN 
                           => n1771);
   U1893 : NAND2_X1 port map( A1 => n1810, A2 => n261, ZN => N2483);
   U1894 : NAND3_X1 port map( A1 => n1775, A2 => n1772, A3 => n1807, ZN => 
                           n1810);
   U1895 : NOR3_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(2), A3 => n1811, ZN 
                           => n1775);
   U1896 : NAND2_X1 port map( A1 => n1812, A2 => n261, ZN => N2419);
   U1897 : NAND3_X1 port map( A1 => n1777, A2 => n1, A3 => n1807, ZN => n1812);
   U1898 : NOR3_X1 port map( A1 => n1809, A2 => ADD_WR(2), A3 => n1811, ZN => 
                           n1777);
   U1899 : NAND2_X1 port map( A1 => n1813, A2 => n261, ZN => N2355);
   U1900 : NAND3_X1 port map( A1 => n1779, A2 => n1, A3 => n1807, ZN => n1813);
   U1901 : NOR3_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(1), A3 => n1814, ZN 
                           => n1779);
   U1902 : NAND2_X1 port map( A1 => n1815, A2 => n261, ZN => N2291);
   U1903 : NAND3_X1 port map( A1 => n1781, A2 => n1, A3 => n1807, ZN => n1815);
   U1904 : NOR3_X1 port map( A1 => n1809, A2 => ADD_WR(1), A3 => n1814, ZN => 
                           n1781);
   U1905 : NAND2_X1 port map( A1 => n1816, A2 => n261, ZN => N2227);
   U1906 : NAND3_X1 port map( A1 => n1783, A2 => n1, A3 => n1807, ZN => n1816);
   U1907 : NOR3_X1 port map( A1 => n1811, A2 => ADD_WR(0), A3 => n1814, ZN => 
                           n1783);
   U1908 : AND2_X1 port map( A1 => DATAIN(31), A2 => n261, ZN => N4148);
   U1909 : AND2_X1 port map( A1 => DATAIN(30), A2 => n329, ZN => N4146);
   U1910 : AND2_X1 port map( A1 => DATAIN(29), A2 => n329, ZN => N4144);
   U1911 : AND2_X1 port map( A1 => DATAIN(28), A2 => n329, ZN => N4142);
   U1912 : AND2_X1 port map( A1 => DATAIN(27), A2 => n329, ZN => N4140);
   U1913 : AND2_X1 port map( A1 => DATAIN(26), A2 => n329, ZN => N4138);
   U1914 : AND2_X1 port map( A1 => DATAIN(25), A2 => n329, ZN => N4136);
   U1915 : AND2_X1 port map( A1 => DATAIN(24), A2 => n329, ZN => N4134);
   U1916 : AND2_X1 port map( A1 => DATAIN(23), A2 => n329, ZN => N4132);
   U1917 : AND2_X1 port map( A1 => DATAIN(22), A2 => n329, ZN => N4130);
   U1918 : AND2_X1 port map( A1 => DATAIN(21), A2 => n329, ZN => N4128);
   U1919 : AND2_X1 port map( A1 => DATAIN(20), A2 => n295, ZN => N4126);
   U1920 : AND2_X1 port map( A1 => DATAIN(19), A2 => n295, ZN => N4124);
   U1921 : AND2_X1 port map( A1 => DATAIN(18), A2 => n295, ZN => N4122);
   U1922 : AND2_X1 port map( A1 => DATAIN(17), A2 => n295, ZN => N4120);
   U1923 : AND2_X1 port map( A1 => DATAIN(16), A2 => n295, ZN => N4118);
   U1924 : AND2_X1 port map( A1 => DATAIN(15), A2 => n295, ZN => N4116);
   U1925 : AND2_X1 port map( A1 => DATAIN(14), A2 => n295, ZN => N4114);
   U1926 : AND2_X1 port map( A1 => DATAIN(13), A2 => n295, ZN => N4112);
   U1927 : AND2_X1 port map( A1 => DATAIN(12), A2 => n295, ZN => N4110);
   U1928 : AND2_X1 port map( A1 => DATAIN(11), A2 => n295, ZN => N4108);
   U1929 : AND2_X1 port map( A1 => DATAIN(10), A2 => n295, ZN => N4106);
   U1930 : AND2_X1 port map( A1 => DATAIN(9), A2 => n295, ZN => N4104);
   U1931 : AND2_X1 port map( A1 => DATAIN(8), A2 => n295, ZN => N4102);
   U1932 : AND2_X1 port map( A1 => DATAIN(7), A2 => n295, ZN => N4100);
   U1933 : AND2_X1 port map( A1 => DATAIN(6), A2 => n295, ZN => N4098);
   U1934 : AND2_X1 port map( A1 => DATAIN(5), A2 => n295, ZN => N4096);
   U1935 : AND2_X1 port map( A1 => DATAIN(4), A2 => n261, ZN => N4094);
   U1936 : AND2_X1 port map( A1 => DATAIN(3), A2 => n261, ZN => N4092);
   U1937 : AND2_X1 port map( A1 => DATAIN(2), A2 => n261, ZN => N4090);
   U1938 : AND2_X1 port map( A1 => DATAIN(1), A2 => n261, ZN => N4088);
   U1939 : AND2_X1 port map( A1 => DATAIN(0), A2 => n261, ZN => N4086);
   U1940 : NAND2_X1 port map( A1 => n1817, A2 => n261, ZN => N2163);
   U1941 : NAND3_X1 port map( A1 => n1785, A2 => n1, A3 => n1807, ZN => n1817);
   U1942 : AND2_X1 port map( A1 => ADD_WR(4), A2 => ADD_WR(3), ZN => n1807);
   U1943 : AND2_X1 port map( A1 => WR, A2 => ENABLE, ZN => n1772);
   U1944 : NOR3_X1 port map( A1 => n1811, A2 => n1809, A3 => n1814, ZN => n1785
                           );
   U1945 : INV_X1 port map( A => ADD_WR(2), ZN => n1814);
   U1946 : INV_X1 port map( A => ADD_WR(0), ZN => n1809);
   U1947 : INV_X1 port map( A => ADD_WR(1), ZN => n1811);
   U3 : NOR2_X2 port map( A1 => n1140, A2 => ADD_RD2(1), ZN => n1105);
   U4 : NOR2_X2 port map( A1 => n1768, A2 => ADD_RD1(1), ZN => n1745);
   U5 : CLKBUF_X1 port map( A => n1772, Z => n1);
   U6 : AND2_X2 port map( A1 => n1759, A2 => n1744, ZN => n1181);
   U7 : AND2_X2 port map( A1 => n1764, A2 => n1744, ZN => n1191);
   U8 : AND2_X2 port map( A1 => n1739, A2 => n1740, ZN => n1152);
   U9 : AND2_X2 port map( A1 => n1745, A2 => n1750, ZN => n1167);
   U10 : AND2_X2 port map( A1 => n1740, A2 => n1750, ZN => n1162);
   U11 : AND2_X2 port map( A1 => n1759, A2 => n1740, ZN => n1176);
   U12 : AND2_X2 port map( A1 => n1764, A2 => n1740, ZN => n1186);
   U13 : NAND2_X2 port map( A1 => n1125, A2 => n1105, ZN => n49);
   U14 : AND2_X2 port map( A1 => n1739, A2 => n1744, ZN => n1157);
   U15 : NAND2_X2 port map( A1 => n1097, A2 => n1105, ZN => n17);
   U16 : NAND2_X2 port map( A1 => n1100, A2 => n1112, ZN => n24);
   U17 : NAND2_X2 port map( A1 => n1134, A2 => n1105, ZN => n63);
   U18 : NAND2_X2 port map( A1 => n1112, A2 => n1104, ZN => n31);
   U19 : NAND2_X2 port map( A1 => n1134, A2 => n1100, ZN => n56);
   U20 : NAND2_X2 port map( A1 => n1097, A2 => n1100, ZN => n10);
   U21 : NAND2_X2 port map( A1 => n1760, A2 => n1742, ZN => n1172);
   U22 : NAND2_X2 port map( A1 => n1759, A2 => n1745, ZN => n1178);
   U23 : NAND2_X2 port map( A1 => n1750, A2 => n1744, ZN => n1164);
   U24 : NAND2_X2 port map( A1 => n1742, A2 => n1750, ZN => n1159);
   U25 : NAND2_X2 port map( A1 => n1764, A2 => n1742, ZN => n1183);
   U26 : NAND2_X2 port map( A1 => n1739, A2 => n1742, ZN => n1149);
   U27 : NAND2_X2 port map( A1 => n1764, A2 => n1745, ZN => n1188);
   U28 : NAND2_X2 port map( A1 => n1739, A2 => n1745, ZN => n1154);
   U29 : AND2_X2 port map( A1 => n1097, A2 => n1098, ZN => n14);
   U30 : AND2_X2 port map( A1 => n1125, A2 => n1098, ZN => n46);
   U31 : AND2_X2 port map( A1 => n1097, A2 => n1104, ZN => n21);
   U32 : AND2_X2 port map( A1 => n1134, A2 => n1104, ZN => n67);
   U33 : AND2_X2 port map( A1 => n1105, A2 => n1112, ZN => n35);
   U34 : AND2_X2 port map( A1 => n1134, A2 => n1098, ZN => n60);
   U47 : AND2_X2 port map( A1 => n1098, A2 => n1112, ZN => n28);
   U66 : NAND2_X2 port map( A1 => n1765, A2 => n1745, ZN => n1187);
   U85 : AND2_X2 port map( A1 => n1125, A2 => n1104, ZN => n53);
   U104 : NAND2_X2 port map( A1 => n1741, A2 => n1742, ZN => n1148);
   U123 : NAND2_X2 port map( A1 => n1744, A2 => n1751, ZN => n1163);
   U142 : NAND2_X2 port map( A1 => n1765, A2 => n1742, ZN => n1182);
   U161 : NAND2_X2 port map( A1 => n1760, A2 => n1745, ZN => n1177);
   U180 : NAND2_X2 port map( A1 => n1741, A2 => n1745, ZN => n1153);
   U199 : NAND2_X2 port map( A1 => n1742, A2 => n1751, ZN => n1158);
   U218 : AND2_X2 port map( A1 => n1740, A2 => n1751, ZN => n1161);
   U237 : AND2_X2 port map( A1 => n1745, A2 => n1751, ZN => n1166);
   U256 : AND2_X2 port map( A1 => n1760, A2 => n1740, ZN => n1175);
   U275 : AND2_X2 port map( A1 => n1741, A2 => n1744, ZN => n1156);
   U294 : AND2_X2 port map( A1 => n1741, A2 => n1740, ZN => n1151);
   U313 : AND2_X2 port map( A1 => n1760, A2 => n1744, ZN => n1180);
   U332 : AND2_X2 port map( A1 => n1765, A2 => n1740, ZN => n1185);
   U351 : AND2_X2 port map( A1 => n1765, A2 => n1744, ZN => n1190);
   U370 : AND2_X2 port map( A1 => n1126, A2 => n1104, ZN => n52);
   U389 : AND2_X2 port map( A1 => n1099, A2 => n1098, ZN => n13);
   U408 : AND2_X2 port map( A1 => n1099, A2 => n1104, ZN => n20);
   U427 : AND2_X2 port map( A1 => n1126, A2 => n1098, ZN => n45);
   U446 : AND2_X2 port map( A1 => n1135, A2 => n1098, ZN => n59);
   U465 : AND2_X2 port map( A1 => n1135, A2 => n1104, ZN => n66);
   U484 : AND2_X2 port map( A1 => n1098, A2 => n1113, ZN => n27);
   U503 : AND2_X2 port map( A1 => n1105, A2 => n1113, ZN => n34);
   U522 : NAND2_X2 port map( A1 => n1104, A2 => n1113, ZN => n29);
   U541 : NAND2_X2 port map( A1 => n1126, A2 => n1105, ZN => n47);
   U560 : NAND2_X2 port map( A1 => n1135, A2 => n1100, ZN => n54);
   U579 : NAND2_X2 port map( A1 => n1100, A2 => n1113, ZN => n22);
   U598 : NAND2_X2 port map( A1 => n1099, A2 => n1105, ZN => n15);
   U617 : NAND2_X2 port map( A1 => n1135, A2 => n1105, ZN => n61);
   U629 : NAND2_X2 port map( A1 => n1126, A2 => n1100, ZN => n40);
   U630 : NAND2_X2 port map( A1 => n1099, A2 => n1100, ZN => n8);
   U639 : OAI21_X1 port map( B1 => n40, B2 => n41, A => n44, ZN => n39);
   U644 : OAI21_X1 port map( B1 => n40, B2 => n90, A => n92, ZN => n89);
   U645 : OAI21_X1 port map( B1 => n40, B2 => n124, A => n126, ZN => n123);
   U646 : OAI21_X1 port map( B1 => n40, B2 => n158, A => n160, ZN => n157);
   U647 : OAI21_X1 port map( B1 => n40, B2 => n192, A => n194, ZN => n191);
   U650 : OAI21_X1 port map( B1 => n40, B2 => n226, A => n228, ZN => n225);
   U651 : OAI21_X1 port map( B1 => n40, B2 => n260, A => n262, ZN => n259);
   U652 : OAI21_X1 port map( B1 => n40, B2 => n294, A => n296, ZN => n293);
   U654 : OAI21_X1 port map( B1 => n40, B2 => n328, A => n330, ZN => n327);
   U658 : OAI21_X1 port map( B1 => n40, B2 => n362, A => n364, ZN => n361);
   U660 : OAI21_X1 port map( B1 => n40, B2 => n396, A => n398, ZN => n395);
   U661 : OAI21_X1 port map( B1 => n40, B2 => n430, A => n432, ZN => n429);
   U662 : OAI21_X1 port map( B1 => n40, B2 => n464, A => n466, ZN => n463);
   U663 : OAI21_X1 port map( B1 => n40, B2 => n498, A => n500, ZN => n497);
   U666 : OAI21_X1 port map( B1 => n40, B2 => n532, A => n534, ZN => n531);
   U667 : OAI21_X1 port map( B1 => n40, B2 => n566, A => n568, ZN => n565);
   U668 : OAI21_X1 port map( B1 => n40, B2 => n600, A => n602, ZN => n599);
   U670 : OAI21_X1 port map( B1 => n40, B2 => n634, A => n636, ZN => n633);
   U675 : OAI21_X1 port map( B1 => n40, B2 => n668, A => n670, ZN => n667);
   U676 : OAI21_X1 port map( B1 => n40, B2 => n702, A => n704, ZN => n701);
   U678 : OAI21_X1 port map( B1 => n40, B2 => n736, A => n738, ZN => n735);
   U679 : OAI21_X1 port map( B1 => n40, B2 => n770, A => n772, ZN => n769);
   U683 : OAI21_X1 port map( B1 => n40, B2 => n804, A => n806, ZN => n803);
   U684 : OAI21_X1 port map( B1 => n40, B2 => n838, A => n840, ZN => n837);
   U687 : OAI21_X1 port map( B1 => n40, B2 => n872, A => n874, ZN => n871);
   U690 : OAI21_X1 port map( B1 => n40, B2 => n906, A => n908, ZN => n905);
   U691 : OAI21_X1 port map( B1 => n40, B2 => n940, A => n942, ZN => n939);
   U716 : OAI21_X1 port map( B1 => n40, B2 => n974, A => n976, ZN => n973);
   U750 : OAI21_X1 port map( B1 => n40, B2 => n1008, A => n1010, ZN => n1007);
   U784 : OAI21_X1 port map( B1 => n40, B2 => n1042, A => n1044, ZN => n1041);
   U818 : OAI21_X1 port map( B1 => n40, B2 => n1076, A => n1078, ZN => n1075);
   U852 : OAI21_X1 port map( B1 => n40, B2 => n1122, A => n1124, ZN => n1121);
   U886 : OAI21_X1 port map( B1 => n41, B2 => n1172, A => n1174, ZN => n1171);
   U920 : OAI21_X1 port map( B1 => n90, B2 => n1172, A => n1206, ZN => n1205);
   U954 : OAI21_X1 port map( B1 => n124, B2 => n1172, A => n1224, ZN => n1223);
   U988 : OAI21_X1 port map( B1 => n158, B2 => n1172, A => n1242, ZN => n1241);
   U1022 : OAI21_X1 port map( B1 => n192, B2 => n1172, A => n1260, ZN => n1259)
                           ;
   U1056 : OAI21_X1 port map( B1 => n226, B2 => n1172, A => n1278, ZN => n1277)
                           ;
   U1090 : OAI21_X1 port map( B1 => n260, B2 => n1172, A => n1296, ZN => n1295)
                           ;
   U1124 : OAI21_X1 port map( B1 => n294, B2 => n1172, A => n1314, ZN => n1313)
                           ;
   U1158 : OAI21_X1 port map( B1 => n328, B2 => n1172, A => n1332, ZN => n1331)
                           ;
   U1192 : OAI21_X1 port map( B1 => n362, B2 => n1172, A => n1350, ZN => n1349)
                           ;
   U1226 : OAI21_X1 port map( B1 => n396, B2 => n1172, A => n1368, ZN => n1367)
                           ;
   U1260 : OAI21_X1 port map( B1 => n430, B2 => n1172, A => n1386, ZN => n1385)
                           ;
   U1294 : OAI21_X1 port map( B1 => n464, B2 => n1172, A => n1404, ZN => n1403)
                           ;
   U1328 : OAI21_X1 port map( B1 => n498, B2 => n1172, A => n1422, ZN => n1421)
                           ;
   U1362 : OAI21_X1 port map( B1 => n532, B2 => n1172, A => n1440, ZN => n1439)
                           ;
   U1396 : OAI21_X1 port map( B1 => n566, B2 => n1172, A => n1458, ZN => n1457)
                           ;
   U1430 : OAI21_X1 port map( B1 => n600, B2 => n1172, A => n1476, ZN => n1475)
                           ;
   U1464 : OAI21_X1 port map( B1 => n634, B2 => n1172, A => n1494, ZN => n1493)
                           ;
   U1498 : OAI21_X1 port map( B1 => n668, B2 => n1172, A => n1512, ZN => n1511)
                           ;
   U1532 : OAI21_X1 port map( B1 => n702, B2 => n1172, A => n1530, ZN => n1529)
                           ;
   U1566 : OAI21_X1 port map( B1 => n736, B2 => n1172, A => n1548, ZN => n1547)
                           ;
   U1600 : OAI21_X1 port map( B1 => n770, B2 => n1172, A => n1566, ZN => n1565)
                           ;
   U1634 : OAI21_X1 port map( B1 => n804, B2 => n1172, A => n1584, ZN => n1583)
                           ;
   U1668 : OAI21_X1 port map( B1 => n838, B2 => n1172, A => n1602, ZN => n1601)
                           ;
   U1702 : OAI21_X1 port map( B1 => n872, B2 => n1172, A => n1620, ZN => n1619)
                           ;
   U1736 : OAI21_X1 port map( B1 => n906, B2 => n1172, A => n1638, ZN => n1637)
                           ;
   U1755 : OAI21_X1 port map( B1 => n940, B2 => n1172, A => n1656, ZN => n1655)
                           ;
   U1756 : OAI21_X1 port map( B1 => n974, B2 => n1172, A => n1674, ZN => n1673)
                           ;
   U1757 : OAI21_X1 port map( B1 => n1008, B2 => n1172, A => n1692, ZN => n1691
                           );
   U1759 : OAI21_X1 port map( B1 => n1042, B2 => n1172, A => n1710, ZN => n1709
                           );
   U1763 : OAI21_X1 port map( B1 => n1076, B2 => n1172, A => n1728, ZN => n1727
                           );
   U1764 : OAI21_X1 port map( B1 => n1122, B2 => n1172, A => n1758, ZN => n1757
                           );
   U631 : CLKBUF_X1 port map( A => RESET, Z => n193);
   U632 : CLKBUF_X1 port map( A => RESET, Z => n227);
   U635 : CLKBUF_X1 port map( A => RESET, Z => n261);
   U636 : CLKBUF_X1 port map( A => RESET, Z => n295);
   U637 : CLKBUF_X1 port map( A => RESET, Z => n329);

end SYN_A;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity alu_NUMBIT32 is

   port( DATA1, DATA2 : in std_logic_vector (31 downto 0);  FUNC : in 
         std_logic_vector (0 to 4);  OUTALU : out std_logic_vector (31 downto 
         0));

end alu_NUMBIT32;

architecture SYN_STRUCT of alu_NUMBIT32 is

   component BUF_X8
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI222_X4
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component shifter
      port( R : in std_logic_vector (31 downto 0);  Offset : in 
            std_logic_vector (4 downto 0);  Conf : in std_logic_vector (0 to 1)
            ;  Shift_OUT : out std_logic_vector (31 downto 0));
   end component;
   
   component ComparatorUnit
      port( A_MSB, B_MSB : in std_logic;  SUBIN : in std_logic_vector (31 
            downto 0);  COUT, SIGN_UNSIGN : in std_logic;  OP : in 
            std_logic_vector (0 to 2);  CU_OUT : out std_logic_vector (31 
            downto 0));
   end component;
   
   component logicunit
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  LU_OUT : out std_logic_vector (31 
            downto 0));
   end component;
   
   component P4addersub_N32
      port( A, B : in std_logic_vector (31 downto 0);  sub_add : in std_logic; 
            Y : out std_logic_vector (31 downto 0);  Cout : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal sub_add, Sel_2_port, Conf_1_port, Conf_0_port, Comp_OP_1_port, 
      Comp_OP_0_port, sign_unsign, OUT_adder_31_port, OUT_adder_30_port, 
      OUT_adder_29_port, OUT_adder_28_port, OUT_adder_27_port, 
      OUT_adder_26_port, OUT_adder_25_port, OUT_adder_24_port, 
      OUT_adder_23_port, OUT_adder_22_port, OUT_adder_21_port, 
      OUT_adder_20_port, OUT_adder_19_port, OUT_adder_18_port, 
      OUT_adder_17_port, OUT_adder_16_port, OUT_adder_15_port, 
      OUT_adder_14_port, OUT_adder_13_port, OUT_adder_12_port, 
      OUT_adder_11_port, OUT_adder_10_port, OUT_adder_9_port, OUT_adder_8_port,
      OUT_adder_7_port, OUT_adder_6_port, OUT_adder_5_port, OUT_adder_4_port, 
      OUT_adder_3_port, OUT_adder_2_port, OUT_adder_1_port, OUT_adder_0_port, 
      LU_out_31_port, LU_out_30_port, LU_out_29_port, LU_out_28_port, 
      LU_out_27_port, LU_out_26_port, LU_out_25_port, LU_out_24_port, 
      LU_out_23_port, LU_out_22_port, LU_out_21_port, LU_out_20_port, 
      LU_out_19_port, LU_out_18_port, LU_out_17_port, LU_out_16_port, 
      LU_out_15_port, LU_out_14_port, LU_out_13_port, LU_out_12_port, 
      LU_out_11_port, LU_out_10_port, LU_out_9_port, LU_out_8_port, 
      LU_out_7_port, LU_out_6_port, LU_out_5_port, LU_out_4_port, LU_out_3_port
      , LU_out_2_port, LU_out_1_port, LU_out_0_port, SHIFT_OUT_31_port, 
      SHIFT_OUT_30_port, SHIFT_OUT_29_port, SHIFT_OUT_28_port, 
      SHIFT_OUT_27_port, SHIFT_OUT_26_port, SHIFT_OUT_25_port, 
      SHIFT_OUT_24_port, SHIFT_OUT_23_port, SHIFT_OUT_22_port, 
      SHIFT_OUT_21_port, SHIFT_OUT_20_port, SHIFT_OUT_19_port, 
      SHIFT_OUT_18_port, SHIFT_OUT_17_port, SHIFT_OUT_16_port, 
      SHIFT_OUT_15_port, SHIFT_OUT_14_port, SHIFT_OUT_13_port, 
      SHIFT_OUT_12_port, SHIFT_OUT_11_port, SHIFT_OUT_10_port, SHIFT_OUT_9_port
      , SHIFT_OUT_8_port, SHIFT_OUT_7_port, SHIFT_OUT_6_port, SHIFT_OUT_5_port,
      SHIFT_OUT_4_port, SHIFT_OUT_3_port, SHIFT_OUT_2_port, SHIFT_OUT_1_port, 
      SHIFT_OUT_0_port, CU_OUT_0_port, Adder_Cout, n104, n205, n305, n306, n308
      , n310, n311, n312, n314, n315, n316, n317, n318, n319, n320, n321, n322,
      n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, 
      n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, 
      n347, n348, n352, n353, n355, n356, n360, n359, n358, n357, n354, n349, 
      n313, n309, n307, n361, n362, n363, n364, n365, n366, n367, n368, n369, 
      n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, net126648, 
      net126649, net126650, net126651, net126652, net126653, net126654, 
      net126655, net126656, net126657, net126658, net126659, net126660, 
      net126661, net126662, net126663, net126664, net126665, net126666, 
      net126667, net126668, net126669, net126670, net126671, net126672, 
      net126673, net126674, net126675, net126676, net126677, net126678 : 
      std_logic;

begin
   
   U233 : CLKBUF_X2 port map( A => n104, Z => n306);
   U241 : INV_X1 port map( A => n315, ZN => OUTALU(9));
   U242 : AOI222_X1 port map( A1 => OUT_adder_9_port, A2 => n316, B1 => 
                           LU_out_9_port, B2 => n317, C1 => SHIFT_OUT_9_port, 
                           C2 => n318, ZN => n315);
   U243 : INV_X1 port map( A => n319, ZN => OUTALU(8));
   U244 : AOI222_X1 port map( A1 => OUT_adder_8_port, A2 => n316, B1 => 
                           LU_out_8_port, B2 => n317, C1 => SHIFT_OUT_8_port, 
                           C2 => n318, ZN => n319);
   U245 : INV_X1 port map( A => n320, ZN => OUTALU(7));
   U246 : AOI222_X1 port map( A1 => OUT_adder_7_port, A2 => n316, B1 => 
                           LU_out_7_port, B2 => n317, C1 => SHIFT_OUT_7_port, 
                           C2 => n318, ZN => n320);
   U247 : INV_X1 port map( A => n321, ZN => OUTALU(6));
   U248 : AOI222_X1 port map( A1 => OUT_adder_6_port, A2 => n316, B1 => 
                           LU_out_6_port, B2 => n317, C1 => SHIFT_OUT_6_port, 
                           C2 => n318, ZN => n321);
   U249 : INV_X1 port map( A => n322, ZN => OUTALU(5));
   U250 : AOI222_X1 port map( A1 => OUT_adder_5_port, A2 => n316, B1 => 
                           LU_out_5_port, B2 => n317, C1 => SHIFT_OUT_5_port, 
                           C2 => n318, ZN => n322);
   U251 : INV_X1 port map( A => n323, ZN => OUTALU(4));
   U252 : AOI222_X1 port map( A1 => OUT_adder_4_port, A2 => n316, B1 => 
                           LU_out_4_port, B2 => n317, C1 => SHIFT_OUT_4_port, 
                           C2 => n318, ZN => n323);
   U253 : INV_X1 port map( A => n324, ZN => OUTALU(3));
   U254 : AOI222_X1 port map( A1 => n368, A2 => n316, B1 => LU_out_3_port, B2 
                           => n317, C1 => SHIFT_OUT_3_port, C2 => n318, ZN => 
                           n324);
   U255 : INV_X1 port map( A => n325, ZN => OUTALU(31));
   U256 : AOI222_X1 port map( A1 => OUT_adder_31_port, A2 => n316, B1 => 
                           LU_out_31_port, B2 => n317, C1 => SHIFT_OUT_31_port,
                           C2 => n318, ZN => n325);
   U257 : INV_X1 port map( A => n326, ZN => OUTALU(30));
   U259 : INV_X1 port map( A => n327, ZN => OUTALU(2));
   U260 : AOI222_X1 port map( A1 => OUT_adder_2_port, A2 => n316, B1 => 
                           LU_out_2_port, B2 => n317, C1 => SHIFT_OUT_2_port, 
                           C2 => n318, ZN => n327);
   U261 : INV_X1 port map( A => n328, ZN => OUTALU(29));
   U263 : INV_X1 port map( A => n329, ZN => OUTALU(28));
   U265 : INV_X1 port map( A => n330, ZN => OUTALU(27));
   U266 : AOI222_X1 port map( A1 => n378, A2 => n316, B1 => LU_out_27_port, B2 
                           => n317, C1 => SHIFT_OUT_27_port, C2 => n318, ZN => 
                           n330);
   U267 : INV_X1 port map( A => n331, ZN => OUTALU(26));
   U269 : INV_X1 port map( A => n332, ZN => OUTALU(25));
   U270 : AOI222_X1 port map( A1 => OUT_adder_25_port, A2 => n316, B1 => 
                           LU_out_25_port, B2 => n317, C1 => SHIFT_OUT_25_port,
                           C2 => n318, ZN => n332);
   U271 : INV_X1 port map( A => n333, ZN => OUTALU(24));
   U273 : INV_X1 port map( A => n334, ZN => OUTALU(23));
   U274 : AOI222_X1 port map( A1 => OUT_adder_23_port, A2 => n316, B1 => 
                           LU_out_23_port, B2 => n317, C1 => SHIFT_OUT_23_port,
                           C2 => n318, ZN => n334);
   U275 : INV_X1 port map( A => n335, ZN => OUTALU(22));
   U276 : AOI222_X1 port map( A1 => OUT_adder_22_port, A2 => n316, B1 => 
                           LU_out_22_port, B2 => n317, C1 => SHIFT_OUT_22_port,
                           C2 => n318, ZN => n335);
   U277 : INV_X1 port map( A => n336, ZN => OUTALU(21));
   U279 : INV_X1 port map( A => n337, ZN => OUTALU(20));
   U281 : INV_X1 port map( A => n338, ZN => OUTALU(1));
   U282 : AOI222_X1 port map( A1 => OUT_adder_1_port, A2 => n316, B1 => 
                           LU_out_1_port, B2 => n317, C1 => SHIFT_OUT_1_port, 
                           C2 => n318, ZN => n338);
   U283 : INV_X1 port map( A => n339, ZN => OUTALU(19));
   U284 : AOI222_X1 port map( A1 => OUT_adder_19_port, A2 => n316, B1 => 
                           LU_out_19_port, B2 => n317, C1 => SHIFT_OUT_19_port,
                           C2 => n318, ZN => n339);
   U285 : INV_X1 port map( A => n340, ZN => OUTALU(18));
   U286 : AOI222_X1 port map( A1 => OUT_adder_18_port, A2 => n316, B1 => 
                           LU_out_18_port, B2 => n317, C1 => SHIFT_OUT_18_port,
                           C2 => n318, ZN => n340);
   U287 : INV_X1 port map( A => n341, ZN => OUTALU(17));
   U288 : AOI222_X1 port map( A1 => OUT_adder_17_port, A2 => n316, B1 => 
                           LU_out_17_port, B2 => n317, C1 => SHIFT_OUT_17_port,
                           C2 => n318, ZN => n341);
   U289 : INV_X1 port map( A => n342, ZN => OUTALU(16));
   U291 : INV_X1 port map( A => n343, ZN => OUTALU(15));
   U292 : AOI222_X1 port map( A1 => OUT_adder_15_port, A2 => n316, B1 => 
                           LU_out_15_port, B2 => n317, C1 => SHIFT_OUT_15_port,
                           C2 => n318, ZN => n343);
   U293 : INV_X1 port map( A => n344, ZN => OUTALU(14));
   U294 : AOI222_X1 port map( A1 => OUT_adder_14_port, A2 => n316, B1 => 
                           LU_out_14_port, B2 => n317, C1 => SHIFT_OUT_14_port,
                           C2 => n318, ZN => n344);
   U295 : INV_X1 port map( A => n345, ZN => OUTALU(13));
   U296 : AOI222_X1 port map( A1 => OUT_adder_13_port, A2 => n316, B1 => 
                           LU_out_13_port, B2 => n317, C1 => SHIFT_OUT_13_port,
                           C2 => n318, ZN => n345);
   U297 : INV_X1 port map( A => n346, ZN => OUTALU(12));
   U298 : AOI222_X1 port map( A1 => OUT_adder_12_port, A2 => n316, B1 => 
                           LU_out_12_port, B2 => n317, C1 => SHIFT_OUT_12_port,
                           C2 => n318, ZN => n346);
   U299 : INV_X1 port map( A => n347, ZN => OUTALU(11));
   U300 : AOI222_X1 port map( A1 => OUT_adder_11_port, A2 => n316, B1 => 
                           LU_out_11_port, B2 => n317, C1 => SHIFT_OUT_11_port,
                           C2 => n318, ZN => n347);
   U301 : INV_X1 port map( A => n348, ZN => OUTALU(10));
   U302 : AOI222_X1 port map( A1 => OUT_adder_10_port, A2 => n316, B1 => 
                           LU_out_10_port, B2 => n317, C1 => SHIFT_OUT_10_port,
                           C2 => n318, ZN => n348);
   U305 : NAND3_X1 port map( A1 => n352, A2 => n308, A3 => n353, ZN => n314);
   U309 : OAI21_X1 port map( B1 => n311, B2 => n312, A => n356, ZN => n205);
   U310 : INV_X1 port map( A => n352, ZN => n311);
   U318 : NOR2_X1 port map( A1 => FUNC(0), A2 => FUNC(1), ZN => n353);
   U321 : AOI21_X1 port map( B1 => n312, B2 => n356, A => n308, ZN => 
                           Comp_OP_0_port);
   U327 : NOR2_X1 port map( A1 => n360, A2 => FUNC(0), ZN => n355);
   U328 : INV_X1 port map( A => FUNC(1), ZN => n360);
   P4addersub_0 : P4addersub_N32 port map( A(31) => DATA1(31), A(30) => 
                           DATA1(30), A(29) => DATA1(29), A(28) => n367, A(27) 
                           => DATA1(27), A(26) => DATA1(26), A(25) => DATA1(25)
                           , A(24) => DATA1(24), A(23) => DATA1(23), A(22) => 
                           DATA1(22), A(21) => DATA1(21), A(20) => DATA1(20), 
                           A(19) => DATA1(19), A(18) => DATA1(18), A(17) => 
                           DATA1(17), A(16) => DATA1(16), A(15) => DATA1(15), 
                           A(14) => DATA1(14), A(13) => DATA1(13), A(12) => 
                           DATA1(12), A(11) => DATA1(11), A(10) => DATA1(10), 
                           A(9) => DATA1(9), A(8) => DATA1(8), A(7) => DATA1(7)
                           , A(6) => DATA1(6), A(5) => DATA1(5), A(4) => 
                           DATA1(4), A(3) => DATA1(3), A(2) => DATA1(2), A(1) 
                           => DATA1(1), A(0) => DATA1(0), B(31) => DATA2(31), 
                           B(30) => DATA2(30), B(29) => DATA2(29), B(28) => 
                           DATA2(28), B(27) => DATA2(27), B(26) => DATA2(26), 
                           B(25) => DATA2(25), B(24) => DATA2(24), B(23) => 
                           DATA2(23), B(22) => DATA2(22), B(21) => DATA2(21), 
                           B(20) => DATA2(20), B(19) => DATA2(19), B(18) => 
                           DATA2(18), B(17) => DATA2(17), B(16) => DATA2(16), 
                           B(15) => DATA2(15), B(14) => DATA2(14), B(13) => 
                           DATA2(13), B(12) => DATA2(12), B(11) => DATA2(11), 
                           B(10) => DATA2(10), B(9) => DATA2(9), B(8) => 
                           DATA2(8), B(7) => DATA2(7), B(6) => DATA2(6), B(5) 
                           => DATA2(5), B(4) => DATA2(4), B(3) => DATA2(3), 
                           B(2) => DATA2(2), B(1) => DATA2(1), B(0) => DATA2(0)
                           , sub_add => n305, Y(31) => OUT_adder_31_port, Y(30)
                           => OUT_adder_30_port, Y(29) => OUT_adder_29_port, 
                           Y(28) => OUT_adder_28_port, Y(27) => 
                           OUT_adder_27_port, Y(26) => OUT_adder_26_port, Y(25)
                           => OUT_adder_25_port, Y(24) => OUT_adder_24_port, 
                           Y(23) => OUT_adder_23_port, Y(22) => 
                           OUT_adder_22_port, Y(21) => OUT_adder_21_port, Y(20)
                           => OUT_adder_20_port, Y(19) => OUT_adder_19_port, 
                           Y(18) => OUT_adder_18_port, Y(17) => 
                           OUT_adder_17_port, Y(16) => OUT_adder_16_port, Y(15)
                           => OUT_adder_15_port, Y(14) => OUT_adder_14_port, 
                           Y(13) => OUT_adder_13_port, Y(12) => 
                           OUT_adder_12_port, Y(11) => OUT_adder_11_port, Y(10)
                           => OUT_adder_10_port, Y(9) => OUT_adder_9_port, Y(8)
                           => OUT_adder_8_port, Y(7) => OUT_adder_7_port, Y(6) 
                           => OUT_adder_6_port, Y(5) => OUT_adder_5_port, Y(4) 
                           => OUT_adder_4_port, Y(3) => OUT_adder_3_port, Y(2) 
                           => OUT_adder_2_port, Y(1) => OUT_adder_1_port, Y(0) 
                           => OUT_adder_0_port, Cout => Adder_Cout);
   logicunit_0 : logicunit port map( A(31) => DATA1(31), A(30) => DATA1(30), 
                           A(29) => DATA1(29), A(28) => n367, A(27) => 
                           DATA1(27), A(26) => DATA1(26), A(25) => DATA1(25), 
                           A(24) => DATA1(24), A(23) => n366, A(22) => 
                           DATA1(22), A(21) => DATA1(21), A(20) => DATA1(20), 
                           A(19) => DATA1(19), A(18) => DATA1(18), A(17) => 
                           DATA1(17), A(16) => DATA1(16), A(15) => n375, A(14) 
                           => DATA1(14), A(13) => n369, A(12) => DATA1(12), 
                           A(11) => n373, A(10) => DATA1(10), A(9) => n374, 
                           A(8) => DATA1(8), A(7) => n370, A(6) => DATA1(6), 
                           A(5) => n372, A(4) => DATA1(4), A(3) => n376, A(2) 
                           => DATA1(2), A(1) => n371, A(0) => n377, B(31) => 
                           DATA2(31), B(30) => DATA2(30), B(29) => DATA2(29), 
                           B(28) => DATA2(28), B(27) => DATA2(27), B(26) => 
                           DATA2(26), B(25) => DATA2(25), B(24) => DATA2(24), 
                           B(23) => DATA2(23), B(22) => DATA2(22), B(21) => 
                           DATA2(21), B(20) => DATA2(20), B(19) => DATA2(19), 
                           B(18) => DATA2(18), B(17) => DATA2(17), B(16) => 
                           DATA2(16), B(15) => DATA2(15), B(14) => DATA2(14), 
                           B(13) => DATA2(13), B(12) => DATA2(12), B(11) => 
                           DATA2(11), B(10) => DATA2(10), B(9) => DATA2(9), 
                           B(8) => DATA2(8), B(7) => DATA2(7), B(6) => DATA2(6)
                           , B(5) => DATA2(5), B(4) => DATA2(4), B(3) => 
                           DATA2(3), B(2) => DATA2(2), B(1) => DATA2(1), B(0) 
                           => DATA2(0), SEL(2) => Sel_2_port, SEL(1) => n306, 
                           SEL(0) => n306, LU_OUT(31) => LU_out_31_port, 
                           LU_OUT(30) => LU_out_30_port, LU_OUT(29) => 
                           LU_out_29_port, LU_OUT(28) => LU_out_28_port, 
                           LU_OUT(27) => LU_out_27_port, LU_OUT(26) => 
                           LU_out_26_port, LU_OUT(25) => LU_out_25_port, 
                           LU_OUT(24) => LU_out_24_port, LU_OUT(23) => 
                           LU_out_23_port, LU_OUT(22) => LU_out_22_port, 
                           LU_OUT(21) => LU_out_21_port, LU_OUT(20) => 
                           LU_out_20_port, LU_OUT(19) => LU_out_19_port, 
                           LU_OUT(18) => LU_out_18_port, LU_OUT(17) => 
                           LU_out_17_port, LU_OUT(16) => LU_out_16_port, 
                           LU_OUT(15) => LU_out_15_port, LU_OUT(14) => 
                           LU_out_14_port, LU_OUT(13) => LU_out_13_port, 
                           LU_OUT(12) => LU_out_12_port, LU_OUT(11) => 
                           LU_out_11_port, LU_OUT(10) => LU_out_10_port, 
                           LU_OUT(9) => LU_out_9_port, LU_OUT(8) => 
                           LU_out_8_port, LU_OUT(7) => LU_out_7_port, LU_OUT(6)
                           => LU_out_6_port, LU_OUT(5) => LU_out_5_port, 
                           LU_OUT(4) => LU_out_4_port, LU_OUT(3) => 
                           LU_out_3_port, LU_OUT(2) => LU_out_2_port, LU_OUT(1)
                           => LU_out_1_port, LU_OUT(0) => LU_out_0_port);
   ComparatorUnit_0 : ComparatorUnit port map( A_MSB => DATA1(31), B_MSB => 
                           DATA2(31), SUBIN(31) => OUT_adder_31_port, SUBIN(30)
                           => OUT_adder_30_port, SUBIN(29) => OUT_adder_29_port
                           , SUBIN(28) => OUT_adder_28_port, SUBIN(27) => 
                           OUT_adder_27_port, SUBIN(26) => OUT_adder_26_port, 
                           SUBIN(25) => OUT_adder_25_port, SUBIN(24) => 
                           OUT_adder_24_port, SUBIN(23) => OUT_adder_23_port, 
                           SUBIN(22) => OUT_adder_22_port, SUBIN(21) => 
                           OUT_adder_21_port, SUBIN(20) => OUT_adder_20_port, 
                           SUBIN(19) => OUT_adder_19_port, SUBIN(18) => 
                           OUT_adder_18_port, SUBIN(17) => OUT_adder_17_port, 
                           SUBIN(16) => OUT_adder_16_port, SUBIN(15) => 
                           OUT_adder_15_port, SUBIN(14) => OUT_adder_14_port, 
                           SUBIN(13) => OUT_adder_13_port, SUBIN(12) => 
                           OUT_adder_12_port, SUBIN(11) => OUT_adder_11_port, 
                           SUBIN(10) => OUT_adder_10_port, SUBIN(9) => 
                           OUT_adder_9_port, SUBIN(8) => OUT_adder_8_port, 
                           SUBIN(7) => OUT_adder_7_port, SUBIN(6) => 
                           OUT_adder_6_port, SUBIN(5) => OUT_adder_5_port, 
                           SUBIN(4) => OUT_adder_4_port, SUBIN(3) => 
                           OUT_adder_3_port, SUBIN(2) => OUT_adder_2_port, 
                           SUBIN(1) => OUT_adder_1_port, SUBIN(0) => 
                           OUT_adder_0_port, COUT => Adder_Cout, SIGN_UNSIGN =>
                           sign_unsign, OP(0) => n205, OP(1) => Comp_OP_1_port,
                           OP(2) => Comp_OP_0_port, CU_OUT(31) => net126648, 
                           CU_OUT(30) => net126649, CU_OUT(29) => net126650, 
                           CU_OUT(28) => net126651, CU_OUT(27) => net126652, 
                           CU_OUT(26) => net126653, CU_OUT(25) => net126654, 
                           CU_OUT(24) => net126655, CU_OUT(23) => net126656, 
                           CU_OUT(22) => net126657, CU_OUT(21) => net126658, 
                           CU_OUT(20) => net126659, CU_OUT(19) => net126660, 
                           CU_OUT(18) => net126661, CU_OUT(17) => net126662, 
                           CU_OUT(16) => net126663, CU_OUT(15) => net126664, 
                           CU_OUT(14) => net126665, CU_OUT(13) => net126666, 
                           CU_OUT(12) => net126667, CU_OUT(11) => net126668, 
                           CU_OUT(10) => net126669, CU_OUT(9) => net126670, 
                           CU_OUT(8) => net126671, CU_OUT(7) => net126672, 
                           CU_OUT(6) => net126673, CU_OUT(5) => net126674, 
                           CU_OUT(4) => net126675, CU_OUT(3) => net126676, 
                           CU_OUT(2) => net126677, CU_OUT(1) => net126678, 
                           CU_OUT(0) => CU_OUT_0_port);
   shifter_0 : shifter port map( R(31) => DATA1(31), R(30) => DATA1(30), R(29) 
                           => DATA1(29), R(28) => n367, R(27) => DATA1(27), 
                           R(26) => DATA1(26), R(25) => DATA1(25), R(24) => 
                           DATA1(24), R(23) => n366, R(22) => DATA1(22), R(21) 
                           => DATA1(21), R(20) => DATA1(20), R(19) => DATA1(19)
                           , R(18) => DATA1(18), R(17) => DATA1(17), R(16) => 
                           DATA1(16), R(15) => n375, R(14) => DATA1(14), R(13) 
                           => n369, R(12) => DATA1(12), R(11) => n373, R(10) =>
                           DATA1(10), R(9) => n374, R(8) => DATA1(8), R(7) => 
                           n370, R(6) => DATA1(6), R(5) => n372, R(4) => 
                           DATA1(4), R(3) => n376, R(2) => DATA1(2), R(1) => 
                           n371, R(0) => n377, Offset(4) => DATA2(4), Offset(3)
                           => DATA2(3), Offset(2) => DATA2(2), Offset(1) => 
                           DATA2(1), Offset(0) => DATA2(0), Conf(0) => 
                           Conf_1_port, Conf(1) => Conf_0_port, Shift_OUT(31) 
                           => SHIFT_OUT_31_port, Shift_OUT(30) => 
                           SHIFT_OUT_30_port, Shift_OUT(29) => 
                           SHIFT_OUT_29_port, Shift_OUT(28) => 
                           SHIFT_OUT_28_port, Shift_OUT(27) => 
                           SHIFT_OUT_27_port, Shift_OUT(26) => 
                           SHIFT_OUT_26_port, Shift_OUT(25) => 
                           SHIFT_OUT_25_port, Shift_OUT(24) => 
                           SHIFT_OUT_24_port, Shift_OUT(23) => 
                           SHIFT_OUT_23_port, Shift_OUT(22) => 
                           SHIFT_OUT_22_port, Shift_OUT(21) => 
                           SHIFT_OUT_21_port, Shift_OUT(20) => 
                           SHIFT_OUT_20_port, Shift_OUT(19) => 
                           SHIFT_OUT_19_port, Shift_OUT(18) => 
                           SHIFT_OUT_18_port, Shift_OUT(17) => 
                           SHIFT_OUT_17_port, Shift_OUT(16) => 
                           SHIFT_OUT_16_port, Shift_OUT(15) => 
                           SHIFT_OUT_15_port, Shift_OUT(14) => 
                           SHIFT_OUT_14_port, Shift_OUT(13) => 
                           SHIFT_OUT_13_port, Shift_OUT(12) => 
                           SHIFT_OUT_12_port, Shift_OUT(11) => 
                           SHIFT_OUT_11_port, Shift_OUT(10) => 
                           SHIFT_OUT_10_port, Shift_OUT(9) => SHIFT_OUT_9_port,
                           Shift_OUT(8) => SHIFT_OUT_8_port, Shift_OUT(7) => 
                           SHIFT_OUT_7_port, Shift_OUT(6) => SHIFT_OUT_6_port, 
                           Shift_OUT(5) => SHIFT_OUT_5_port, Shift_OUT(4) => 
                           SHIFT_OUT_4_port, Shift_OUT(3) => SHIFT_OUT_3_port, 
                           Shift_OUT(2) => SHIFT_OUT_2_port, Shift_OUT(1) => 
                           SHIFT_OUT_1_port, Shift_OUT(0) => SHIFT_OUT_0_port);
   U326 : INV_X1 port map( A => n355, ZN => n312);
   U320 : NAND2_X1 port map( A1 => FUNC(3), A2 => n355, ZN => n310);
   U240 : INV_X1 port map( A => n313, ZN => Sel_2_port);
   U239 : OAI21_X1 port map( B1 => n308, B2 => n313, A => n314, ZN => n104);
   U322 : INV_X1 port map( A => FUNC(4), ZN => n308);
   U317 : NAND3_X1 port map( A1 => n353, A2 => FUNC(2), A3 => FUNC(3), ZN => 
                           n358);
   U238 : OAI22_X1 port map( A1 => FUNC(2), A2 => n310, B1 => n311, B2 => n312,
                           ZN => sign_unsign);
   U315 : NOR2_X1 port map( A1 => n308, A2 => n358, ZN => Conf_1_port);
   U316 : NOR2_X1 port map( A1 => FUNC(4), A2 => n358, ZN => Conf_0_port);
   U308 : NOR2_X1 port map( A1 => n355, A2 => n205, ZN => n309);
   U235 : NAND2_X2 port map( A1 => n313, A2 => n314, ZN => n317);
   U325 : INV_X1 port map( A => FUNC(3), ZN => n357);
   U306 : NAND3_X1 port map( A1 => n353, A2 => n354, A3 => FUNC(3), ZN => n313)
                           ;
   U311 : NOR2_X1 port map( A1 => n354, A2 => FUNC(3), ZN => n352);
   U323 : NAND4_X1 port map( A1 => FUNC(0), A2 => n357, A3 => n354, A4 => n360,
                           ZN => n356);
   U324 : INV_X1 port map( A => FUNC(2), ZN => n354);
   U237 : OAI21_X1 port map( B1 => n307, B2 => n308, A => n309, ZN => sub_add);
   U313 : NAND3_X1 port map( A1 => n357, A2 => n354, A3 => n353, ZN => n307);
   U314 : NAND3_X1 port map( A1 => n353, A2 => FUNC(2), A3 => FUNC(4), ZN => 
                           n359);
   U234 : NAND2_X2 port map( A1 => n358, A2 => n359, ZN => n318);
   U236 : INV_X2 port map( A => n307, ZN => n316);
   U312 : AOI22_X1 port map( A1 => SHIFT_OUT_0_port, A2 => n318, B1 => 
                           OUT_adder_0_port, B2 => n316, ZN => n349);
   U232 : AOI222_X4 port map( A1 => OUT_adder_28_port, A2 => n316, B1 => 
                           LU_out_28_port, B2 => n317, C1 => SHIFT_OUT_28_port,
                           C2 => n318, ZN => n329);
   U258 : CLKBUF_X1 port map( A => OUT_adder_26_port, Z => n364);
   U262 : OAI221_X1 port map( B1 => n361, B2 => n362, C1 => n363, C2 => n309, A
                           => n349, ZN => OUTALU(0));
   U264 : INV_X1 port map( A => LU_out_0_port, ZN => n361);
   U268 : INV_X1 port map( A => n317, ZN => n362);
   U272 : INV_X1 port map( A => CU_OUT_0_port, ZN => n363);
   U278 : CLKBUF_X1 port map( A => OUT_adder_16_port, Z => n365);
   U280 : AOI222_X4 port map( A1 => n364, A2 => n316, B1 => LU_out_26_port, B2 
                           => n317, C1 => SHIFT_OUT_26_port, C2 => n318, ZN => 
                           n331);
   U290 : AOI222_X4 port map( A1 => n365, A2 => n316, B1 => LU_out_16_port, B2 
                           => n317, C1 => SHIFT_OUT_16_port, C2 => n318, ZN => 
                           n342);
   U303 : CLKBUF_X1 port map( A => DATA1(23), Z => n366);
   U304 : BUF_X2 port map( A => DATA1(28), Z => n367);
   U307 : AOI222_X4 port map( A1 => OUT_adder_21_port, A2 => n316, B1 => 
                           LU_out_21_port, B2 => n317, C1 => SHIFT_OUT_21_port,
                           C2 => n318, ZN => n336);
   U319 : AOI222_X4 port map( A1 => OUT_adder_29_port, A2 => n316, B1 => 
                           LU_out_29_port, B2 => n317, C1 => SHIFT_OUT_29_port,
                           C2 => n318, ZN => n328);
   U329 : CLKBUF_X1 port map( A => OUT_adder_30_port, Z => n379);
   U330 : CLKBUF_X1 port map( A => OUT_adder_3_port, Z => n368);
   U331 : CLKBUF_X1 port map( A => DATA1(13), Z => n369);
   U332 : CLKBUF_X1 port map( A => DATA1(7), Z => n370);
   U333 : CLKBUF_X1 port map( A => DATA1(1), Z => n371);
   U334 : CLKBUF_X1 port map( A => DATA1(5), Z => n372);
   U335 : CLKBUF_X1 port map( A => DATA1(11), Z => n373);
   U336 : CLKBUF_X1 port map( A => DATA1(9), Z => n374);
   U337 : CLKBUF_X1 port map( A => DATA1(15), Z => n375);
   U338 : CLKBUF_X1 port map( A => DATA1(3), Z => n376);
   U339 : INV_X2 port map( A => n310, ZN => Comp_OP_1_port);
   U340 : CLKBUF_X1 port map( A => DATA1(0), Z => n377);
   U341 : AOI222_X4 port map( A1 => OUT_adder_24_port, A2 => n316, B1 => 
                           LU_out_24_port, B2 => n317, C1 => SHIFT_OUT_24_port,
                           C2 => n318, ZN => n333);
   U342 : AOI222_X4 port map( A1 => OUT_adder_20_port, A2 => n316, B1 => 
                           LU_out_20_port, B2 => n317, C1 => SHIFT_OUT_20_port,
                           C2 => n318, ZN => n337);
   U343 : CLKBUF_X1 port map( A => OUT_adder_27_port, Z => n378);
   U344 : AOI222_X4 port map( A1 => n379, A2 => n316, B1 => LU_out_30_port, B2 
                           => n317, C1 => SHIFT_OUT_30_port, C2 => n318, ZN => 
                           n326);
   U345 : BUF_X8 port map( A => sub_add, Z => n305);

end SYN_STRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P4addersub_N32 is

   port( A, B : in std_logic_vector (31 downto 0);  sub_add : in std_logic;  Y 
         : out std_logic_vector (31 downto 0);  Cout : out std_logic);

end P4addersub_N32;

architecture SYN_struct_architecture of P4addersub_N32 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component sumgen_N_blocks8
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector
            (7 downto 0);  S : out std_logic_vector (31 downto 0));
   end component;
   
   component STCG_N32_L5
      port( A, B : in std_logic_vector (31 downto 0);  cin : in std_logic;  
            cout : out std_logic_vector (7 downto 0));
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal B_subadd_31_port, B_subadd_30_port, B_subadd_29_port, 
      B_subadd_26_port, B_subadd_25_port, B_subadd_4_port, carry_7_port, 
      carry_6_port, carry_5_port, carry_4_port, carry_3_port, carry_2_port, 
      carry_1_port, net6007, net6009, net6012, net6021, net6024, n1, n2, n3, n4
      , n5, n6, n7, n8, n9, n10, n11, n13, n14, n15, n16, n19, n21, n22, n25, 
      n26, n38, n43, n44, n45, n46, n47, n48, n49, n50, n51 : std_logic;

begin
   
   U65 : XOR2_X1 port map( A => sub_add, B => B(13), Z => net6024);
   U66 : XOR2_X1 port map( A => sub_add, B => B(23), Z => net6021);
   U67 : XOR2_X1 port map( A => sub_add, B => B(7), Z => net6012);
   U68 : XOR2_X1 port map( A => sub_add, B => B(11), Z => net6009);
   U69 : XOR2_X1 port map( A => sub_add, B => B(15), Z => net6007);
   U70 : XOR2_X1 port map( A => sub_add, B => B(17), Z => n9);
   U71 : XOR2_X1 port map( A => sub_add, B => B(20), Z => n8);
   U72 : XOR2_X1 port map( A => sub_add, B => B(1), Z => n7);
   U73 : XOR2_X1 port map( A => sub_add, B => B(22), Z => n6);
   U74 : XOR2_X1 port map( A => sub_add, B => B(8), Z => n5);
   U75 : XOR2_X1 port map( A => sub_add, B => B(14), Z => n4);
   U76 : XOR2_X1 port map( A => sub_add, B => B(0), Z => n38);
   U77 : XOR2_X1 port map( A => sub_add, B => B(10), Z => n3);
   U78 : XOR2_X1 port map( A => sub_add, B => B(19), Z => n26);
   U79 : XOR2_X1 port map( A => sub_add, B => B(16), Z => n25);
   U80 : XOR2_X1 port map( A => sub_add, B => B(5), Z => n22);
   U81 : XOR2_X1 port map( A => sub_add, B => B(9), Z => n21);
   U82 : XOR2_X1 port map( A => sub_add, B => B(6), Z => n2);
   U83 : XOR2_X1 port map( A => sub_add, B => B(27), Z => n19);
   U84 : XOR2_X1 port map( A => sub_add, B => B(3), Z => n16);
   U85 : XOR2_X1 port map( A => sub_add, B => B(2), Z => n15);
   U86 : XOR2_X1 port map( A => sub_add, B => B(24), Z => n14);
   U87 : XOR2_X1 port map( A => sub_add, B => B(18), Z => n13);
   U88 : XOR2_X1 port map( A => sub_add, B => B(21), Z => n11);
   U89 : XOR2_X1 port map( A => sub_add, B => B(12), Z => n10);
   U90 : XOR2_X1 port map( A => sub_add, B => B(28), Z => n1);
   U91 : XOR2_X1 port map( A => sub_add, B => B(4), Z => B_subadd_4_port);
   U92 : XOR2_X1 port map( A => sub_add, B => B(31), Z => B_subadd_31_port);
   U93 : XOR2_X1 port map( A => sub_add, B => B(30), Z => B_subadd_30_port);
   U94 : XOR2_X1 port map( A => sub_add, B => B(29), Z => B_subadd_29_port);
   U95 : XOR2_X1 port map( A => sub_add, B => B(26), Z => B_subadd_26_port);
   U96 : XOR2_X1 port map( A => sub_add, B => B(25), Z => B_subadd_25_port);
   STCG_1 : STCG_N32_L5 port map( A(31) => A(31), A(30) => A(30), A(29) => 
                           A(29), A(28) => A(28), A(27) => A(27), A(26) => 
                           A(26), A(25) => A(25), A(24) => A(24), A(23) => 
                           A(23), A(22) => A(22), A(21) => A(21), A(20) => 
                           A(20), A(19) => A(19), A(18) => A(18), A(17) => 
                           A(17), A(16) => A(16), A(15) => A(15), A(14) => 
                           A(14), A(13) => A(13), A(12) => A(12), A(11) => 
                           A(11), A(10) => A(10), A(9) => A(9), A(8) => A(8), 
                           A(7) => A(7), A(6) => A(6), A(5) => A(5), A(4) => 
                           A(4), A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(31) => B_subadd_31_port, B(30) => 
                           B_subadd_30_port, B(29) => B_subadd_29_port, B(28) 
                           => n1, B(27) => n19, B(26) => B_subadd_26_port, 
                           B(25) => B_subadd_25_port, B(24) => n14, B(23) => 
                           net6021, B(22) => n6, B(21) => n11, B(20) => n8, 
                           B(19) => n26, B(18) => n13, B(17) => n9, B(16) => 
                           n25, B(15) => net6007, B(14) => n4, B(13) => net6024
                           , B(12) => n10, B(11) => net6009, B(10) => n3, B(9) 
                           => n21, B(8) => n5, B(7) => net6012, B(6) => n2, 
                           B(5) => n22, B(4) => B_subadd_4_port, B(3) => n16, 
                           B(2) => n15, B(1) => n7, B(0) => n38, cin => sub_add
                           , cout(7) => Cout, cout(6) => carry_7_port, cout(5) 
                           => carry_6_port, cout(4) => carry_5_port, cout(3) =>
                           carry_4_port, cout(2) => carry_3_port, cout(1) => 
                           carry_2_port, cout(0) => carry_1_port);
   sumgen_1 : sumgen_N_blocks8 port map( A(31) => A(31), A(30) => A(30), A(29) 
                           => A(29), A(28) => A(28), A(27) => A(27), A(26) => 
                           A(26), A(25) => A(25), A(24) => A(24), A(23) => 
                           A(23), A(22) => A(22), A(21) => A(21), A(20) => 
                           A(20), A(19) => A(19), A(18) => A(18), A(17) => 
                           A(17), A(16) => A(16), A(15) => n50, A(14) => A(14),
                           A(13) => n46, A(12) => A(12), A(11) => n47, A(10) =>
                           A(10), A(9) => n45, A(8) => A(8), A(7) => n49, A(6) 
                           => A(6), A(5) => n44, A(4) => A(4), A(3) => n48, 
                           A(2) => A(2), A(1) => n43, A(0) => n51, B(31) => 
                           B_subadd_31_port, B(30) => B_subadd_30_port, B(29) 
                           => B_subadd_29_port, B(28) => n1, B(27) => n19, 
                           B(26) => B_subadd_26_port, B(25) => B_subadd_25_port
                           , B(24) => n14, B(23) => net6021, B(22) => n6, B(21)
                           => n11, B(20) => n8, B(19) => n26, B(18) => n13, 
                           B(17) => n9, B(16) => n25, B(15) => net6007, B(14) 
                           => n4, B(13) => net6024, B(12) => n10, B(11) => 
                           net6009, B(10) => n3, B(9) => n21, B(8) => n5, B(7) 
                           => net6012, B(6) => n2, B(5) => n22, B(4) => 
                           B_subadd_4_port, B(3) => n16, B(2) => n15, B(1) => 
                           n7, B(0) => n38, Ci(7) => carry_7_port, Ci(6) => 
                           carry_6_port, Ci(5) => carry_5_port, Ci(4) => 
                           carry_4_port, Ci(3) => carry_3_port, Ci(2) => 
                           carry_2_port, Ci(1) => carry_1_port, Ci(0) => 
                           sub_add, S(31) => Y(31), S(30) => Y(30), S(29) => 
                           Y(29), S(28) => Y(28), S(27) => Y(27), S(26) => 
                           Y(26), S(25) => Y(25), S(24) => Y(24), S(23) => 
                           Y(23), S(22) => Y(22), S(21) => Y(21), S(20) => 
                           Y(20), S(19) => Y(19), S(18) => Y(18), S(17) => 
                           Y(17), S(16) => Y(16), S(15) => Y(15), S(14) => 
                           Y(14), S(13) => Y(13), S(12) => Y(12), S(11) => 
                           Y(11), S(10) => Y(10), S(9) => Y(9), S(8) => Y(8), 
                           S(7) => Y(7), S(6) => Y(6), S(5) => Y(5), S(4) => 
                           Y(4), S(3) => Y(3), S(2) => Y(2), S(1) => Y(1), S(0)
                           => Y(0));
   U97 : BUF_X2 port map( A => A(9), Z => n45);
   U98 : CLKBUF_X1 port map( A => A(1), Z => n43);
   U99 : CLKBUF_X1 port map( A => A(5), Z => n44);
   U100 : CLKBUF_X1 port map( A => A(13), Z => n46);
   U101 : CLKBUF_X1 port map( A => A(11), Z => n47);
   U102 : BUF_X2 port map( A => A(0), Z => n51);
   U103 : CLKBUF_X1 port map( A => A(3), Z => n48);
   U104 : CLKBUF_X1 port map( A => A(7), Z => n49);
   U105 : CLKBUF_X1 port map( A => A(15), Z => n50);

end SYN_struct_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity HazardUnit_NUMBIT32_ADDRESS_WIDTH_RF5_OP_CODE_SIZE6 is

   port( CLK, RST : in std_logic;  RS1, RS2 : in std_logic_vector (4 downto 0);
         REGWRITE_DX, MEMREAD_DX : in std_logic;  RD : in std_logic_vector (4 
         downto 0);  OPCODE : in std_logic_vector (5 downto 0);  STALL : out 
         std_logic);

end HazardUnit_NUMBIT32_ADDRESS_WIDTH_RF5_OP_CODE_SIZE6;

architecture SYN_beh of HazardUnit_NUMBIT32_ADDRESS_WIDTH_RF5_OP_CODE_SIZE6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N9, N10, N11, N12, N13, n1, n2, n3, n4, n5, n6, n7, n8, n9_port, 
      n10_port, n11_port, n12_port, n13_port, n14, n15, n16, n17, n18, n19, n20
      , n21, n22, n23, n24, net114859, net114860, net114861 : std_logic;

begin
   
   RD_DX_reg_4_inst : DFF_X1 port map( D => N13, CK => CLK, Q => net114861, QN 
                           => n6);
   RD_DX_reg_3_inst : DFF_X1 port map( D => N12, CK => CLK, Q => net114860, QN 
                           => n5);
   RD_DX_reg_2_inst : DFF_X1 port map( D => N11, CK => CLK, Q => net114859, QN 
                           => n9_port);
   RD_DX_reg_1_inst : DFF_X1 port map( D => N10, CK => CLK, Q => n2, QN => n8);
   RD_DX_reg_0_inst : DFF_X1 port map( D => N9, CK => CLK, Q => n1, QN => n7);
   U3 : AND2_X1 port map( A1 => n3, A2 => n4, ZN => n18);
   U4 : XOR2_X1 port map( A => n6, B => RS1(4), Z => n3);
   U5 : XOR2_X1 port map( A => RS1(2), B => n9_port, Z => n4);
   U6 : AND4_X2 port map( A1 => n15, A2 => n16, A3 => n17, A4 => n18, ZN => 
                           n12_port);
   U7 : NAND2_X1 port map( A1 => n10_port, A2 => n11_port, ZN => STALL);
   U8 : NAND4_X1 port map( A1 => OPCODE(2), A2 => n12_port, A3 => REGWRITE_DX, 
                           A4 => n13_port, ZN => n11_port);
   U9 : NOR4_X1 port map( A1 => OPCODE(5), A2 => OPCODE(4), A3 => OPCODE(3), A4
                           => OPCODE(1), ZN => n13_port);
   U10 : OAI21_X1 port map( B1 => n14, B2 => n12_port, A => MEMREAD_DX, ZN => 
                           n10_port);
   U11 : XOR2_X1 port map( A => n7, B => RS1(0), Z => n17);
   U12 : XOR2_X1 port map( A => n8, B => RS1(1), Z => n16);
   U13 : XOR2_X1 port map( A => n5, B => RS1(3), Z => n15);
   U14 : NOR3_X1 port map( A1 => n19, A2 => n20, A3 => n21, ZN => n14);
   U15 : XNOR2_X1 port map( A => n6, B => RS2(4), ZN => n21);
   U16 : XNOR2_X1 port map( A => n9_port, B => RS2(2), ZN => n20);
   U17 : NAND3_X1 port map( A1 => n22, A2 => n23, A3 => n24, ZN => n19);
   U18 : XOR2_X1 port map( A => n7, B => RS2(0), Z => n24);
   U19 : XOR2_X1 port map( A => n8, B => RS2(1), Z => n23);
   U20 : XOR2_X1 port map( A => n5, B => RS2(3), Z => n22);
   U21 : AND2_X1 port map( A1 => RST, A2 => RD(0), ZN => N9);
   U22 : AND2_X1 port map( A1 => RD(4), A2 => RST, ZN => N13);
   U23 : AND2_X1 port map( A1 => RD(3), A2 => RST, ZN => N12);
   U24 : AND2_X1 port map( A1 => RD(2), A2 => RST, ZN => N11);
   U25 : AND2_X1 port map( A1 => RD(1), A2 => RST, ZN => N10);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity BTB_PC_SIZE32_BTBSIZE5 is

   port( Reset, Clk, Enable : in std_logic;  PC_read : in std_logic_vector (31 
         downto 0);  WR : in std_logic;  PC_write : in std_logic_vector (31 
         downto 0);  SetT_NT : in std_logic;  Set_target : in std_logic_vector 
         (31 downto 0);  OUT_PC_target : out std_logic_vector (31 downto 0);  
         OUTT_NT, prevT_NT : out std_logic);

end BTB_PC_SIZE32_BTBSIZE5;

architecture SYN_Behavioral of BTB_PC_SIZE32_BTBSIZE5 is

   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component BTB_PC_SIZE32_BTBSIZE5_DW01_cmp6_0
      port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, 
            GT, EQ, LE, GE, NE : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X8
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X2
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal OUTT_NT_port, prevT_NT_port, pc_target_2_31_port, pc_target_2_30_port
      , pc_target_2_29_port, pc_target_2_28_port, pc_target_2_27_port, 
      pc_target_2_26_port, pc_target_2_25_port, pc_target_2_24_port, 
      pc_target_2_23_port, pc_target_2_22_port, pc_target_2_21_port, 
      pc_target_2_20_port, pc_target_2_19_port, pc_target_2_18_port, 
      pc_target_2_17_port, pc_target_2_16_port, pc_target_2_15_port, 
      pc_target_2_14_port, pc_target_2_13_port, pc_target_2_12_port, 
      pc_target_2_11_port, pc_target_2_10_port, pc_target_2_9_port, 
      pc_target_2_8_port, pc_target_2_7_port, pc_target_2_6_port, 
      pc_target_2_5_port, pc_target_2_4_port, pc_target_2_3_port, 
      pc_target_2_2_port, pc_target_2_1_port, pc_target_2_0_port, 
      pc_target_3_31_port, pc_target_3_30_port, pc_target_3_29_port, 
      pc_target_3_28_port, pc_target_3_27_port, pc_target_3_26_port, 
      pc_target_3_25_port, pc_target_3_24_port, pc_target_3_23_port, 
      pc_target_3_22_port, pc_target_3_21_port, pc_target_3_20_port, 
      pc_target_3_19_port, pc_target_3_18_port, pc_target_3_17_port, 
      pc_target_3_16_port, pc_target_3_15_port, pc_target_3_14_port, 
      pc_target_3_13_port, pc_target_3_12_port, pc_target_3_11_port, 
      pc_target_3_10_port, pc_target_3_9_port, pc_target_3_8_port, 
      pc_target_3_7_port, pc_target_3_6_port, pc_target_3_5_port, 
      pc_target_3_4_port, pc_target_3_3_port, pc_target_3_2_port, 
      pc_target_3_1_port, pc_target_3_0_port, pc_target_6_31_port, 
      pc_target_6_30_port, pc_target_6_29_port, pc_target_6_28_port, 
      pc_target_6_27_port, pc_target_6_26_port, pc_target_6_25_port, 
      pc_target_6_24_port, pc_target_6_23_port, pc_target_6_22_port, 
      pc_target_6_21_port, pc_target_6_20_port, pc_target_6_19_port, 
      pc_target_6_18_port, pc_target_6_17_port, pc_target_6_16_port, 
      pc_target_6_15_port, pc_target_6_14_port, pc_target_6_13_port, 
      pc_target_6_12_port, pc_target_6_11_port, pc_target_6_10_port, 
      pc_target_6_9_port, pc_target_6_8_port, pc_target_6_7_port, 
      pc_target_6_6_port, pc_target_6_5_port, pc_target_6_4_port, 
      pc_target_6_3_port, pc_target_6_2_port, pc_target_6_1_port, 
      pc_target_6_0_port, pc_target_7_31_port, pc_target_7_30_port, 
      pc_target_7_29_port, pc_target_7_28_port, pc_target_7_27_port, 
      pc_target_7_26_port, pc_target_7_25_port, pc_target_7_24_port, 
      pc_target_7_23_port, pc_target_7_22_port, pc_target_7_21_port, 
      pc_target_7_20_port, pc_target_7_19_port, pc_target_7_18_port, 
      pc_target_7_17_port, pc_target_7_16_port, pc_target_7_15_port, 
      pc_target_7_14_port, pc_target_7_13_port, pc_target_7_12_port, 
      pc_target_7_11_port, pc_target_7_10_port, pc_target_7_9_port, 
      pc_target_7_8_port, pc_target_7_7_port, pc_target_7_6_port, 
      pc_target_7_5_port, pc_target_7_4_port, pc_target_7_3_port, 
      pc_target_7_2_port, pc_target_7_1_port, pc_target_7_0_port, 
      pc_target_10_31_port, pc_target_10_30_port, pc_target_10_29_port, 
      pc_target_10_28_port, pc_target_10_27_port, pc_target_10_26_port, 
      pc_target_10_25_port, pc_target_10_24_port, pc_target_10_23_port, 
      pc_target_10_22_port, pc_target_10_21_port, pc_target_10_20_port, 
      pc_target_10_19_port, pc_target_10_18_port, pc_target_10_17_port, 
      pc_target_10_16_port, pc_target_10_15_port, pc_target_10_14_port, 
      pc_target_10_13_port, pc_target_10_12_port, pc_target_10_11_port, 
      pc_target_10_10_port, pc_target_10_9_port, pc_target_10_8_port, 
      pc_target_10_7_port, pc_target_10_6_port, pc_target_10_5_port, 
      pc_target_10_4_port, pc_target_10_3_port, pc_target_10_2_port, 
      pc_target_10_1_port, pc_target_10_0_port, pc_target_11_31_port, 
      pc_target_11_30_port, pc_target_11_29_port, pc_target_11_28_port, 
      pc_target_11_27_port, pc_target_11_26_port, pc_target_11_25_port, 
      pc_target_11_24_port, pc_target_11_23_port, pc_target_11_22_port, 
      pc_target_11_21_port, pc_target_11_20_port, pc_target_11_19_port, 
      pc_target_11_18_port, pc_target_11_17_port, pc_target_11_16_port, 
      pc_target_11_15_port, pc_target_11_14_port, pc_target_11_13_port, 
      pc_target_11_12_port, pc_target_11_11_port, pc_target_11_10_port, 
      pc_target_11_9_port, pc_target_11_8_port, pc_target_11_7_port, 
      pc_target_11_6_port, pc_target_11_5_port, pc_target_11_4_port, 
      pc_target_11_3_port, pc_target_11_2_port, pc_target_11_1_port, 
      pc_target_11_0_port, pc_target_14_31_port, pc_target_14_30_port, 
      pc_target_14_29_port, pc_target_14_28_port, pc_target_14_27_port, 
      pc_target_14_26_port, pc_target_14_25_port, pc_target_14_24_port, 
      pc_target_14_23_port, pc_target_14_22_port, pc_target_14_21_port, 
      pc_target_14_20_port, pc_target_14_19_port, pc_target_14_18_port, 
      pc_target_14_17_port, pc_target_14_16_port, pc_target_14_15_port, 
      pc_target_14_14_port, pc_target_14_13_port, pc_target_14_12_port, 
      pc_target_14_11_port, pc_target_14_10_port, pc_target_14_9_port, 
      pc_target_14_8_port, pc_target_14_7_port, pc_target_14_6_port, 
      pc_target_14_5_port, pc_target_14_4_port, pc_target_14_3_port, 
      pc_target_14_2_port, pc_target_14_1_port, pc_target_14_0_port, 
      pc_target_15_31_port, pc_target_15_30_port, pc_target_15_29_port, 
      pc_target_15_28_port, pc_target_15_27_port, pc_target_15_26_port, 
      pc_target_15_25_port, pc_target_15_24_port, pc_target_15_23_port, 
      pc_target_15_22_port, pc_target_15_21_port, pc_target_15_20_port, 
      pc_target_15_19_port, pc_target_15_18_port, pc_target_15_17_port, 
      pc_target_15_16_port, pc_target_15_15_port, pc_target_15_14_port, 
      pc_target_15_13_port, pc_target_15_12_port, pc_target_15_11_port, 
      pc_target_15_10_port, pc_target_15_9_port, pc_target_15_8_port, 
      pc_target_15_7_port, pc_target_15_6_port, pc_target_15_5_port, 
      pc_target_15_4_port, pc_target_15_3_port, pc_target_15_2_port, 
      pc_target_15_1_port, pc_target_15_0_port, pc_target_16_22_port, 
      pc_target_18_31_port, pc_target_18_30_port, pc_target_18_29_port, 
      pc_target_18_28_port, pc_target_18_27_port, pc_target_18_26_port, 
      pc_target_18_25_port, pc_target_18_24_port, pc_target_18_23_port, 
      pc_target_18_22_port, pc_target_18_21_port, pc_target_18_20_port, 
      pc_target_18_19_port, pc_target_18_18_port, pc_target_18_17_port, 
      pc_target_18_16_port, pc_target_18_15_port, pc_target_18_14_port, 
      pc_target_18_13_port, pc_target_18_12_port, pc_target_18_11_port, 
      pc_target_18_10_port, pc_target_18_9_port, pc_target_18_8_port, 
      pc_target_18_7_port, pc_target_18_6_port, pc_target_18_5_port, 
      pc_target_18_4_port, pc_target_18_3_port, pc_target_18_2_port, 
      pc_target_18_1_port, pc_target_18_0_port, pc_target_19_31_port, 
      pc_target_19_30_port, pc_target_19_29_port, pc_target_19_28_port, 
      pc_target_19_27_port, pc_target_19_26_port, pc_target_19_25_port, 
      pc_target_19_24_port, pc_target_19_23_port, pc_target_19_22_port, 
      pc_target_19_21_port, pc_target_19_20_port, pc_target_19_19_port, 
      pc_target_19_18_port, pc_target_19_17_port, pc_target_19_16_port, 
      pc_target_19_15_port, pc_target_19_14_port, pc_target_19_13_port, 
      pc_target_19_12_port, pc_target_19_11_port, pc_target_19_10_port, 
      pc_target_19_9_port, pc_target_19_8_port, pc_target_19_7_port, 
      pc_target_19_6_port, pc_target_19_5_port, pc_target_19_4_port, 
      pc_target_19_3_port, pc_target_19_2_port, pc_target_19_1_port, 
      pc_target_19_0_port, pc_target_20_31_port, pc_target_20_30_port, 
      pc_target_20_29_port, pc_target_20_28_port, pc_target_20_27_port, 
      pc_target_20_26_port, pc_target_20_25_port, pc_target_20_24_port, 
      pc_target_20_23_port, pc_target_20_22_port, pc_target_20_21_port, 
      pc_target_20_20_port, pc_target_20_19_port, pc_target_20_18_port, 
      pc_target_20_17_port, pc_target_20_16_port, pc_target_20_15_port, 
      pc_target_20_14_port, pc_target_20_13_port, pc_target_20_12_port, 
      pc_target_20_11_port, pc_target_20_10_port, pc_target_20_9_port, 
      pc_target_20_8_port, pc_target_20_7_port, pc_target_20_6_port, 
      pc_target_20_5_port, pc_target_20_4_port, pc_target_20_3_port, 
      pc_target_20_2_port, pc_target_20_1_port, pc_target_20_0_port, 
      pc_target_21_31_port, pc_target_21_30_port, pc_target_21_29_port, 
      pc_target_21_28_port, pc_target_21_27_port, pc_target_21_26_port, 
      pc_target_21_25_port, pc_target_21_24_port, pc_target_21_23_port, 
      pc_target_21_22_port, pc_target_21_21_port, pc_target_21_20_port, 
      pc_target_21_19_port, pc_target_21_18_port, pc_target_21_17_port, 
      pc_target_21_16_port, pc_target_21_15_port, pc_target_21_14_port, 
      pc_target_21_13_port, pc_target_21_12_port, pc_target_21_11_port, 
      pc_target_21_10_port, pc_target_21_9_port, pc_target_21_8_port, 
      pc_target_21_7_port, pc_target_21_6_port, pc_target_21_5_port, 
      pc_target_21_4_port, pc_target_21_3_port, pc_target_21_2_port, 
      pc_target_21_1_port, pc_target_21_0_port, pc_target_26_31_port, 
      pc_target_26_30_port, pc_target_26_29_port, pc_target_26_28_port, 
      pc_target_26_27_port, pc_target_26_26_port, pc_target_26_25_port, 
      pc_target_26_24_port, pc_target_26_23_port, pc_target_26_22_port, 
      pc_target_26_21_port, pc_target_26_20_port, pc_target_26_19_port, 
      pc_target_26_18_port, pc_target_26_17_port, pc_target_26_16_port, 
      pc_target_26_15_port, pc_target_26_14_port, pc_target_26_13_port, 
      pc_target_26_12_port, pc_target_26_11_port, pc_target_26_10_port, 
      pc_target_26_9_port, pc_target_26_8_port, pc_target_26_7_port, 
      pc_target_26_6_port, pc_target_26_5_port, pc_target_26_4_port, 
      pc_target_26_3_port, pc_target_26_2_port, pc_target_26_1_port, 
      pc_target_26_0_port, pc_target_27_31_port, pc_target_27_30_port, 
      pc_target_27_29_port, pc_target_27_28_port, pc_target_27_27_port, 
      pc_target_27_26_port, pc_target_27_25_port, pc_target_27_24_port, 
      pc_target_27_23_port, pc_target_27_22_port, pc_target_27_21_port, 
      pc_target_27_20_port, pc_target_27_19_port, pc_target_27_18_port, 
      pc_target_27_17_port, pc_target_27_16_port, pc_target_27_15_port, 
      pc_target_27_14_port, pc_target_27_13_port, pc_target_27_12_port, 
      pc_target_27_11_port, pc_target_27_10_port, pc_target_27_9_port, 
      pc_target_27_8_port, pc_target_27_7_port, pc_target_27_6_port, 
      pc_target_27_5_port, pc_target_27_4_port, pc_target_27_3_port, 
      pc_target_27_2_port, pc_target_27_1_port, pc_target_27_0_port, 
      pc_target_30_31_port, pc_target_30_30_port, pc_target_30_29_port, 
      pc_target_30_28_port, pc_target_30_27_port, pc_target_30_26_port, 
      pc_target_30_25_port, pc_target_30_24_port, pc_target_30_23_port, 
      pc_target_30_22_port, pc_target_30_21_port, pc_target_30_20_port, 
      pc_target_30_19_port, pc_target_30_18_port, pc_target_30_17_port, 
      pc_target_30_16_port, pc_target_30_15_port, pc_target_30_14_port, 
      pc_target_30_13_port, pc_target_30_12_port, pc_target_30_11_port, 
      pc_target_30_10_port, pc_target_30_9_port, pc_target_30_8_port, 
      pc_target_30_7_port, pc_target_30_6_port, pc_target_30_5_port, 
      pc_target_30_4_port, pc_target_30_3_port, pc_target_30_2_port, 
      pc_target_30_1_port, pc_target_30_0_port, pc_target_31_31_port, 
      pc_target_31_30_port, pc_target_31_29_port, pc_target_31_28_port, 
      pc_target_31_27_port, pc_target_31_26_port, pc_target_31_25_port, 
      pc_target_31_24_port, pc_target_31_23_port, pc_target_31_22_port, 
      pc_target_31_21_port, pc_target_31_20_port, pc_target_31_19_port, 
      pc_target_31_18_port, pc_target_31_17_port, pc_target_31_16_port, 
      pc_target_31_15_port, pc_target_31_14_port, pc_target_31_13_port, 
      pc_target_31_12_port, pc_target_31_11_port, pc_target_31_10_port, 
      pc_target_31_9_port, pc_target_31_8_port, pc_target_31_7_port, 
      pc_target_31_6_port, pc_target_31_5_port, pc_target_31_4_port, 
      pc_target_31_3_port, pc_target_31_2_port, pc_target_31_1_port, 
      pc_target_31_0_port, N96, N97, N98, N99, N100, N101, N102, N103, N104, 
      N105, N106, N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, 
      N117, N118, N119, N120, N121, N122, N123, N124, N125, N126, N127, 
      pc_lut_2_31_port, pc_lut_2_30_port, pc_lut_2_29_port, pc_lut_2_28_port, 
      pc_lut_2_27_port, pc_lut_2_26_port, pc_lut_2_25_port, pc_lut_2_24_port, 
      pc_lut_2_23_port, pc_lut_2_22_port, pc_lut_2_21_port, pc_lut_2_20_port, 
      pc_lut_2_19_port, pc_lut_2_18_port, pc_lut_2_17_port, pc_lut_2_16_port, 
      pc_lut_2_15_port, pc_lut_2_14_port, pc_lut_2_13_port, pc_lut_2_12_port, 
      pc_lut_2_11_port, pc_lut_2_10_port, pc_lut_2_9_port, pc_lut_2_8_port, 
      pc_lut_2_7_port, pc_lut_2_6_port, pc_lut_2_5_port, pc_lut_2_1_port, 
      pc_lut_3_31_port, pc_lut_3_30_port, pc_lut_3_29_port, pc_lut_3_28_port, 
      pc_lut_3_27_port, pc_lut_3_26_port, pc_lut_3_25_port, pc_lut_3_24_port, 
      pc_lut_3_23_port, pc_lut_3_22_port, pc_lut_3_21_port, pc_lut_3_20_port, 
      pc_lut_3_19_port, pc_lut_3_18_port, pc_lut_3_17_port, pc_lut_3_16_port, 
      pc_lut_3_15_port, pc_lut_3_14_port, pc_lut_3_13_port, pc_lut_3_12_port, 
      pc_lut_3_11_port, pc_lut_3_10_port, pc_lut_3_9_port, pc_lut_3_8_port, 
      pc_lut_3_7_port, pc_lut_3_6_port, pc_lut_3_5_port, pc_lut_3_1_port, 
      pc_lut_3_0_port, pc_lut_6_31_port, pc_lut_6_30_port, pc_lut_6_29_port, 
      pc_lut_6_28_port, pc_lut_6_27_port, pc_lut_6_26_port, pc_lut_6_25_port, 
      pc_lut_6_24_port, pc_lut_6_23_port, pc_lut_6_22_port, pc_lut_6_21_port, 
      pc_lut_6_20_port, pc_lut_6_19_port, pc_lut_6_18_port, pc_lut_6_17_port, 
      pc_lut_6_16_port, pc_lut_6_15_port, pc_lut_6_14_port, pc_lut_6_13_port, 
      pc_lut_6_12_port, pc_lut_6_11_port, pc_lut_6_10_port, pc_lut_6_9_port, 
      pc_lut_6_8_port, pc_lut_6_7_port, pc_lut_6_6_port, pc_lut_6_5_port, 
      pc_lut_6_2_port, pc_lut_6_1_port, pc_lut_7_31_port, pc_lut_7_30_port, 
      pc_lut_7_29_port, pc_lut_7_28_port, pc_lut_7_27_port, pc_lut_7_26_port, 
      pc_lut_7_25_port, pc_lut_7_24_port, pc_lut_7_23_port, pc_lut_7_22_port, 
      pc_lut_7_21_port, pc_lut_7_20_port, pc_lut_7_19_port, pc_lut_7_18_port, 
      pc_lut_7_17_port, pc_lut_7_16_port, pc_lut_7_15_port, pc_lut_7_14_port, 
      pc_lut_7_13_port, pc_lut_7_12_port, pc_lut_7_11_port, pc_lut_7_10_port, 
      pc_lut_7_9_port, pc_lut_7_8_port, pc_lut_7_7_port, pc_lut_7_6_port, 
      pc_lut_7_5_port, pc_lut_7_2_port, pc_lut_7_1_port, pc_lut_7_0_port, 
      pc_lut_10_31_port, pc_lut_10_30_port, pc_lut_10_29_port, 
      pc_lut_10_28_port, pc_lut_10_27_port, pc_lut_10_26_port, 
      pc_lut_10_25_port, pc_lut_10_24_port, pc_lut_10_23_port, 
      pc_lut_10_22_port, pc_lut_10_21_port, pc_lut_10_20_port, 
      pc_lut_10_19_port, pc_lut_10_18_port, pc_lut_10_17_port, 
      pc_lut_10_16_port, pc_lut_10_15_port, pc_lut_10_14_port, 
      pc_lut_10_13_port, pc_lut_10_12_port, pc_lut_10_11_port, 
      pc_lut_10_10_port, pc_lut_10_9_port, pc_lut_10_8_port, pc_lut_10_7_port, 
      pc_lut_10_6_port, pc_lut_10_5_port, pc_lut_10_3_port, pc_lut_10_1_port, 
      pc_lut_11_31_port, pc_lut_11_30_port, pc_lut_11_29_port, 
      pc_lut_11_28_port, pc_lut_11_27_port, pc_lut_11_26_port, 
      pc_lut_11_25_port, pc_lut_11_24_port, pc_lut_11_23_port, 
      pc_lut_11_22_port, pc_lut_11_21_port, pc_lut_11_20_port, 
      pc_lut_11_19_port, pc_lut_11_18_port, pc_lut_11_17_port, 
      pc_lut_11_16_port, pc_lut_11_15_port, pc_lut_11_14_port, 
      pc_lut_11_13_port, pc_lut_11_12_port, pc_lut_11_11_port, 
      pc_lut_11_10_port, pc_lut_11_9_port, pc_lut_11_8_port, pc_lut_11_7_port, 
      pc_lut_11_6_port, pc_lut_11_5_port, pc_lut_11_3_port, pc_lut_11_1_port, 
      pc_lut_11_0_port, pc_lut_14_31_port, pc_lut_14_30_port, pc_lut_14_29_port
      , pc_lut_14_28_port, pc_lut_14_27_port, pc_lut_14_26_port, 
      pc_lut_14_25_port, pc_lut_14_24_port, pc_lut_14_23_port, 
      pc_lut_14_22_port, pc_lut_14_21_port, pc_lut_14_20_port, 
      pc_lut_14_19_port, pc_lut_14_18_port, pc_lut_14_17_port, 
      pc_lut_14_16_port, pc_lut_14_15_port, pc_lut_14_14_port, 
      pc_lut_14_13_port, pc_lut_14_12_port, pc_lut_14_11_port, 
      pc_lut_14_10_port, pc_lut_14_9_port, pc_lut_14_8_port, pc_lut_14_7_port, 
      pc_lut_14_6_port, pc_lut_14_5_port, pc_lut_14_3_port, pc_lut_14_2_port, 
      pc_lut_14_1_port, pc_lut_15_31_port, pc_lut_15_30_port, pc_lut_15_29_port
      , pc_lut_15_28_port, pc_lut_15_27_port, pc_lut_15_26_port, 
      pc_lut_15_25_port, pc_lut_15_24_port, pc_lut_15_23_port, 
      pc_lut_15_22_port, pc_lut_15_21_port, pc_lut_15_20_port, 
      pc_lut_15_19_port, pc_lut_15_18_port, pc_lut_15_17_port, 
      pc_lut_15_16_port, pc_lut_15_15_port, pc_lut_15_14_port, 
      pc_lut_15_13_port, pc_lut_15_12_port, pc_lut_15_11_port, 
      pc_lut_15_10_port, pc_lut_15_9_port, pc_lut_15_8_port, pc_lut_15_7_port, 
      pc_lut_15_6_port, pc_lut_15_5_port, pc_lut_15_3_port, pc_lut_15_2_port, 
      pc_lut_15_1_port, pc_lut_15_0_port, pc_lut_18_31_port, pc_lut_18_30_port,
      pc_lut_18_29_port, pc_lut_18_28_port, pc_lut_18_27_port, 
      pc_lut_18_26_port, pc_lut_18_25_port, pc_lut_18_24_port, 
      pc_lut_18_23_port, pc_lut_18_22_port, pc_lut_18_21_port, 
      pc_lut_18_20_port, pc_lut_18_19_port, pc_lut_18_18_port, 
      pc_lut_18_17_port, pc_lut_18_16_port, pc_lut_18_15_port, 
      pc_lut_18_14_port, pc_lut_18_13_port, pc_lut_18_12_port, 
      pc_lut_18_11_port, pc_lut_18_10_port, pc_lut_18_9_port, pc_lut_18_8_port,
      pc_lut_18_7_port, pc_lut_18_6_port, pc_lut_18_5_port, pc_lut_18_4_port, 
      pc_lut_18_1_port, pc_lut_19_31_port, pc_lut_19_30_port, pc_lut_19_29_port
      , pc_lut_19_28_port, pc_lut_19_27_port, pc_lut_19_26_port, 
      pc_lut_19_25_port, pc_lut_19_24_port, pc_lut_19_23_port, 
      pc_lut_19_22_port, pc_lut_19_21_port, pc_lut_19_20_port, 
      pc_lut_19_19_port, pc_lut_19_18_port, pc_lut_19_17_port, 
      pc_lut_19_16_port, pc_lut_19_15_port, pc_lut_19_14_port, 
      pc_lut_19_13_port, pc_lut_19_12_port, pc_lut_19_11_port, 
      pc_lut_19_10_port, pc_lut_19_9_port, pc_lut_19_8_port, pc_lut_19_7_port, 
      pc_lut_19_6_port, pc_lut_19_5_port, pc_lut_19_4_port, pc_lut_19_1_port, 
      pc_lut_19_0_port, pc_lut_20_31_port, pc_lut_20_30_port, pc_lut_20_29_port
      , pc_lut_20_28_port, pc_lut_20_27_port, pc_lut_20_26_port, 
      pc_lut_20_25_port, pc_lut_20_24_port, pc_lut_20_23_port, 
      pc_lut_20_22_port, pc_lut_20_21_port, pc_lut_20_20_port, 
      pc_lut_20_19_port, pc_lut_20_18_port, pc_lut_20_17_port, 
      pc_lut_20_16_port, pc_lut_20_15_port, pc_lut_20_14_port, 
      pc_lut_20_13_port, pc_lut_20_12_port, pc_lut_20_11_port, 
      pc_lut_20_10_port, pc_lut_20_9_port, pc_lut_20_8_port, pc_lut_20_7_port, 
      pc_lut_20_6_port, pc_lut_20_5_port, pc_lut_20_4_port, pc_lut_20_2_port, 
      pc_lut_21_31_port, pc_lut_21_30_port, pc_lut_21_29_port, 
      pc_lut_21_28_port, pc_lut_21_27_port, pc_lut_21_26_port, 
      pc_lut_21_25_port, pc_lut_21_24_port, pc_lut_21_23_port, 
      pc_lut_21_22_port, pc_lut_21_21_port, pc_lut_21_20_port, 
      pc_lut_21_19_port, pc_lut_21_18_port, pc_lut_21_17_port, 
      pc_lut_21_16_port, pc_lut_21_15_port, pc_lut_21_14_port, 
      pc_lut_21_13_port, pc_lut_21_12_port, pc_lut_21_11_port, 
      pc_lut_21_10_port, pc_lut_21_9_port, pc_lut_21_8_port, pc_lut_21_7_port, 
      pc_lut_21_6_port, pc_lut_21_5_port, pc_lut_21_4_port, pc_lut_21_2_port, 
      pc_lut_21_0_port, pc_lut_26_31_port, pc_lut_26_30_port, pc_lut_26_29_port
      , pc_lut_26_28_port, pc_lut_26_27_port, pc_lut_26_26_port, 
      pc_lut_26_25_port, pc_lut_26_24_port, pc_lut_26_23_port, 
      pc_lut_26_22_port, pc_lut_26_21_port, pc_lut_26_20_port, 
      pc_lut_26_19_port, pc_lut_26_18_port, pc_lut_26_17_port, 
      pc_lut_26_16_port, pc_lut_26_15_port, pc_lut_26_14_port, 
      pc_lut_26_13_port, pc_lut_26_12_port, pc_lut_26_11_port, 
      pc_lut_26_10_port, pc_lut_26_9_port, pc_lut_26_8_port, pc_lut_26_7_port, 
      pc_lut_26_6_port, pc_lut_26_5_port, pc_lut_26_4_port, pc_lut_26_3_port, 
      pc_lut_26_1_port, pc_lut_27_31_port, pc_lut_27_30_port, pc_lut_27_29_port
      , pc_lut_27_28_port, pc_lut_27_27_port, pc_lut_27_26_port, 
      pc_lut_27_25_port, pc_lut_27_24_port, pc_lut_27_23_port, 
      pc_lut_27_22_port, pc_lut_27_21_port, pc_lut_27_20_port, 
      pc_lut_27_19_port, pc_lut_27_18_port, pc_lut_27_17_port, 
      pc_lut_27_16_port, pc_lut_27_15_port, pc_lut_27_14_port, 
      pc_lut_27_13_port, pc_lut_27_12_port, pc_lut_27_11_port, 
      pc_lut_27_10_port, pc_lut_27_9_port, pc_lut_27_8_port, pc_lut_27_7_port, 
      pc_lut_27_6_port, pc_lut_27_5_port, pc_lut_27_4_port, pc_lut_27_3_port, 
      pc_lut_27_1_port, pc_lut_27_0_port, pc_lut_30_31_port, pc_lut_30_30_port,
      pc_lut_30_29_port, pc_lut_30_28_port, pc_lut_30_27_port, 
      pc_lut_30_26_port, pc_lut_30_25_port, pc_lut_30_24_port, 
      pc_lut_30_23_port, pc_lut_30_22_port, pc_lut_30_21_port, 
      pc_lut_30_20_port, pc_lut_30_19_port, pc_lut_30_18_port, 
      pc_lut_30_17_port, pc_lut_30_16_port, pc_lut_30_15_port, 
      pc_lut_30_14_port, pc_lut_30_13_port, pc_lut_30_12_port, 
      pc_lut_30_11_port, pc_lut_30_10_port, pc_lut_30_9_port, pc_lut_30_8_port,
      pc_lut_30_7_port, pc_lut_30_6_port, pc_lut_30_5_port, pc_lut_30_4_port, 
      pc_lut_30_3_port, pc_lut_30_2_port, pc_lut_30_1_port, pc_lut_31_31_port, 
      pc_lut_31_30_port, pc_lut_31_29_port, pc_lut_31_28_port, 
      pc_lut_31_27_port, pc_lut_31_26_port, pc_lut_31_25_port, 
      pc_lut_31_24_port, pc_lut_31_23_port, pc_lut_31_22_port, 
      pc_lut_31_21_port, pc_lut_31_20_port, pc_lut_31_19_port, 
      pc_lut_31_18_port, pc_lut_31_17_port, pc_lut_31_16_port, 
      pc_lut_31_15_port, pc_lut_31_14_port, pc_lut_31_13_port, 
      pc_lut_31_12_port, pc_lut_31_11_port, pc_lut_31_10_port, pc_lut_31_9_port
      , pc_lut_31_8_port, pc_lut_31_7_port, pc_lut_31_6_port, pc_lut_31_5_port,
      pc_lut_31_4_port, pc_lut_31_3_port, pc_lut_31_2_port, pc_lut_31_1_port, 
      pc_lut_31_0_port, N188, N189, N190, N191, N192, N193, N194, N195, N196, 
      N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, 
      N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, 
      n1, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33
      , n34, n35, n36, n37, n38, n39, n40, n42, n43, n44, n45, n46, n47, n48, 
      n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63
      , n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
      n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92
      , n93, n94, n95, n96_port, n97_port, n98_port, n99_port, n100_port, 
      n101_port, n102_port, n103_port, n104_port, n105_port, n106_port, 
      n107_port, n108_port, n109_port, n110_port, n111_port, n112_port, 
      n113_port, n114_port, n115_port, n116_port, n117_port, n118_port, 
      n119_port, n120_port, n121_port, n122_port, n123_port, n124_port, 
      n125_port, n126_port, n127_port, n128, n129, n130, n131, n132, n133, n134
      , n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n181, n182, n183, 
      n184, n185, n186, n187, n188_port, n189_port, n190_port, n191_port, 
      n192_port, n193_port, n194_port, n195_port, n196_port, n197_port, 
      n198_port, n199_port, n200_port, n201_port, n202_port, n203_port, 
      n204_port, n205_port, n206_port, n207_port, n208_port, n209_port, 
      n210_port, n211_port, n212_port, n213_port, n214_port, n215_port, 
      n216_port, n217_port, n218_port, n219_port, n220_port, n221, n222, n223, 
      n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, 
      n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
      n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n284, 
      n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, 
      n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, 
      n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, 
      n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, 
      n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, 
      n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, 
      n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, 
      n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, 
      n381, n382, n383, n384, n385, n386, n388, n389, n390, n391, n392, n393, 
      n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, 
      n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, 
      n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, 
      n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, 
      n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, 
      n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, 
      n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, 
      n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, 
      n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, 
      n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, 
      n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n526, 
      n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, 
      n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, 
      n551, n552, n553, n554, n555, n556, n557, n559, n560, n561, n562, n563, 
      n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, 
      n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, 
      n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, 
      n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, 
      n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, 
      n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, 
      n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, 
      n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, 
      n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, 
      n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, 
      n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, 
      n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, 
      n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, 
      n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, 
      n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, 
      n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, 
      n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, 
      n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, 
      n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, 
      n793, n794, n795, n796, n797, n798, n799, n800, n801, n803, n804, n805, 
      n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, 
      n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, 
      n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, 
      n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, 
      n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, 
      n866, n867, n868, n869, n870, n872, n873, n874, n875, n876, n877, n878, 
      n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, 
      n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, 
      n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, 
      n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, 
      n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, 
      n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, 
      n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, 
      n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n974, n975, 
      n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, 
      n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, 
      n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, 
      n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, 
      n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, 
      n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, 
      n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, 
      n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, 
      n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, 
      n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, 
      n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, 
      n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, 
      n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, 
      n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, 
      n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, 
      n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, 
      n1140, n1141, n1142, n1143, n1144, n1146, n1147, n1148, n1149, n1150, 
      n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, 
      n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, 
      n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, 
      n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, 
      n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, 
      n1201, n1202, n1203, n1204, n1205, n1206, n1208, n1209, n1210, n1211, 
      n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, 
      n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, 
      n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1241, n1242, 
      n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, 
      n1253, n1254, n1255, n1257, n1258, n1260, n1261, n1262, n1263, n1264, 
      n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, 
      n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, 
      n1286, n1287, n1288, n1289, n1290, n1291, n1294, n1295, n1296, n1297, 
      n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, 
      n1308, n1309, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, 
      n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, 
      n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, 
      n1339, n1340, n1341, n1342, n1343, n1345, n1346, n1347, n1348, n1349, 
      n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, 
      n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, 
      n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, 
      n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, 
      n1390, n1391, n1393, n1395, n1396, n1397, n1398, n1399, n1400, n1401, 
      n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, 
      n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, 
      n1422, n1423, n1424, n1425, n1429, n1430, n1431, n1432, n1433, n1434, 
      n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, 
      n1445, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, 
      n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1464, n1465, n1466, 
      n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, 
      n1477, n1478, n1479, n1480, n1482, n1483, n1484, n1485, n1486, n1487, 
      n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1497, n1499, 
      n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, 
      n1510, n1511, n1512, n1514, n1515, n1516, n1517, n1518, n1519, n1520, 
      n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, 
      n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, 
      n1541, n1542, n1543, n1544, n1546, n1547, n1548, n1549, n1550, n1551, 
      n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, 
      n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, 
      n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, 
      n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, 
      n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, 
      n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1612, 
      n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, 
      n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, 
      n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, 
      n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, 
      n1653, n1654, n1655, n1657, n1660, n1661, n1662, n1663, n1664, n1665, 
      n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, 
      n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, 
      n1686, n1687, n1688, n1689, n1694, n1695, n1696, n1697, n1698, n1699, 
      n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1710, 
      n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, 
      n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, 
      n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, 
      n1741, n1742, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, 
      n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, 
      n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, 
      n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, 
      n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1791, n1792, 
      n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, 
      n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, 
      n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, 
      n1825, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, 
      n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, 
      n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, 
      n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, 
      n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, 
      n1877, n1878, n1879, n1880, n1882, n1883, n1884, n1885, n1886, n1887, 
      n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, 
      n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, 
      n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, 
      n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1927, n1929, n1930, 
      n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, 
      n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, 
      n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1963, n1964, 
      n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, 
      n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, 
      n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, 
      n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, 
      n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2014, n2015, 
      n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, 
      n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, 
      n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, 
      n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, 
      n2056, n2058, n2059, n2062, n2063, n2064, n2065, n2066, n2067, n2068, 
      n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, 
      n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, 
      n2089, n2090, n2092, n2096, n2097, n2098, n2099, n2100, n2101, n2102, 
      n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2113, 
      n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, 
      n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, 
      n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, 
      n2144, n2145, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, 
      n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, 
      n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, 
      n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, 
      n2185, n2186, n2187, n2188, n2191, n2194, n2195, n2196, n2197, n2198, 
      n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, 
      n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, 
      n2219, n2220, n2221, n2222, n2228, n2229, n2230, n2231, n2232, n2233, 
      n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, 
      n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, 
      n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, 
      n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, 
      n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, 
      n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, 
      n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, 
      n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, 
      n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, 
      n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, 
      n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, 
      n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, 
      n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, 
      n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2374, 
      n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, 
      n2386, n2389, n2391, n2392, n2394, n2397, n2399, n2400, n2401, n2404, 
      n2405, n2406, n2407, n2412, n2413, n2414, n2415, n2419, n2420, n2421, 
      n2422, n2423, n2424, n2425, n2426, n2427, n2436, n2437, n2438, n2439, 
      n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, 
      n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, 
      n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, 
      n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, 
      n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, 
      n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, 
      n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, 
      n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, 
      n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, 
      n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, 
      n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, 
      n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, 
      n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, 
      n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, 
      n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, 
      n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, 
      n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, 
      n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, 
      n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, 
      n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, 
      n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, 
      n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, 
      n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, 
      n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, 
      n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, 
      n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, 
      n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, 
      n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, 
      n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, 
      n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, 
      n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, 
      n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, 
      n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, 
      n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, 
      n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, 
      n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, 
      n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, 
      n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, 
      n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, 
      n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, 
      n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, 
      n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, 
      n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, 
      n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, 
      n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, 
      n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, 
      n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, 
      n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, 
      n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, 
      n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, 
      n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, 
      n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, 
      n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, 
      n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, 
      n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, 
      n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, 
      n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, 
      n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, 
      n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, 
      n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, 
      n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, 
      n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, 
      n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, 
      n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, 
      n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, 
      n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, 
      n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, 
      n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, 
      n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, 
      n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, 
      n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, 
      n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, 
      n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, 
      n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, 
      n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, 
      n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, 
      n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, 
      n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, 
      n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, 
      n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, 
      n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, 
      n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, 
      n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, 
      n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, 
      n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, 
      n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, 
      n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, 
      n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, 
      n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, 
      n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, 
      n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, 
      n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, 
      n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, 
      n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, 
      n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, 
      n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, 
      n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, 
      n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, 
      n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, 
      n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, 
      n3440, n3441, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, 
      n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, 
      n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, 
      n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, 
      n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, 
      n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, 
      n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, 
      n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, 
      n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, 
      n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, 
      n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, 
      n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, 
      n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, 
      n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, 
      n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, 
      n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, 
      n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, 
      n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, 
      n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, 
      n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, 
      n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, 
      n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, 
      n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, 
      n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, 
      n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, 
      n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, 
      n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, 
      n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, 
      n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, 
      n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, 
      n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, 
      n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, 
      n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, 
      n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, 
      n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, 
      n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, 
      n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, 
      n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, 
      n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, 
      n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, 
      n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, 
      n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, 
      n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, 
      n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, 
      n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, 
      n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, 
      n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, 
      n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, 
      n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, 
      n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, 
      n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, 
      n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, 
      n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, 
      n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, 
      n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, 
      n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, 
      n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, 
      n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, 
      n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, 
      n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, 
      n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, 
      n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, 
      n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, 
      n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, 
      n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, 
      n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, 
      n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, 
      n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, 
      n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, 
      n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, 
      n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, 
      n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, 
      n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, 
      n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, 
      n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, 
      n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, 
      n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, 
      n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, 
      n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, 
      n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, 
      n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, 
      n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, 
      n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, 
      n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, 
      n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, 
      n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, 
      n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, 
      n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, 
      n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, 
      n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, 
      n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, 
      n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, 
      n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, 
      n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, 
      n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, 
      n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, 
      n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, 
      n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, 
      n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, 
      n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, 
      n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, 
      n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, 
      n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, 
      n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, 
      n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, 
      n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, 
      n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, 
      n6558, n6559, n6560, n6562, n6563, n6564, n6565, n6566, n6567, n6568, 
      n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, 
      n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, 
      n6589, n6590, n6591, n6592, n6593, n6595, n6596, n6597, n6598, n6599, 
      n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, 
      n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, 
      n6620, n6621, n6622, n6623, n6624, n6627, n6628, n6629, n6630, n6631, 
      n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, 
      n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, 
      n6652, n6653, n6654, n6655, n6657, n6658, n6659, n6660, n6661, n6662, 
      n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, 
      n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, 
      n6683, n6684, n6685, n6686, n6687, n6690, n6691, n6692, n6693, n6694, 
      n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, 
      n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, 
      n6715, n6716, n6717, n6718, n6719, n6721, n6723, n6724, n6725, n6726, 
      n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, 
      n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, 
      n6747, n6748, n6749, n6750, n6751, n6755, n6756, n6757, n6758, n6759, 
      n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, 
      n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, 
      n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6788, n6789, n6790, 
      n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, 
      n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, 
      n6811, n6812, n6813, n6814, n6815, n6816, n6818, n6820, n6821, n6822, 
      n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, 
      n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, 
      n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6852, n6853, n6854, 
      n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, 
      n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, 
      n6875, n6876, n6877, n6878, n6879, n6880, n6884, n6885, n6886, n6887, 
      n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, 
      n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, 
      n6908, n6909, n6910, n6911, n6913, n6914, n6916, n6917, n6918, n6919, 
      n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, 
      n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, 
      n6940, n6941, n6942, n6943, n6946, n6948, n6949, n6950, n6951, n6952, 
      n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, 
      n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, 
      n6973, n6974, n6975, n6977, n6980, n6981, n6982, n6983, n6984, n6985, 
      n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, 
      n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, 
      n7006, n7007, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, 
      n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, 
      n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7040, 
      n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, 
      n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, 
      n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, 
      n7072, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, 
      n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, 
      n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, 
      n7104, n7105, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, 
      n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, 
      n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, 
      n7136, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, 
      n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, 
      n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7169, 
      n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, 
      n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, 
      n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7202, 
      n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, 
      n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, 
      n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7233, n7235, 
      n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, 
      n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, 
      n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7267, n7268, n7269, 
      n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, 
      n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, 
      n7290, n7291, n7292, n7293, n7294, n7296, n7297, n7298, n7300, n7301, 
      n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, 
      n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, 
      n7322, n7323, n7324, n7325, n7326, n7328, n7330, n7332, n7333, n7334, 
      n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, 
      n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, 
      n7355, n7356, n7357, n7358, n7360, n7361, n7364, n7365, n7366, n7367, 
      n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, 
      n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, 
      n7388, n7389, n7390, n7392, n7396, n7397, n7398, n7399, n7400, n7401, 
      n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, 
      n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, 
      n7422, n7425, n7426, n7428, n7429, n7430, n7431, n7432, n7433, n7434, 
      n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, 
      n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, 
      n7458, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, 
      n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, 
      n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7489, n7492, 
      n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, 
      n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, 
      n7513, n7514, n7515, n7516, n7517, n7518, n7524, n7525, n7526, n7527, 
      n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n2,
      n3, n283, n525, n558, n768, n802, n871, n973, n1240, n1256, n1259, n1275,
      n1292, n1293, n1344, n1392, n1394, n1426, n1427, n1428, n1446, n1463, 
      n1481, n1496, n1498, n1611, n1656, n1658, n1659, n1690, n1691, n1692, 
      n1693, n1709, n1743, n1790, n1793, n1824, n1826, n1827, n1881, n1925, 
      n1926, n1928, n1959, n1960, n1961, n1962, n2013, n2057, n2060, n2061, 
      n2091, n2093, n2094, n2095, n2112, n2146, n2189, n2190, n2192, n2193, 
      n2223, n2224, n2225, n2226, n2227, n2373, n2385, n2387, n2388, n2390, 
      n2393, n2395, n2396, n2398, n2402, n2403, n2408, n2409, n2410, n2411, 
      n2416, n2417, n2418, n2428, n2429, n2430, n2431, n2432, n2433, n2434, 
      n2435, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, 
      n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, 
      n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, 
      n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, 
      n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, 
      n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, 
      n3501, n3502, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, 
      n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, 
      n3536, n3537, n3538, net113295, net113296, net113297, net113298, 
      net113299, net113300, net113301, net113302, net113303, net113304, 
      net113305, net113306, net113307, net113308, net113309, net113310, 
      net113311, net113312, net113313, net113314, net113315, net113316, 
      net113317, net113318, net113319, net113320, net113321, net113322, 
      net113323, net113324, net113325, net113326, net113327, net113328, 
      net113329, net113330, net113331, net113332, net113333, net113334, 
      net113335, net113336, net113337, net113338, net113339, net113340, 
      net113341, net113342, net113343, net113344, net113345, net113346, 
      net113347, net113348, net113349, net113350, net113351, net113352, 
      net113353, net113354, net113355, net113356, net113357, net113358, 
      net113359, net113360, net113361, net113362, net113363, net113364, 
      net113365, net113366, net113367, net113368, net113369, net113372, 
      net113375, net113377, net113378, net113379, net113380, net113381, 
      net113382, net113383, net113384, net113385, net113386, net113387, 
      net113388, net113389, net113390, net113391, net113392, net113393, 
      net113394, net113395, net113396, net113397, net113398, net113399, 
      net113400, net113403, net113406, net113408, net113409, net113410, 
      net113411, net113412, net113413, net113414, net113415, net113416, 
      net113417, net113418, net113419, net113420, net113421, net113422, 
      net113423, net113424, net113425, net113426, net113427, net113428, 
      net113429, net113430, net113431, net113432, net113433, net113434, 
      net113435, net113436, net113437, net113438, net113439, net113440, 
      net113441, net113442, net113443, net113444, net113445, net113446, 
      net113447, net113448, net113449, net113450, net113451, net113452, 
      net113453, net113454, net113455, net113456, net113457, net113458, 
      net113459, net113460, net113461, net113462, net113463, net113464, 
      net113465, net113466, net113467, net113468, net113469, net113470, 
      net113471, net113472, net113473, net113474, net113475, net113476, 
      net113477, net113478, net113479, net113480, net113481, net113482, 
      net113483, net113484, net113485, net113486, net113487, net113488, 
      net113489, net113490, net113491, net113492, net113493, net113494, 
      net113495, net113496, net113497, net113498, net113499, net113500, 
      net113501, net113502, net113503, net113504, net113505, net113506, 
      net113507, net113508, net113509, net113510, net113511, net113512, 
      net113513, net113514, net113515, net113516, net113517, net113518, 
      net113519, net113520, net113521, net113522, net113523, net113524, 
      net113525, net113526, net113528, net113531, net113532, net113533, 
      net113534, net113535, net113536, net113537, net113538, net113539, 
      net113540, net113541, net113542, net113543, net113544, net113545, 
      net113546, net113547, net113548, net113549, net113550, net113551, 
      net113552, net113553, net113554, net113555, net113558, net113561, 
      net113563, net113564, net113565, net113566, net113567, net113568, 
      net113569, net113570, net113571, net113572, net113573, net113574, 
      net113575, net113576, net113577, net113578, net113579, net113580, 
      net113581, net113582, net113583, net113584, net113585, net113586, 
      net113589, net113592, net113594, net113595, net113596, net113597, 
      net113598, net113599, net113600, net113601, net113602, net113603, 
      net113604, net113605, net113606, net113607, net113608, net113609, 
      net113610, net113611, net113612, net113613, net113614, net113615, 
      net113616, net113617, net113618, net113619, net113620, net113621, 
      net113622, net113623, net113624, net113625, net113626, net113627, 
      net113628, net113629, net113630, net113631, net113632, net113633, 
      net113634, net113635, net113636, net113637, net113638, net113639, 
      net113640, net113641, net113642, net113643, net113644, net113645, 
      net113646, net113647, net113648, net113649, net113650, net113651, 
      net113652, net113653, net113654, net113655, net113656, net113657, 
      net113658, net113659, net113660, net113661, net113662, net113663, 
      net113664, net113665, net113666, net113667, net113668, net113669, 
      net113670, net113671, net113672, net113673, net113674, net113675, 
      net113676, net113677, net113678, net113679, net113680, net113681, 
      net113682, net113683, net113684, net113685, net113686, net113687, 
      net113688, net113689, net113690, net113691, net113692, net113693, 
      net113694, net113695, net113696, net113697, net113698, net113699, 
      net113700, net113701, net113702, net113703, net113704, net113705, 
      net113706, net113707, net113708, net113709, net113710, net113711, 
      net113712, net113713, net113714, net113715, net113716, net113717, 
      net113718, net113719, net113720, net113721, net113722, net113723, 
      net113724, net113725, net113726, net113727, net113728, net113729, 
      net113730, net113731, net113732, net113733, net113734, net113735, 
      net113736, net113737, net113738, net113739, net113741, net113744, 
      net113745, net113746, net113747, net113748, net113749, net113750, 
      net113751, net113752, net113753, net113754, net113755, net113756, 
      net113757, net113758, net113759, net113760, net113762, net113763, 
      net113764, net113765, net113766, net113767, net113768, net113769, 
      net113770, net113771, net113772, net113773, net113774, net113775, 
      net113776, net113777, net113778, net113779, net113780, net113781, 
      net113782, net113783, net113784, net113785, net113786, net113787, 
      net113788, net113789, net113790, net113791, net113792, net113793, 
      net113794, net113795, net113796, net113797, net113798, net113799, 
      net113800, net113801, net113802, net113803, net113804, net113805, 
      net113806, net113807, net113808, net113809, net113810, net113811, 
      net113812, net113813, net113814, net113815, net113816, net113817, 
      net113818, net113819, net113820, net113821, net113822, net113823, 
      net113824, net113825, net113826, net113827, net113828, net113829, 
      net113830, net113831, net113832, net113833, net113834, net113835, 
      net113836, net113837, net113838, net113839, net113840, net113841, 
      net113842, net113843, net113844, net113845, net113846, net113847, 
      net113848, net113849, net113850, net113851, net113852, net113853, 
      net113856, net113859, net113861, net113862, net113863, net113864, 
      net113865, net113866, net113867, net113868, net113869, net113870, 
      net113871, net113872, net113873, net113874, net113875, net113876, 
      net113877, net113878, net113879, net113880, net113881, net113882, 
      net113883, net113884, net113887, net113890, net113892, net113893, 
      net113894, net113895, net113896, net113897, net113898, net113899, 
      net113900, net113901, net113902, net113903, net113904, net113905, 
      net113906, net113907, net113908, net113909, net113910, net113911, 
      net113912, net113913, net113914, net113915, net113916, net113917, 
      net113918, net113919, net113920, net113921, net113922, net113923, 
      net113924, net113925, net113926, net113927, net113928, net113929, 
      net113930, net113931, net113932, net113933, net113934, net113935, 
      net113936, net113937, net113938, net113939, net113940, net113941, 
      net113942, net113943, net113944, net113945, net113946, net113947, 
      net113948, net113949, net113950, net113951, net113952, net113953, 
      net113954, net113955, net113956, net113957, net113958, net113959, 
      net113960, net113961, net113962, net113963, net113964, net113965, 
      net113966, net113967, net113968, net113969, net113970, net113971, 
      net113972, net113973, net113974, net113975, net113977, net113980, 
      net113981, net113982, net113983, net113984, net113985, net113986, 
      net113987, net113988, net113989, net113990, net113991, net113992, 
      net113993, net113994, net113995, net113996, net113997, net113998, 
      net113999, net114000, net114001, net114002, net114003, net114004, 
      net114005, net114006, net114007, net114008, net114009, net114010, 
      net114011, net114012, net114013, net114014, net114015, net114016, 
      net114017, net114018, net114019, net114020, net114021, net114022, 
      net114023, net114024, net114037, net114038, net114039, net114040, 
      net114041, net114042, net114043, net114057, net114058, net114059, 
      net114060, net114061, net114062, net114063, net114064, net114065, 
      net114066, net114067, net114068, net114069, net114070, net114071, 
      net114072, net114073, net114074, net114075, net114076, net114077, 
      net114078, net114079, net114080, net114081, net114082, net114083, 
      net114084, net114085, net114086, net114087, net114088, net114089, 
      net114090, net114091, net114092, net114093, net114094, net114095, 
      net114096, net114097, net114098, net114100, net114103, net114104, 
      net114105, net114106, net114107, net114108, net114109, net114110, 
      net114111, net114112, net114113, net114114, net114115, net114116, 
      net114117, net114118, net114119, net114120, net114121, net114122, 
      net114123, net114124, net114125, net114126, net114127, net114128, 
      net114129, net114130, net114131, net114132, net114133, net114134, 
      net114135, net114136, net114137, net114138, net114139, net114140, 
      net114141, net114142, net114143, net114144, net114145, net114146, 
      net114147, net114148, net114149, net114152, net114155, net114157, 
      net114158, net114159, net114160, net114161, net114162, net114163, 
      net114164, net114165, net114166, net114167, net114168, net114169, 
      net114170, net114171, net114172, net114173, net114174, net114175, 
      net114176, net114177, net114178, net114179, net114180, net114183, 
      net114186, net114188, net114189, net114190, net114191, net114192, 
      net114193, net114194, net114195, net114196, net114197, net114198, 
      net114199, net114200, net114206, net114207, net114208, net114209, 
      net114295, net114296, net114297, net114298, net114299, net114300, 
      net114301, net114302, net114303, net114304, net114305, net114306, 
      net114307, net114308, net114309, net114310, net114311, net114312, 
      net114313, net114314, net114315, net114316, net114317, net114318, 
      net114319, net114320, net114321, net114322, net114323, net114324, 
      net114325, net114326, net114327, net114328, net114329, net114330, 
      net114331, net114332, net114333, net114334, net114335, net114336, 
      net114337, net114338, net114339, net114340, net114341, net114342, 
      net114343, net114344, net114345, net114346, net114347, net114348, 
      net114349, net114350, net114351, net114352, net114353, net114354, 
      net114355, net114356, net114357, net114358, net114359, net114360, 
      net114361, net114362, net114363, net114364, net114365, net114366, 
      net114367, net114368, net114369, net114370, net114371, net114372, 
      net114373, net114374, net114375, net114376, net114377, net114378, 
      net114379, net114380, net114381, net114382, net114383, net114384, 
      net114385, net114386, net114387, net114388, net114389, net114390, 
      net114391, net114392, net114393, net114394, net114395, net114396, 
      net114397, net114398, net114399, net114400, net114401, net114402, 
      net114403, net114404, net114405, net114406, net114407, net114408, 
      net114409, net114410, net114411, net114412, net114413, net114414, 
      net114415, net114416, net114417, net114418, net114419, net114433, 
      net114434, net114435, net114450, net114451, net114452, net114453, 
      net114454, net114455, net114456, net114457, net114458, net114459, 
      net114460, net114461, net114462, net114463, net114464, net114465, 
      net114466, net114467, net114468, net114469, net114470, net114471, 
      net114472, net114473, net114474, net114475, net114476, net114477, 
      net114478, net114479, net114480, net114481, net114482, net114483, 
      net114484, net114485, net114486, net114487, net114488, net114489, 
      net114490, net114491, net114492, net114493, net114494, net114495, 
      net114496, net114497, net114498, net114499, net114500, net114501, 
      net114502, net114503, net114504, net114505, net114506, net114507, 
      net114508, net114563, net114564, net114565, net114566, net114567, 
      net114568, net114569, net114570, net114571, net114572, net114573, 
      net114574, net114575, net114576, net114577, net114578, net114579, 
      net114580, net114581, net114582, net114583, net114584, net114585, 
      net114586, net114587, net114588, net114589, net114590, net114591, 
      net114592, net114593, net114594, net114595, net114596, net114597, 
      net114598, net114599, net114600, net114601, net114602, net114603, 
      net114604, net114605, net114606, net114607, net114608, net114609, 
      net114610, net114611, net114612, net114613, net114614, net114615, 
      net114616, net114617, net114618, net114619, net114620, net114621, 
      net114635, net114636, net114637, net114652, net114653, net114654, 
      net114655, net114656, net114657, net114658, net114659, net114660, 
      net114661, net114662, net114663, net114664, net114665, net114666, 
      net114667, net114668, net114669, net114670, net114671, net114672, 
      net114673, net114674, net114675, net114676, net114677, net114678, 
      net114679, net114680, net114681, net114682, net114683, net114684, 
      net114685, net114686, net114687, net114688, net114689, net114690, 
      net114691, net114692, net114693, net114694, net114695, net114696, 
      net114697, net114698, net114699, net114700, net114701, net114702, 
      net114703, net114704, net114705, net114706, net114707, net114708, 
      net114709, net114710, net114724, net114725, net114726, net114741, 
      net114742, net114743, net114744, net114745, net114746, net114747, 
      net114748, net114749, net114750, net114751, net114752, net114753, 
      net114754, net114755, net114756, net114757, net114758, net114759, 
      net114760, net114761, net114762, net114763, net114764, net114765, 
      net114766, net114767, net114768, net114769, net114770, net114771, 
      net114772, net114773, net114774, net114775, net114776, net114777, 
      net114778, net114779, net114780, net114781, net114782, net114783, 
      net114784, net114785, net114786, net114787, net114788, net114789, 
      net114790, net114791, net114792, net114793, net114794, net114795, 
      net114796, net114797, net114798, net114799, net114800, net114801, 
      net114802, net114803, net114804, net114805, net114806, net114807, 
      net114808, net114809, net114810, net114811, net114812, net114813, 
      net114814, net114815, net114816, net114817, net114818, net114819, 
      net114820, net114821, net114822, net114823, net114824, net114825, 
      net114826, net114827, net114828, net114829, net114830, net114831, 
      net114832, net114833, net114834, net114835, net114836, net114837, 
      net114838, net114839, net114840, net114841, net114842, net114843, 
      net114844, net114845, net114846, net114847, net114848, net114849, 
      net114850, net114851, net114852, net114853, net114854, net114855, 
      net114856, net114857, net114858, n3744, n3745, n3746, n3747, n3748, n3749
      , n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, 
      n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, 
      n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, 
      n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, 
      n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, 
      n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, 
      n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, 
      n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, 
      n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, 
      n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, 
      n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, 
      n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, 
      n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, 
      n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, 
      n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, 
      n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, 
      n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, 
      n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, 
      n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, 
      n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, 
      n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, 
      n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, 
      n3970, n3971, n3972, n3973, n3974, n3975, n3976, n_1006, n_1007, n_1008, 
      n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, n_1017, 
      n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, 
      n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, 
      n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, 
      n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, 
      n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, 
      n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, 
      n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, 
      n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, 
      n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, 
      n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, 
      n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116 : 
      std_logic;

begin
   OUTT_NT <= OUTT_NT_port;
   prevT_NT <= prevT_NT_port;
   
   n1 <= '0';
   prevT_NTs_reg : DFFR_X1 port map( D => OUTT_NT_port, CK => Clk, RN => n3894,
                           Q => prevT_NT_port, QN => net114858);
   pc_lut_reg_0_31_inst : DFFR_X1 port map( D => n7537, CK => Clk, RN => n3895,
                           Q => net114857, QN => n2241);
   pc_lut_reg_0_29_inst : DFFR_X1 port map( D => n7536, CK => Clk, RN => n3895,
                           Q => net114856, QN => n2240);
   pc_lut_reg_0_27_inst : DFFR_X1 port map( D => n7535, CK => Clk, RN => n3895,
                           Q => net114855, QN => n2239);
   pc_lut_reg_0_25_inst : DFFR_X1 port map( D => n7534, CK => Clk, RN => n3895,
                           Q => net114854, QN => n2238);
   pc_lut_reg_0_23_inst : DFFR_X1 port map( D => n7533, CK => Clk, RN => n3895,
                           Q => net114853, QN => n2237);
   pc_lut_reg_0_21_inst : DFFR_X1 port map( D => n7532, CK => Clk, RN => n3895,
                           Q => net114852, QN => n2236);
   pc_lut_reg_0_19_inst : DFFR_X1 port map( D => n7531, CK => Clk, RN => n3895,
                           Q => net114851, QN => n2235);
   pc_lut_reg_0_17_inst : DFFR_X1 port map( D => n7530, CK => Clk, RN => n3895,
                           Q => net114850, QN => n2234);
   pc_lut_reg_0_15_inst : DFFR_X1 port map( D => n7529, CK => Clk, RN => n3895,
                           Q => net114849, QN => n2233);
   pc_lut_reg_0_13_inst : DFFR_X1 port map( D => n7528, CK => Clk, RN => n3895,
                           Q => net114848, QN => n2232);
   pc_lut_reg_0_11_inst : DFFR_X1 port map( D => n7527, CK => Clk, RN => n3895,
                           Q => net114847, QN => n2231);
   pc_lut_reg_0_9_inst : DFFR_X1 port map( D => n7526, CK => Clk, RN => n3895, 
                           Q => net114846, QN => n2230);
   pc_lut_reg_0_7_inst : DFFR_X1 port map( D => n7525, CK => Clk, RN => n3895, 
                           Q => net114845, QN => n2229);
   pc_lut_reg_0_5_inst : DFFR_X1 port map( D => n7524, CK => Clk, RN => n3858, 
                           Q => net114844, QN => n2228);
   pc_lut_reg_0_6_inst : DFFR_X1 port map( D => n7518, CK => Clk, RN => n3895, 
                           Q => net114843, QN => n2222);
   pc_lut_reg_0_8_inst : DFFR_X1 port map( D => n7517, CK => Clk, RN => n3895, 
                           Q => net114842, QN => n2221);
   pc_lut_reg_0_10_inst : DFFR_X1 port map( D => n7516, CK => Clk, RN => n3896,
                           Q => net114841, QN => n2220);
   pc_lut_reg_0_12_inst : DFFR_X1 port map( D => n7515, CK => Clk, RN => n3896,
                           Q => net114840, QN => n2219);
   pc_lut_reg_0_14_inst : DFFR_X1 port map( D => n7514, CK => Clk, RN => n3896,
                           Q => net114839, QN => n2218);
   pc_lut_reg_0_16_inst : DFFR_X1 port map( D => n7513, CK => Clk, RN => n3896,
                           Q => net114838, QN => n2217);
   pc_lut_reg_0_18_inst : DFFR_X1 port map( D => n7512, CK => Clk, RN => n3861,
                           Q => net114837, QN => n2216);
   pc_lut_reg_0_20_inst : DFFR_X1 port map( D => n7511, CK => Clk, RN => n3896,
                           Q => net114836, QN => n2215);
   pc_lut_reg_0_22_inst : DFFR_X1 port map( D => n7510, CK => Clk, RN => n3896,
                           Q => net114835, QN => n2214);
   pc_lut_reg_0_24_inst : DFFR_X1 port map( D => n7509, CK => Clk, RN => n3896,
                           Q => net114834, QN => n2213);
   pc_lut_reg_0_26_inst : DFFR_X1 port map( D => n7508, CK => Clk, RN => n3916,
                           Q => net114833, QN => n2212);
   pc_lut_reg_0_28_inst : DFFR_X1 port map( D => n7507, CK => Clk, RN => n3912,
                           Q => net114832, QN => n2211);
   pc_lut_reg_0_30_inst : DFFR_X1 port map( D => n7506, CK => Clk, RN => n3912,
                           Q => net114831, QN => n2209);
   pc_lut_reg_1_31_inst : DFFR_X1 port map( D => n7505, CK => Clk, RN => n3913,
                           Q => net114830, QN => n2207);
   pc_lut_reg_1_29_inst : DFFR_X1 port map( D => n7504, CK => Clk, RN => n3913,
                           Q => net114829, QN => n2206);
   pc_lut_reg_1_27_inst : DFFR_X1 port map( D => n7503, CK => Clk, RN => n3913,
                           Q => net114828, QN => n2205);
   pc_lut_reg_1_25_inst : DFFR_X1 port map( D => n7502, CK => Clk, RN => n3913,
                           Q => net114827, QN => n2204);
   pc_lut_reg_1_23_inst : DFFR_X1 port map( D => n7501, CK => Clk, RN => n3913,
                           Q => net114826, QN => n2203);
   pc_lut_reg_1_21_inst : DFFR_X1 port map( D => n7500, CK => Clk, RN => n3913,
                           Q => net114825, QN => n2202);
   pc_lut_reg_1_19_inst : DFFR_X1 port map( D => n7499, CK => Clk, RN => n3913,
                           Q => net114824, QN => n2201);
   pc_lut_reg_1_17_inst : DFFR_X1 port map( D => n7498, CK => Clk, RN => n3913,
                           Q => net114823, QN => n2200);
   pc_lut_reg_1_15_inst : DFFR_X1 port map( D => n7497, CK => Clk, RN => n3913,
                           Q => net114822, QN => n2199);
   pc_lut_reg_1_13_inst : DFFR_X1 port map( D => n7496, CK => Clk, RN => n3913,
                           Q => net114821, QN => n2198);
   pc_lut_reg_1_11_inst : DFFR_X1 port map( D => n7495, CK => Clk, RN => n3913,
                           Q => net114820, QN => n2197);
   pc_lut_reg_1_9_inst : DFFR_X1 port map( D => n7494, CK => Clk, RN => n3913, 
                           Q => net114819, QN => n2196);
   pc_lut_reg_1_7_inst : DFFR_X1 port map( D => n7493, CK => Clk, RN => n3913, 
                           Q => net114818, QN => n2195);
   pc_lut_reg_1_5_inst : DFFR_X1 port map( D => n7492, CK => Clk, RN => n3858, 
                           Q => net114817, QN => n2194);
   pc_lut_reg_1_0_inst : DFFR_X1 port map( D => n7489, CK => Clk, RN => n3913, 
                           Q => net114816, QN => n2191);
   pc_lut_reg_1_6_inst : DFFR_X1 port map( D => n7486, CK => Clk, RN => n3913, 
                           Q => net114815, QN => n2188);
   pc_lut_reg_1_8_inst : DFFR_X1 port map( D => n7485, CK => Clk, RN => n3914, 
                           Q => net114814, QN => n2187);
   pc_lut_reg_1_10_inst : DFFR_X1 port map( D => n7484, CK => Clk, RN => n3914,
                           Q => net114813, QN => n2186);
   pc_lut_reg_1_12_inst : DFFR_X1 port map( D => n7483, CK => Clk, RN => n3914,
                           Q => net114812, QN => n2185);
   pc_lut_reg_1_14_inst : DFFR_X1 port map( D => n7482, CK => Clk, RN => n3914,
                           Q => net114811, QN => n2184);
   pc_lut_reg_1_16_inst : DFFR_X1 port map( D => n7481, CK => Clk, RN => n3914,
                           Q => net114810, QN => n2183);
   pc_lut_reg_1_18_inst : DFFR_X1 port map( D => n7480, CK => Clk, RN => n3861,
                           Q => net114809, QN => n2182);
   pc_lut_reg_1_20_inst : DFFR_X1 port map( D => n7479, CK => Clk, RN => n3914,
                           Q => net114808, QN => n2181);
   pc_lut_reg_1_22_inst : DFFR_X1 port map( D => n7478, CK => Clk, RN => n3914,
                           Q => net114807, QN => n2180);
   pc_lut_reg_1_24_inst : DFFR_X1 port map( D => n7477, CK => Clk, RN => n3914,
                           Q => net114806, QN => n2179);
   pc_lut_reg_1_26_inst : DFFR_X1 port map( D => n7476, CK => Clk, RN => n3914,
                           Q => net114805, QN => n2178);
   pc_lut_reg_1_28_inst : DFFR_X1 port map( D => n7475, CK => Clk, RN => n3914,
                           Q => net114804, QN => n2177);
   pc_lut_reg_1_30_inst : DFFR_X1 port map( D => n7474, CK => Clk, RN => n3914,
                           Q => net114803, QN => n2175);
   pc_lut_reg_2_31_inst : DFFR_X1 port map( D => n7473, CK => Clk, RN => n3914,
                           Q => pc_lut_2_31_port, QN => n2173);
   pc_lut_reg_2_29_inst : DFFR_X1 port map( D => n7472, CK => Clk, RN => n3914,
                           Q => pc_lut_2_29_port, QN => n2172);
   pc_lut_reg_2_27_inst : DFFR_X1 port map( D => n7471, CK => Clk, RN => n3914,
                           Q => pc_lut_2_27_port, QN => n2171);
   pc_lut_reg_2_25_inst : DFFR_X1 port map( D => n7470, CK => Clk, RN => n3914,
                           Q => pc_lut_2_25_port, QN => n2170);
   pc_lut_reg_2_23_inst : DFFR_X1 port map( D => n7469, CK => Clk, RN => n3915,
                           Q => pc_lut_2_23_port, QN => n2169);
   pc_lut_reg_2_21_inst : DFFR_X1 port map( D => n7468, CK => Clk, RN => n3915,
                           Q => pc_lut_2_21_port, QN => n2168);
   pc_lut_reg_2_19_inst : DFFR_X1 port map( D => n7467, CK => Clk, RN => n3915,
                           Q => pc_lut_2_19_port, QN => n2167);
   pc_lut_reg_2_17_inst : DFFR_X1 port map( D => n7466, CK => Clk, RN => n3915,
                           Q => pc_lut_2_17_port, QN => n2166);
   pc_lut_reg_2_15_inst : DFFR_X1 port map( D => n7465, CK => Clk, RN => n3915,
                           Q => pc_lut_2_15_port, QN => n2165);
   pc_lut_reg_2_13_inst : DFFR_X1 port map( D => n7464, CK => Clk, RN => n3915,
                           Q => pc_lut_2_13_port, QN => n2164);
   pc_lut_reg_2_11_inst : DFFR_X1 port map( D => n7463, CK => Clk, RN => n3915,
                           Q => pc_lut_2_11_port, QN => n2163);
   pc_lut_reg_2_9_inst : DFFR_X1 port map( D => n7462, CK => Clk, RN => n3915, 
                           Q => pc_lut_2_9_port, QN => n2162);
   pc_lut_reg_2_7_inst : DFFR_X1 port map( D => n7461, CK => Clk, RN => n3915, 
                           Q => pc_lut_2_7_port, QN => n2161);
   pc_lut_reg_2_5_inst : DFFR_X1 port map( D => n7460, CK => Clk, RN => n3858, 
                           Q => pc_lut_2_5_port, QN => n2160);
   pc_lut_reg_2_1_inst : DFFR_X1 port map( D => n7458, CK => Clk, RN => n3915, 
                           Q => pc_lut_2_1_port, QN => net114802);
   pc_lut_reg_2_6_inst : DFFR_X1 port map( D => n7454, CK => Clk, RN => n3915, 
                           Q => pc_lut_2_6_port, QN => n2158);
   pc_lut_reg_2_8_inst : DFFR_X1 port map( D => n7453, CK => Clk, RN => n3915, 
                           Q => pc_lut_2_8_port, QN => n2157);
   pc_lut_reg_2_10_inst : DFFR_X1 port map( D => n7452, CK => Clk, RN => n3915,
                           Q => pc_lut_2_10_port, QN => n2156);
   pc_lut_reg_2_12_inst : DFFR_X1 port map( D => n7451, CK => Clk, RN => n3915,
                           Q => pc_lut_2_12_port, QN => n2155);
   pc_lut_reg_2_14_inst : DFFR_X1 port map( D => n7450, CK => Clk, RN => n3915,
                           Q => pc_lut_2_14_port, QN => n2154);
   pc_lut_reg_2_16_inst : DFFR_X1 port map( D => n7449, CK => Clk, RN => n3916,
                           Q => pc_lut_2_16_port, QN => n2153);
   pc_lut_reg_2_18_inst : DFFR_X1 port map( D => n7448, CK => Clk, RN => n3861,
                           Q => pc_lut_2_18_port, QN => n2152);
   pc_lut_reg_2_20_inst : DFFR_X1 port map( D => n7447, CK => Clk, RN => n3916,
                           Q => pc_lut_2_20_port, QN => n2151);
   pc_lut_reg_2_22_inst : DFFR_X1 port map( D => n7446, CK => Clk, RN => n3916,
                           Q => pc_lut_2_22_port, QN => n2150);
   pc_lut_reg_2_24_inst : DFFR_X1 port map( D => n7445, CK => Clk, RN => n3916,
                           Q => pc_lut_2_24_port, QN => n2149);
   pc_lut_reg_2_26_inst : DFFR_X1 port map( D => n7444, CK => Clk, RN => n3916,
                           Q => pc_lut_2_26_port, QN => n2148);
   pc_lut_reg_2_28_inst : DFFR_X1 port map( D => n7443, CK => Clk, RN => n3916,
                           Q => pc_lut_2_28_port, QN => n2147);
   pc_lut_reg_2_30_inst : DFFR_X1 port map( D => n7442, CK => Clk, RN => n3916,
                           Q => pc_lut_2_30_port, QN => n2145);
   pc_lut_reg_3_31_inst : DFFR_X1 port map( D => n7441, CK => Clk, RN => n3916,
                           Q => pc_lut_3_31_port, QN => n2140);
   pc_lut_reg_3_29_inst : DFFR_X1 port map( D => n7440, CK => Clk, RN => n3916,
                           Q => pc_lut_3_29_port, QN => n2139);
   pc_lut_reg_3_27_inst : DFFR_X1 port map( D => n7439, CK => Clk, RN => n3916,
                           Q => pc_lut_3_27_port, QN => n2138);
   pc_lut_reg_3_25_inst : DFFR_X1 port map( D => n7438, CK => Clk, RN => n3916,
                           Q => pc_lut_3_25_port, QN => n2137);
   pc_lut_reg_3_23_inst : DFFR_X1 port map( D => n7437, CK => Clk, RN => n3916,
                           Q => pc_lut_3_23_port, QN => n2136);
   pc_lut_reg_3_21_inst : DFFR_X1 port map( D => n7436, CK => Clk, RN => n3916,
                           Q => pc_lut_3_21_port, QN => n2135);
   pc_lut_reg_3_19_inst : DFFR_X1 port map( D => n7435, CK => Clk, RN => n3916,
                           Q => pc_lut_3_19_port, QN => n2134);
   pc_lut_reg_3_17_inst : DFFR_X1 port map( D => n7434, CK => Clk, RN => n3917,
                           Q => pc_lut_3_17_port, QN => n2133);
   pc_lut_reg_3_15_inst : DFFR_X1 port map( D => n7433, CK => Clk, RN => n3917,
                           Q => pc_lut_3_15_port, QN => n2132);
   pc_lut_reg_3_13_inst : DFFR_X1 port map( D => n7432, CK => Clk, RN => n3917,
                           Q => pc_lut_3_13_port, QN => n2131);
   pc_lut_reg_3_11_inst : DFFR_X1 port map( D => n7431, CK => Clk, RN => n3917,
                           Q => pc_lut_3_11_port, QN => n2130);
   pc_lut_reg_3_9_inst : DFFR_X1 port map( D => n7430, CK => Clk, RN => n3917, 
                           Q => pc_lut_3_9_port, QN => n2129);
   pc_lut_reg_3_7_inst : DFFR_X1 port map( D => n7429, CK => Clk, RN => n3917, 
                           Q => pc_lut_3_7_port, QN => n2128);
   pc_lut_reg_3_5_inst : DFFR_X1 port map( D => n7428, CK => Clk, RN => n3858, 
                           Q => pc_lut_3_5_port, QN => n2127);
   pc_lut_reg_3_1_inst : DFFR_X1 port map( D => n7426, CK => Clk, RN => n3917, 
                           Q => pc_lut_3_1_port, QN => net114801);
   pc_lut_reg_3_0_inst : DFFR_X1 port map( D => n7425, CK => Clk, RN => n3917, 
                           Q => pc_lut_3_0_port, QN => net114800);
   pc_lut_reg_3_6_inst : DFFR_X1 port map( D => n7422, CK => Clk, RN => n3917, 
                           Q => pc_lut_3_6_port, QN => n2124);
   pc_lut_reg_3_8_inst : DFFR_X1 port map( D => n7421, CK => Clk, RN => n3917, 
                           Q => pc_lut_3_8_port, QN => n2123);
   pc_lut_reg_3_10_inst : DFFR_X1 port map( D => n7420, CK => Clk, RN => n3917,
                           Q => pc_lut_3_10_port, QN => n2122);
   pc_lut_reg_3_12_inst : DFFR_X1 port map( D => n7419, CK => Clk, RN => n3917,
                           Q => pc_lut_3_12_port, QN => n2121);
   pc_lut_reg_3_14_inst : DFFR_X1 port map( D => n7418, CK => Clk, RN => n3917,
                           Q => pc_lut_3_14_port, QN => n2120);
   pc_lut_reg_3_16_inst : DFFR_X1 port map( D => n7417, CK => Clk, RN => n3917,
                           Q => pc_lut_3_16_port, QN => n2119);
   pc_lut_reg_3_18_inst : DFFR_X1 port map( D => n7416, CK => Clk, RN => n3861,
                           Q => pc_lut_3_18_port, QN => n2118);
   pc_lut_reg_3_20_inst : DFFR_X1 port map( D => n7415, CK => Clk, RN => n3917,
                           Q => pc_lut_3_20_port, QN => n2117);
   pc_lut_reg_3_22_inst : DFFR_X1 port map( D => n7414, CK => Clk, RN => n3918,
                           Q => pc_lut_3_22_port, QN => n2116);
   pc_lut_reg_3_24_inst : DFFR_X1 port map( D => n7413, CK => Clk, RN => n3918,
                           Q => pc_lut_3_24_port, QN => n2115);
   pc_lut_reg_3_26_inst : DFFR_X1 port map( D => n7412, CK => Clk, RN => n3918,
                           Q => pc_lut_3_26_port, QN => n2114);
   pc_lut_reg_3_28_inst : DFFR_X1 port map( D => n7411, CK => Clk, RN => n3918,
                           Q => pc_lut_3_28_port, QN => n2113);
   pc_lut_reg_3_30_inst : DFFR_X1 port map( D => n7410, CK => Clk, RN => n3918,
                           Q => pc_lut_3_30_port, QN => n2111);
   pc_lut_reg_4_31_inst : DFFR_X1 port map( D => n7409, CK => Clk, RN => n3918,
                           Q => net114799, QN => n2109);
   pc_lut_reg_4_29_inst : DFFR_X1 port map( D => n7408, CK => Clk, RN => n3918,
                           Q => net114798, QN => n2108);
   pc_lut_reg_4_27_inst : DFFR_X1 port map( D => n7407, CK => Clk, RN => n3918,
                           Q => net114797, QN => n2107);
   pc_lut_reg_4_25_inst : DFFR_X1 port map( D => n7406, CK => Clk, RN => n3918,
                           Q => net114796, QN => n2106);
   pc_lut_reg_4_23_inst : DFFR_X1 port map( D => n7405, CK => Clk, RN => n3918,
                           Q => net114795, QN => n2105);
   pc_lut_reg_4_21_inst : DFFR_X1 port map( D => n7404, CK => Clk, RN => n3918,
                           Q => net114794, QN => n2104);
   pc_lut_reg_4_19_inst : DFFR_X1 port map( D => n7403, CK => Clk, RN => n3918,
                           Q => net114793, QN => n2103);
   pc_lut_reg_4_17_inst : DFFR_X1 port map( D => n7402, CK => Clk, RN => n3918,
                           Q => net114792, QN => n2102);
   pc_lut_reg_4_15_inst : DFFR_X1 port map( D => n7401, CK => Clk, RN => n3918,
                           Q => net114791, QN => n2101);
   pc_lut_reg_4_13_inst : DFFR_X1 port map( D => n7400, CK => Clk, RN => n3918,
                           Q => net114790, QN => n2100);
   pc_lut_reg_4_11_inst : DFFR_X1 port map( D => n7399, CK => Clk, RN => n3919,
                           Q => net114789, QN => n2099);
   pc_lut_reg_4_9_inst : DFFR_X1 port map( D => n7398, CK => Clk, RN => n3919, 
                           Q => net114788, QN => n2098);
   pc_lut_reg_4_7_inst : DFFR_X1 port map( D => n7397, CK => Clk, RN => n3919, 
                           Q => net114787, QN => n2097);
   pc_lut_reg_4_5_inst : DFFR_X1 port map( D => n7396, CK => Clk, RN => n3859, 
                           Q => net114786, QN => n2096);
   pc_lut_reg_4_2_inst : DFFR_X1 port map( D => n7392, CK => Clk, RN => n3919, 
                           Q => net114785, QN => n2092);
   pc_lut_reg_4_6_inst : DFFR_X1 port map( D => n7390, CK => Clk, RN => n3919, 
                           Q => net114784, QN => n2090);
   pc_lut_reg_4_8_inst : DFFR_X1 port map( D => n7389, CK => Clk, RN => n3919, 
                           Q => net114783, QN => n2089);
   pc_lut_reg_4_10_inst : DFFR_X1 port map( D => n7388, CK => Clk, RN => n3919,
                           Q => net114782, QN => n2088);
   pc_lut_reg_4_12_inst : DFFR_X1 port map( D => n7387, CK => Clk, RN => n3919,
                           Q => net114781, QN => n2087);
   pc_lut_reg_4_14_inst : DFFR_X1 port map( D => n7386, CK => Clk, RN => n3919,
                           Q => net114780, QN => n2086);
   pc_lut_reg_4_16_inst : DFFR_X1 port map( D => n7385, CK => Clk, RN => n3919,
                           Q => net114779, QN => n2085);
   pc_lut_reg_4_18_inst : DFFR_X1 port map( D => n7384, CK => Clk, RN => n3862,
                           Q => net114778, QN => n2084);
   pc_lut_reg_4_20_inst : DFFR_X1 port map( D => n7383, CK => Clk, RN => n3919,
                           Q => net114777, QN => n2083);
   pc_lut_reg_4_22_inst : DFFR_X1 port map( D => n7382, CK => Clk, RN => n3919,
                           Q => net114776, QN => n2082);
   pc_lut_reg_4_24_inst : DFFR_X1 port map( D => n7381, CK => Clk, RN => n3919,
                           Q => net114775, QN => n2081);
   pc_lut_reg_4_26_inst : DFFR_X1 port map( D => n7380, CK => Clk, RN => n3919,
                           Q => net114774, QN => n2080);
   pc_lut_reg_4_28_inst : DFFR_X1 port map( D => n7379, CK => Clk, RN => n3920,
                           Q => net114773, QN => n2079);
   pc_lut_reg_4_30_inst : DFFR_X1 port map( D => n7378, CK => Clk, RN => n3920,
                           Q => net114772, QN => n2077);
   pc_lut_reg_5_31_inst : DFFR_X1 port map( D => n7377, CK => Clk, RN => n3919,
                           Q => net114771, QN => n2075);
   pc_lut_reg_5_29_inst : DFFR_X1 port map( D => n7376, CK => Clk, RN => n3920,
                           Q => net114770, QN => n2074);
   pc_lut_reg_5_27_inst : DFFR_X1 port map( D => n7375, CK => Clk, RN => n3920,
                           Q => net114769, QN => n2073);
   pc_lut_reg_5_25_inst : DFFR_X1 port map( D => n7374, CK => Clk, RN => n3920,
                           Q => net114768, QN => n2072);
   pc_lut_reg_5_23_inst : DFFR_X1 port map( D => n7373, CK => Clk, RN => n3920,
                           Q => net114767, QN => n2071);
   pc_lut_reg_5_21_inst : DFFR_X1 port map( D => n7372, CK => Clk, RN => n3920,
                           Q => net114766, QN => n2070);
   pc_lut_reg_5_19_inst : DFFR_X1 port map( D => n7371, CK => Clk, RN => n3920,
                           Q => net114765, QN => n2069);
   pc_lut_reg_5_17_inst : DFFR_X1 port map( D => n7370, CK => Clk, RN => n3920,
                           Q => net114764, QN => n2068);
   pc_lut_reg_5_15_inst : DFFR_X1 port map( D => n7369, CK => Clk, RN => n3920,
                           Q => net114763, QN => n2067);
   pc_lut_reg_5_13_inst : DFFR_X1 port map( D => n7368, CK => Clk, RN => n3920,
                           Q => net114762, QN => n2066);
   pc_lut_reg_5_11_inst : DFFR_X1 port map( D => n7367, CK => Clk, RN => n3920,
                           Q => net114761, QN => n2065);
   pc_lut_reg_5_9_inst : DFFR_X1 port map( D => n7366, CK => Clk, RN => n3920, 
                           Q => net114760, QN => n2064);
   pc_lut_reg_5_7_inst : DFFR_X1 port map( D => n7365, CK => Clk, RN => n3920, 
                           Q => net114759, QN => n2063);
   pc_lut_reg_5_5_inst : DFFR_X1 port map( D => n7364, CK => Clk, RN => n3859, 
                           Q => net114758, QN => n2062);
   pc_lut_reg_5_0_inst : DFFR_X1 port map( D => n7361, CK => Clk, RN => n3920, 
                           Q => net114757, QN => n2059);
   pc_lut_reg_5_2_inst : DFFR_X1 port map( D => n7360, CK => Clk, RN => n3908, 
                           Q => net114756, QN => n2058);
   pc_lut_reg_5_6_inst : DFFR_X1 port map( D => n7358, CK => Clk, RN => n3904, 
                           Q => net114755, QN => n2056);
   pc_lut_reg_5_8_inst : DFFR_X1 port map( D => n7357, CK => Clk, RN => n3904, 
                           Q => net114754, QN => n2055);
   pc_lut_reg_5_10_inst : DFFR_X1 port map( D => n7356, CK => Clk, RN => n3904,
                           Q => net114753, QN => n2054);
   pc_lut_reg_5_12_inst : DFFR_X1 port map( D => n7355, CK => Clk, RN => n3904,
                           Q => net114752, QN => n2053);
   pc_lut_reg_5_14_inst : DFFR_X1 port map( D => n7354, CK => Clk, RN => n3904,
                           Q => net114751, QN => n2052);
   pc_lut_reg_5_16_inst : DFFR_X1 port map( D => n7353, CK => Clk, RN => n3905,
                           Q => net114750, QN => n2051);
   pc_lut_reg_5_18_inst : DFFR_X1 port map( D => n7352, CK => Clk, RN => n3862,
                           Q => net114749, QN => n2050);
   pc_lut_reg_5_20_inst : DFFR_X1 port map( D => n7351, CK => Clk, RN => n3905,
                           Q => net114748, QN => n2049);
   pc_lut_reg_5_22_inst : DFFR_X1 port map( D => n7350, CK => Clk, RN => n3905,
                           Q => net114747, QN => n2048);
   pc_lut_reg_5_24_inst : DFFR_X1 port map( D => n7349, CK => Clk, RN => n3905,
                           Q => net114746, QN => n2047);
   pc_lut_reg_5_26_inst : DFFR_X1 port map( D => n7348, CK => Clk, RN => n3905,
                           Q => net114745, QN => n2046);
   pc_lut_reg_5_28_inst : DFFR_X1 port map( D => n7347, CK => Clk, RN => n3905,
                           Q => net114744, QN => n2045);
   pc_lut_reg_5_30_inst : DFFR_X1 port map( D => n7346, CK => Clk, RN => n3905,
                           Q => net114743, QN => n2043);
   pc_lut_reg_6_31_inst : DFFR_X1 port map( D => n7345, CK => Clk, RN => n3905,
                           Q => pc_lut_6_31_port, QN => n2041);
   pc_lut_reg_6_29_inst : DFFR_X1 port map( D => n7344, CK => Clk, RN => n3905,
                           Q => pc_lut_6_29_port, QN => n2040);
   pc_lut_reg_6_27_inst : DFFR_X1 port map( D => n7343, CK => Clk, RN => n3905,
                           Q => pc_lut_6_27_port, QN => n2039);
   pc_lut_reg_6_25_inst : DFFR_X1 port map( D => n7342, CK => Clk, RN => n3905,
                           Q => pc_lut_6_25_port, QN => n2038);
   pc_lut_reg_6_23_inst : DFFR_X1 port map( D => n7341, CK => Clk, RN => n3905,
                           Q => pc_lut_6_23_port, QN => n2037);
   pc_lut_reg_6_21_inst : DFFR_X1 port map( D => n7340, CK => Clk, RN => n3905,
                           Q => pc_lut_6_21_port, QN => n2036);
   pc_lut_reg_6_19_inst : DFFR_X1 port map( D => n7339, CK => Clk, RN => n3905,
                           Q => pc_lut_6_19_port, QN => n2035);
   pc_lut_reg_6_17_inst : DFFR_X1 port map( D => n7338, CK => Clk, RN => n3905,
                           Q => pc_lut_6_17_port, QN => n2034);
   pc_lut_reg_6_15_inst : DFFR_X1 port map( D => n7337, CK => Clk, RN => n3906,
                           Q => pc_lut_6_15_port, QN => n2033);
   pc_lut_reg_6_13_inst : DFFR_X1 port map( D => n7336, CK => Clk, RN => n3906,
                           Q => pc_lut_6_13_port, QN => n2032);
   pc_lut_reg_6_11_inst : DFFR_X1 port map( D => n7335, CK => Clk, RN => n3906,
                           Q => pc_lut_6_11_port, QN => n2031);
   pc_lut_reg_6_9_inst : DFFR_X1 port map( D => n7334, CK => Clk, RN => n3906, 
                           Q => pc_lut_6_9_port, QN => n2030);
   pc_lut_reg_6_7_inst : DFFR_X1 port map( D => n7333, CK => Clk, RN => n3906, 
                           Q => pc_lut_6_7_port, QN => n2029);
   pc_lut_reg_6_5_inst : DFFR_X1 port map( D => n7332, CK => Clk, RN => n3859, 
                           Q => pc_lut_6_5_port, QN => n2028);
   pc_lut_reg_6_1_inst : DFFR_X1 port map( D => n7330, CK => Clk, RN => n3906, 
                           Q => pc_lut_6_1_port, QN => net114742);
   pc_lut_reg_6_2_inst : DFFR_X1 port map( D => n7328, CK => Clk, RN => n3906, 
                           Q => pc_lut_6_2_port, QN => net114741);
   pc_lut_reg_6_6_inst : DFFR_X1 port map( D => n7326, CK => Clk, RN => n3906, 
                           Q => pc_lut_6_6_port, QN => n2025);
   pc_lut_reg_6_8_inst : DFFR_X1 port map( D => n7325, CK => Clk, RN => n3906, 
                           Q => pc_lut_6_8_port, QN => n2024);
   pc_lut_reg_6_10_inst : DFFR_X1 port map( D => n7324, CK => Clk, RN => n3906,
                           Q => pc_lut_6_10_port, QN => n2023);
   pc_lut_reg_6_12_inst : DFFR_X1 port map( D => n7323, CK => Clk, RN => n3906,
                           Q => pc_lut_6_12_port, QN => n2022);
   pc_lut_reg_6_14_inst : DFFR_X1 port map( D => n7322, CK => Clk, RN => n3906,
                           Q => pc_lut_6_14_port, QN => n2021);
   pc_lut_reg_6_16_inst : DFFR_X1 port map( D => n7321, CK => Clk, RN => n3906,
                           Q => pc_lut_6_16_port, QN => n2020);
   pc_lut_reg_6_18_inst : DFFR_X1 port map( D => n7320, CK => Clk, RN => n3862,
                           Q => pc_lut_6_18_port, QN => n2019);
   pc_lut_reg_6_20_inst : DFFR_X1 port map( D => n7319, CK => Clk, RN => n3906,
                           Q => pc_lut_6_20_port, QN => n2018);
   pc_lut_reg_6_22_inst : DFFR_X1 port map( D => n7318, CK => Clk, RN => n3906,
                           Q => pc_lut_6_22_port, QN => n2017);
   pc_lut_reg_6_24_inst : DFFR_X1 port map( D => n7317, CK => Clk, RN => n3907,
                           Q => pc_lut_6_24_port, QN => n2016);
   pc_lut_reg_6_26_inst : DFFR_X1 port map( D => n7316, CK => Clk, RN => n3907,
                           Q => pc_lut_6_26_port, QN => n2015);
   pc_lut_reg_6_28_inst : DFFR_X1 port map( D => n7315, CK => Clk, RN => n3907,
                           Q => pc_lut_6_28_port, QN => n2014);
   pc_lut_reg_6_30_inst : DFFR_X1 port map( D => n7314, CK => Clk, RN => n3907,
                           Q => pc_lut_6_30_port, QN => n2012);
   pc_lut_reg_7_31_inst : DFFR_X1 port map( D => n7313, CK => Clk, RN => n3907,
                           Q => pc_lut_7_31_port, QN => n2009);
   pc_lut_reg_7_29_inst : DFFR_X1 port map( D => n7312, CK => Clk, RN => n3907,
                           Q => pc_lut_7_29_port, QN => n2008);
   pc_lut_reg_7_27_inst : DFFR_X1 port map( D => n7311, CK => Clk, RN => n3907,
                           Q => pc_lut_7_27_port, QN => n2007);
   pc_lut_reg_7_25_inst : DFFR_X1 port map( D => n7310, CK => Clk, RN => n3907,
                           Q => pc_lut_7_25_port, QN => n2006);
   pc_lut_reg_7_23_inst : DFFR_X1 port map( D => n7309, CK => Clk, RN => n3907,
                           Q => pc_lut_7_23_port, QN => n2005);
   pc_lut_reg_7_21_inst : DFFR_X1 port map( D => n7308, CK => Clk, RN => n3907,
                           Q => pc_lut_7_21_port, QN => n2004);
   pc_lut_reg_7_19_inst : DFFR_X1 port map( D => n7307, CK => Clk, RN => n3907,
                           Q => pc_lut_7_19_port, QN => n2003);
   pc_lut_reg_7_17_inst : DFFR_X1 port map( D => n7306, CK => Clk, RN => n3907,
                           Q => pc_lut_7_17_port, QN => n2002);
   pc_lut_reg_7_15_inst : DFFR_X1 port map( D => n7305, CK => Clk, RN => n3907,
                           Q => pc_lut_7_15_port, QN => n2001);
   pc_lut_reg_7_13_inst : DFFR_X1 port map( D => n7304, CK => Clk, RN => n3907,
                           Q => pc_lut_7_13_port, QN => n2000);
   pc_lut_reg_7_11_inst : DFFR_X1 port map( D => n7303, CK => Clk, RN => n3907,
                           Q => pc_lut_7_11_port, QN => n1999);
   pc_lut_reg_7_9_inst : DFFR_X1 port map( D => n7302, CK => Clk, RN => n3908, 
                           Q => pc_lut_7_9_port, QN => n1998);
   pc_lut_reg_7_7_inst : DFFR_X1 port map( D => n7301, CK => Clk, RN => n3908, 
                           Q => pc_lut_7_7_port, QN => n1997);
   pc_lut_reg_7_5_inst : DFFR_X1 port map( D => n7300, CK => Clk, RN => n3859, 
                           Q => pc_lut_7_5_port, QN => n1996);
   pc_lut_reg_7_1_inst : DFFR_X1 port map( D => n7298, CK => Clk, RN => n3908, 
                           Q => pc_lut_7_1_port, QN => net114726);
   pc_lut_reg_7_0_inst : DFFR_X1 port map( D => n7297, CK => Clk, RN => n3908, 
                           Q => pc_lut_7_0_port, QN => net114725);
   pc_lut_reg_7_2_inst : DFFR_X1 port map( D => n7296, CK => Clk, RN => n3908, 
                           Q => pc_lut_7_2_port, QN => net114724);
   pc_lut_reg_7_6_inst : DFFR_X1 port map( D => n7294, CK => Clk, RN => n3908, 
                           Q => pc_lut_7_6_port, QN => n1992);
   pc_lut_reg_7_8_inst : DFFR_X1 port map( D => n7293, CK => Clk, RN => n3908, 
                           Q => pc_lut_7_8_port, QN => n1991);
   pc_lut_reg_7_10_inst : DFFR_X1 port map( D => n7292, CK => Clk, RN => n3908,
                           Q => pc_lut_7_10_port, QN => n1990);
   pc_lut_reg_7_12_inst : DFFR_X1 port map( D => n7291, CK => Clk, RN => n3897,
                           Q => pc_lut_7_12_port, QN => n1989);
   pc_lut_reg_7_14_inst : DFFR_X1 port map( D => n7290, CK => Clk, RN => n3897,
                           Q => pc_lut_7_14_port, QN => n1988);
   pc_lut_reg_7_16_inst : DFFR_X1 port map( D => n7289, CK => Clk, RN => n3897,
                           Q => pc_lut_7_16_port, QN => n1987);
   pc_lut_reg_7_18_inst : DFFR_X1 port map( D => n7288, CK => Clk, RN => n3862,
                           Q => pc_lut_7_18_port, QN => n1986);
   pc_lut_reg_7_20_inst : DFFR_X1 port map( D => n7287, CK => Clk, RN => n3897,
                           Q => pc_lut_7_20_port, QN => n1985);
   pc_lut_reg_7_22_inst : DFFR_X1 port map( D => n7286, CK => Clk, RN => n3897,
                           Q => pc_lut_7_22_port, QN => n1984);
   pc_lut_reg_7_24_inst : DFFR_X1 port map( D => n7285, CK => Clk, RN => n3897,
                           Q => pc_lut_7_24_port, QN => n1983);
   pc_lut_reg_7_26_inst : DFFR_X1 port map( D => n7284, CK => Clk, RN => n3897,
                           Q => pc_lut_7_26_port, QN => n1982);
   pc_lut_reg_7_28_inst : DFFR_X1 port map( D => n7283, CK => Clk, RN => n3897,
                           Q => pc_lut_7_28_port, QN => n1981);
   pc_lut_reg_7_30_inst : DFFR_X1 port map( D => n7282, CK => Clk, RN => n3897,
                           Q => pc_lut_7_30_port, QN => n1979);
   pc_lut_reg_8_31_inst : DFFR_X1 port map( D => n7281, CK => Clk, RN => n3897,
                           Q => net114710, QN => n1977);
   pc_lut_reg_8_29_inst : DFFR_X1 port map( D => n7280, CK => Clk, RN => n3897,
                           Q => net114709, QN => n1976);
   pc_lut_reg_8_27_inst : DFFR_X1 port map( D => n7279, CK => Clk, RN => n3897,
                           Q => net114708, QN => n1975);
   pc_lut_reg_8_25_inst : DFFR_X1 port map( D => n7278, CK => Clk, RN => n3897,
                           Q => net114707, QN => n1974);
   pc_lut_reg_8_23_inst : DFFR_X1 port map( D => n7277, CK => Clk, RN => n3898,
                           Q => net114706, QN => n1973);
   pc_lut_reg_8_21_inst : DFFR_X1 port map( D => n7276, CK => Clk, RN => n3898,
                           Q => net114705, QN => n1972);
   pc_lut_reg_8_19_inst : DFFR_X1 port map( D => n7275, CK => Clk, RN => n3898,
                           Q => net114704, QN => n1971);
   pc_lut_reg_8_17_inst : DFFR_X1 port map( D => n7274, CK => Clk, RN => n3898,
                           Q => net114703, QN => n1970);
   pc_lut_reg_8_15_inst : DFFR_X1 port map( D => n7273, CK => Clk, RN => n3898,
                           Q => net114702, QN => n1969);
   pc_lut_reg_8_13_inst : DFFR_X1 port map( D => n7272, CK => Clk, RN => n3898,
                           Q => net114701, QN => n1968);
   pc_lut_reg_8_11_inst : DFFR_X1 port map( D => n7271, CK => Clk, RN => n3898,
                           Q => net114700, QN => n1967);
   pc_lut_reg_8_9_inst : DFFR_X1 port map( D => n7270, CK => Clk, RN => n3898, 
                           Q => net114699, QN => n1966);
   pc_lut_reg_8_7_inst : DFFR_X1 port map( D => n7269, CK => Clk, RN => n3898, 
                           Q => net114698, QN => n1965);
   pc_lut_reg_8_5_inst : DFFR_X1 port map( D => n7268, CK => Clk, RN => n3859, 
                           Q => net114697, QN => n1964);
   pc_lut_reg_8_3_inst : DFFR_X1 port map( D => n7267, CK => Clk, RN => n3898, 
                           Q => net114696, QN => n1963);
   pc_lut_reg_8_6_inst : DFFR_X1 port map( D => n7262, CK => Clk, RN => n3898, 
                           Q => net114695, QN => n1958);
   pc_lut_reg_8_8_inst : DFFR_X1 port map( D => n7261, CK => Clk, RN => n3898, 
                           Q => net114694, QN => n1957);
   pc_lut_reg_8_10_inst : DFFR_X1 port map( D => n7260, CK => Clk, RN => n3898,
                           Q => net114693, QN => n1956);
   pc_lut_reg_8_12_inst : DFFR_X1 port map( D => n7259, CK => Clk, RN => n3898,
                           Q => net114692, QN => n1955);
   pc_lut_reg_8_14_inst : DFFR_X1 port map( D => n7258, CK => Clk, RN => n3899,
                           Q => net114691, QN => n1954);
   pc_lut_reg_8_16_inst : DFFR_X1 port map( D => n7257, CK => Clk, RN => n3899,
                           Q => net114690, QN => n1953);
   pc_lut_reg_8_18_inst : DFFR_X1 port map( D => n7256, CK => Clk, RN => n3862,
                           Q => net114689, QN => n1952);
   pc_lut_reg_8_20_inst : DFFR_X1 port map( D => n7255, CK => Clk, RN => n3899,
                           Q => net114688, QN => n1951);
   pc_lut_reg_8_22_inst : DFFR_X1 port map( D => n7254, CK => Clk, RN => n3899,
                           Q => net114687, QN => n1950);
   pc_lut_reg_8_24_inst : DFFR_X1 port map( D => n7253, CK => Clk, RN => n3899,
                           Q => net114686, QN => n1949);
   pc_lut_reg_8_26_inst : DFFR_X1 port map( D => n7252, CK => Clk, RN => n3899,
                           Q => net114685, QN => n1948);
   pc_lut_reg_8_28_inst : DFFR_X1 port map( D => n7251, CK => Clk, RN => n3899,
                           Q => net114684, QN => n1947);
   pc_lut_reg_8_30_inst : DFFR_X1 port map( D => n7250, CK => Clk, RN => n3899,
                           Q => net114683, QN => n1945);
   pc_lut_reg_9_31_inst : DFFR_X1 port map( D => n7249, CK => Clk, RN => n3898,
                           Q => net114682, QN => n1943);
   pc_lut_reg_9_29_inst : DFFR_X1 port map( D => n7248, CK => Clk, RN => n3899,
                           Q => net114681, QN => n1942);
   pc_lut_reg_9_27_inst : DFFR_X1 port map( D => n7247, CK => Clk, RN => n3899,
                           Q => net114680, QN => n1941);
   pc_lut_reg_9_25_inst : DFFR_X1 port map( D => n7246, CK => Clk, RN => n3899,
                           Q => net114679, QN => n1940);
   pc_lut_reg_9_23_inst : DFFR_X1 port map( D => n7245, CK => Clk, RN => n3899,
                           Q => net114678, QN => n1939);
   pc_lut_reg_9_21_inst : DFFR_X1 port map( D => n7244, CK => Clk, RN => n3899,
                           Q => net114677, QN => n1938);
   pc_lut_reg_9_19_inst : DFFR_X1 port map( D => n7243, CK => Clk, RN => n3899,
                           Q => net114676, QN => n1937);
   pc_lut_reg_9_17_inst : DFFR_X1 port map( D => n7242, CK => Clk, RN => n3899,
                           Q => net114675, QN => n1936);
   pc_lut_reg_9_15_inst : DFFR_X1 port map( D => n7241, CK => Clk, RN => n3900,
                           Q => net114674, QN => n1935);
   pc_lut_reg_9_13_inst : DFFR_X1 port map( D => n7240, CK => Clk, RN => n3900,
                           Q => net114673, QN => n1934);
   pc_lut_reg_9_11_inst : DFFR_X1 port map( D => n7239, CK => Clk, RN => n3900,
                           Q => net114672, QN => n1933);
   pc_lut_reg_9_9_inst : DFFR_X1 port map( D => n7238, CK => Clk, RN => n3900, 
                           Q => net114671, QN => n1932);
   pc_lut_reg_9_7_inst : DFFR_X1 port map( D => n7237, CK => Clk, RN => n3900, 
                           Q => net114670, QN => n1931);
   pc_lut_reg_9_5_inst : DFFR_X1 port map( D => n7236, CK => Clk, RN => n3859, 
                           Q => net114669, QN => n1930);
   pc_lut_reg_9_3_inst : DFFR_X1 port map( D => n7235, CK => Clk, RN => n3900, 
                           Q => net114668, QN => n1929);
   pc_lut_reg_9_0_inst : DFFR_X1 port map( D => n7233, CK => Clk, RN => n3900, 
                           Q => net114667, QN => n1927);
   pc_lut_reg_9_6_inst : DFFR_X1 port map( D => n7230, CK => Clk, RN => n3900, 
                           Q => net114666, QN => n1924);
   pc_lut_reg_9_8_inst : DFFR_X1 port map( D => n7229, CK => Clk, RN => n3900, 
                           Q => net114665, QN => n1923);
   pc_lut_reg_9_10_inst : DFFR_X1 port map( D => n7228, CK => Clk, RN => n3900,
                           Q => net114664, QN => n1922);
   pc_lut_reg_9_12_inst : DFFR_X1 port map( D => n7227, CK => Clk, RN => n3900,
                           Q => net114663, QN => n1921);
   pc_lut_reg_9_14_inst : DFFR_X1 port map( D => n7226, CK => Clk, RN => n3900,
                           Q => net114662, QN => n1920);
   pc_lut_reg_9_16_inst : DFFR_X1 port map( D => n7225, CK => Clk, RN => n3900,
                           Q => net114661, QN => n1919);
   pc_lut_reg_9_18_inst : DFFR_X1 port map( D => n7224, CK => Clk, RN => n3862,
                           Q => net114660, QN => n1918);
   pc_lut_reg_9_20_inst : DFFR_X1 port map( D => n7223, CK => Clk, RN => n3900,
                           Q => net114659, QN => n1917);
   pc_lut_reg_9_22_inst : DFFR_X1 port map( D => n7222, CK => Clk, RN => n3901,
                           Q => net114658, QN => n1916);
   pc_lut_reg_9_24_inst : DFFR_X1 port map( D => n7221, CK => Clk, RN => n3901,
                           Q => net114657, QN => n1915);
   pc_lut_reg_9_26_inst : DFFR_X1 port map( D => n7220, CK => Clk, RN => n3901,
                           Q => net114656, QN => n1914);
   pc_lut_reg_9_28_inst : DFFR_X1 port map( D => n7219, CK => Clk, RN => n3901,
                           Q => net114655, QN => n1913);
   pc_lut_reg_9_30_inst : DFFR_X1 port map( D => n7218, CK => Clk, RN => n3901,
                           Q => net114654, QN => n1911);
   pc_lut_reg_10_31_inst : DFFR_X1 port map( D => n7217, CK => Clk, RN => n3901
                           , Q => pc_lut_10_31_port, QN => n1909);
   pc_lut_reg_10_29_inst : DFFR_X1 port map( D => n7216, CK => Clk, RN => n3901
                           , Q => pc_lut_10_29_port, QN => n1908);
   pc_lut_reg_10_27_inst : DFFR_X1 port map( D => n7215, CK => Clk, RN => n3901
                           , Q => pc_lut_10_27_port, QN => n1907);
   pc_lut_reg_10_25_inst : DFFR_X1 port map( D => n7214, CK => Clk, RN => n3901
                           , Q => pc_lut_10_25_port, QN => n1906);
   pc_lut_reg_10_23_inst : DFFR_X1 port map( D => n7213, CK => Clk, RN => n3901
                           , Q => pc_lut_10_23_port, QN => n1905);
   pc_lut_reg_10_21_inst : DFFR_X1 port map( D => n7212, CK => Clk, RN => n3901
                           , Q => pc_lut_10_21_port, QN => n1904);
   pc_lut_reg_10_19_inst : DFFR_X1 port map( D => n7211, CK => Clk, RN => n3901
                           , Q => pc_lut_10_19_port, QN => n1903);
   pc_lut_reg_10_17_inst : DFFR_X1 port map( D => n7210, CK => Clk, RN => n3901
                           , Q => pc_lut_10_17_port, QN => n1902);
   pc_lut_reg_10_15_inst : DFFR_X1 port map( D => n7209, CK => Clk, RN => n3901
                           , Q => pc_lut_10_15_port, QN => n1901);
   pc_lut_reg_10_13_inst : DFFR_X1 port map( D => n7208, CK => Clk, RN => n3901
                           , Q => pc_lut_10_13_port, QN => n1900);
   pc_lut_reg_10_11_inst : DFFR_X1 port map( D => n7207, CK => Clk, RN => n3902
                           , Q => pc_lut_10_11_port, QN => n1899);
   pc_lut_reg_10_9_inst : DFFR_X1 port map( D => n7206, CK => Clk, RN => n3902,
                           Q => pc_lut_10_9_port, QN => n1898);
   pc_lut_reg_10_7_inst : DFFR_X1 port map( D => n7205, CK => Clk, RN => n3902,
                           Q => pc_lut_10_7_port, QN => n1897);
   pc_lut_reg_10_5_inst : DFFR_X1 port map( D => n7204, CK => Clk, RN => n3859,
                           Q => pc_lut_10_5_port, QN => n1896);
   pc_lut_reg_10_3_inst : DFFR_X1 port map( D => n7203, CK => Clk, RN => n3902,
                           Q => pc_lut_10_3_port, QN => net114653);
   pc_lut_reg_10_1_inst : DFFR_X1 port map( D => n7202, CK => Clk, RN => n3902,
                           Q => pc_lut_10_1_port, QN => net114652);
   pc_lut_reg_10_6_inst : DFFR_X1 port map( D => n7198, CK => Clk, RN => n3902,
                           Q => pc_lut_10_6_port, QN => n1893);
   pc_lut_reg_10_8_inst : DFFR_X1 port map( D => n7197, CK => Clk, RN => n3902,
                           Q => pc_lut_10_8_port, QN => n1892);
   pc_lut_reg_10_10_inst : DFFR_X1 port map( D => n7196, CK => Clk, RN => n3902
                           , Q => pc_lut_10_10_port, QN => n1891);
   pc_lut_reg_10_12_inst : DFFR_X1 port map( D => n7195, CK => Clk, RN => n3902
                           , Q => pc_lut_10_12_port, QN => n1890);
   pc_lut_reg_10_14_inst : DFFR_X1 port map( D => n7194, CK => Clk, RN => n3902
                           , Q => pc_lut_10_14_port, QN => n1889);
   pc_lut_reg_10_16_inst : DFFR_X1 port map( D => n7193, CK => Clk, RN => n3902
                           , Q => pc_lut_10_16_port, QN => n1888);
   pc_lut_reg_10_18_inst : DFFR_X1 port map( D => n7192, CK => Clk, RN => n3862
                           , Q => pc_lut_10_18_port, QN => n1887);
   pc_lut_reg_10_20_inst : DFFR_X1 port map( D => n7191, CK => Clk, RN => n3902
                           , Q => pc_lut_10_20_port, QN => n1886);
   pc_lut_reg_10_22_inst : DFFR_X1 port map( D => n7190, CK => Clk, RN => n3902
                           , Q => pc_lut_10_22_port, QN => n1885);
   pc_lut_reg_10_24_inst : DFFR_X1 port map( D => n7189, CK => Clk, RN => n3902
                           , Q => pc_lut_10_24_port, QN => n1884);
   pc_lut_reg_10_26_inst : DFFR_X1 port map( D => n7188, CK => Clk, RN => n3902
                           , Q => pc_lut_10_26_port, QN => n1883);
   pc_lut_reg_10_28_inst : DFFR_X1 port map( D => n7187, CK => Clk, RN => n3903
                           , Q => pc_lut_10_28_port, QN => n1882);
   pc_lut_reg_10_30_inst : DFFR_X1 port map( D => n7186, CK => Clk, RN => n3903
                           , Q => pc_lut_10_30_port, QN => n1880);
   pc_lut_reg_11_31_inst : DFFR_X1 port map( D => n7185, CK => Clk, RN => n3903
                           , Q => pc_lut_11_31_port, QN => n1877);
   pc_lut_reg_11_29_inst : DFFR_X1 port map( D => n7184, CK => Clk, RN => n3903
                           , Q => pc_lut_11_29_port, QN => n1876);
   pc_lut_reg_11_27_inst : DFFR_X1 port map( D => n7183, CK => Clk, RN => n3903
                           , Q => pc_lut_11_27_port, QN => n1875);
   pc_lut_reg_11_25_inst : DFFR_X1 port map( D => n7182, CK => Clk, RN => n3903
                           , Q => pc_lut_11_25_port, QN => n1874);
   pc_lut_reg_11_23_inst : DFFR_X1 port map( D => n7181, CK => Clk, RN => n3903
                           , Q => pc_lut_11_23_port, QN => n1873);
   pc_lut_reg_11_21_inst : DFFR_X1 port map( D => n7180, CK => Clk, RN => n3903
                           , Q => pc_lut_11_21_port, QN => n1872);
   pc_lut_reg_11_19_inst : DFFR_X1 port map( D => n7179, CK => Clk, RN => n3903
                           , Q => pc_lut_11_19_port, QN => n1871);
   pc_lut_reg_11_17_inst : DFFR_X1 port map( D => n7178, CK => Clk, RN => n3903
                           , Q => pc_lut_11_17_port, QN => n1870);
   pc_lut_reg_11_15_inst : DFFR_X1 port map( D => n7177, CK => Clk, RN => n3903
                           , Q => pc_lut_11_15_port, QN => n1869);
   pc_lut_reg_11_13_inst : DFFR_X1 port map( D => n7176, CK => Clk, RN => n3903
                           , Q => pc_lut_11_13_port, QN => n1868);
   pc_lut_reg_11_11_inst : DFFR_X1 port map( D => n7175, CK => Clk, RN => n3903
                           , Q => pc_lut_11_11_port, QN => n1867);
   pc_lut_reg_11_9_inst : DFFR_X1 port map( D => n7174, CK => Clk, RN => n3903,
                           Q => pc_lut_11_9_port, QN => n1866);
   pc_lut_reg_11_7_inst : DFFR_X1 port map( D => n7173, CK => Clk, RN => n3903,
                           Q => pc_lut_11_7_port, QN => n1865);
   pc_lut_reg_11_5_inst : DFFR_X1 port map( D => n7172, CK => Clk, RN => n3859,
                           Q => pc_lut_11_5_port, QN => n1864);
   pc_lut_reg_11_3_inst : DFFR_X1 port map( D => n7171, CK => Clk, RN => n3904,
                           Q => pc_lut_11_3_port, QN => net114637);
   pc_lut_reg_11_1_inst : DFFR_X1 port map( D => n7170, CK => Clk, RN => n3904,
                           Q => pc_lut_11_1_port, QN => net114636);
   pc_lut_reg_11_0_inst : DFFR_X1 port map( D => n7169, CK => Clk, RN => n3904,
                           Q => pc_lut_11_0_port, QN => net114635);
   pc_lut_reg_11_6_inst : DFFR_X1 port map( D => n7166, CK => Clk, RN => n3904,
                           Q => pc_lut_11_6_port, QN => n1860);
   pc_lut_reg_11_8_inst : DFFR_X1 port map( D => n7165, CK => Clk, RN => n3904,
                           Q => pc_lut_11_8_port, QN => n1859);
   pc_lut_reg_11_10_inst : DFFR_X1 port map( D => n7164, CK => Clk, RN => n3904
                           , Q => pc_lut_11_10_port, QN => n1858);
   pc_lut_reg_11_12_inst : DFFR_X1 port map( D => n7163, CK => Clk, RN => n3904
                           , Q => pc_lut_11_12_port, QN => n1857);
   pc_lut_reg_11_14_inst : DFFR_X1 port map( D => n7162, CK => Clk, RN => n3904
                           , Q => pc_lut_11_14_port, QN => n1856);
   pc_lut_reg_11_16_inst : DFFR_X1 port map( D => n7161, CK => Clk, RN => n3904
                           , Q => pc_lut_11_16_port, QN => n1855);
   pc_lut_reg_11_18_inst : DFFR_X1 port map( D => n7160, CK => Clk, RN => n3862
                           , Q => pc_lut_11_18_port, QN => n1854);
   pc_lut_reg_11_20_inst : DFFR_X1 port map( D => n7159, CK => Clk, RN => n3892
                           , Q => pc_lut_11_20_port, QN => n1853);
   pc_lut_reg_11_22_inst : DFFR_X1 port map( D => n7158, CK => Clk, RN => n3888
                           , Q => pc_lut_11_22_port, QN => n1852);
   pc_lut_reg_11_24_inst : DFFR_X1 port map( D => n7157, CK => Clk, RN => n3888
                           , Q => pc_lut_11_24_port, QN => n1851);
   pc_lut_reg_11_26_inst : DFFR_X1 port map( D => n7156, CK => Clk, RN => n3888
                           , Q => pc_lut_11_26_port, QN => n1850);
   pc_lut_reg_11_28_inst : DFFR_X1 port map( D => n7155, CK => Clk, RN => n3888
                           , Q => pc_lut_11_28_port, QN => n1849);
   pc_lut_reg_11_30_inst : DFFR_X1 port map( D => n7154, CK => Clk, RN => n3888
                           , Q => pc_lut_11_30_port, QN => n1847);
   pc_lut_reg_12_31_inst : DFFR_X1 port map( D => n7153, CK => Clk, RN => n3888
                           , Q => net114621, QN => n1842);
   pc_lut_reg_12_29_inst : DFFR_X1 port map( D => n7152, CK => Clk, RN => n3888
                           , Q => net114620, QN => n1841);
   pc_lut_reg_12_27_inst : DFFR_X1 port map( D => n7151, CK => Clk, RN => n3888
                           , Q => net114619, QN => n1840);
   pc_lut_reg_12_25_inst : DFFR_X1 port map( D => n7150, CK => Clk, RN => n3888
                           , Q => net114618, QN => n1839);
   pc_lut_reg_12_23_inst : DFFR_X1 port map( D => n7149, CK => Clk, RN => n3888
                           , Q => net114617, QN => n1838);
   pc_lut_reg_12_21_inst : DFFR_X1 port map( D => n7148, CK => Clk, RN => n3888
                           , Q => net114616, QN => n1837);
   pc_lut_reg_12_19_inst : DFFR_X1 port map( D => n7147, CK => Clk, RN => n3889
                           , Q => net114615, QN => n1836);
   pc_lut_reg_12_17_inst : DFFR_X1 port map( D => n7146, CK => Clk, RN => n3889
                           , Q => net114614, QN => n1835);
   pc_lut_reg_12_15_inst : DFFR_X1 port map( D => n7145, CK => Clk, RN => n3889
                           , Q => net114613, QN => n1834);
   pc_lut_reg_12_13_inst : DFFR_X1 port map( D => n7144, CK => Clk, RN => n3889
                           , Q => net114612, QN => n1833);
   pc_lut_reg_12_11_inst : DFFR_X1 port map( D => n7143, CK => Clk, RN => n3889
                           , Q => net114611, QN => n1832);
   pc_lut_reg_12_9_inst : DFFR_X1 port map( D => n7142, CK => Clk, RN => n3889,
                           Q => net114610, QN => n1831);
   pc_lut_reg_12_7_inst : DFFR_X1 port map( D => n7141, CK => Clk, RN => n3889,
                           Q => net114609, QN => n1830);
   pc_lut_reg_12_5_inst : DFFR_X1 port map( D => n7140, CK => Clk, RN => n3859,
                           Q => net114608, QN => n1829);
   pc_lut_reg_12_3_inst : DFFR_X1 port map( D => n7139, CK => Clk, RN => n3889,
                           Q => net114607, QN => n1828);
   pc_lut_reg_12_2_inst : DFFR_X1 port map( D => n7136, CK => Clk, RN => n3889,
                           Q => net114606, QN => n1825);
   pc_lut_reg_12_6_inst : DFFR_X1 port map( D => n7134, CK => Clk, RN => n3889,
                           Q => net114605, QN => n1823);
   pc_lut_reg_12_8_inst : DFFR_X1 port map( D => n7133, CK => Clk, RN => n3889,
                           Q => net114604, QN => n1822);
   pc_lut_reg_12_10_inst : DFFR_X1 port map( D => n7132, CK => Clk, RN => n3889
                           , Q => net114603, QN => n1821);
   pc_lut_reg_12_12_inst : DFFR_X1 port map( D => n7131, CK => Clk, RN => n3889
                           , Q => net114602, QN => n1820);
   pc_lut_reg_12_14_inst : DFFR_X1 port map( D => n7130, CK => Clk, RN => n3889
                           , Q => net114601, QN => n1819);
   pc_lut_reg_12_16_inst : DFFR_X1 port map( D => n7129, CK => Clk, RN => n3889
                           , Q => net114600, QN => n1818);
   pc_lut_reg_12_18_inst : DFFR_X1 port map( D => n7128, CK => Clk, RN => n3862
                           , Q => net114599, QN => n1817);
   pc_lut_reg_12_20_inst : DFFR_X1 port map( D => n7127, CK => Clk, RN => n3890
                           , Q => net114598, QN => n1816);
   pc_lut_reg_12_22_inst : DFFR_X1 port map( D => n7126, CK => Clk, RN => n3890
                           , Q => net114597, QN => n1815);
   pc_lut_reg_12_24_inst : DFFR_X1 port map( D => n7125, CK => Clk, RN => n3890
                           , Q => net114596, QN => n1814);
   pc_lut_reg_12_26_inst : DFFR_X1 port map( D => n7124, CK => Clk, RN => n3890
                           , Q => net114595, QN => n1813);
   pc_lut_reg_12_28_inst : DFFR_X1 port map( D => n7123, CK => Clk, RN => n3890
                           , Q => net114594, QN => n1812);
   pc_lut_reg_12_30_inst : DFFR_X1 port map( D => n7122, CK => Clk, RN => n3890
                           , Q => net114593, QN => n1810);
   pc_lut_reg_13_31_inst : DFFR_X1 port map( D => n7121, CK => Clk, RN => n3890
                           , Q => net114592, QN => n1808);
   pc_lut_reg_13_29_inst : DFFR_X1 port map( D => n7120, CK => Clk, RN => n3890
                           , Q => net114591, QN => n1807);
   pc_lut_reg_13_27_inst : DFFR_X1 port map( D => n7119, CK => Clk, RN => n3890
                           , Q => net114590, QN => n1806);
   pc_lut_reg_13_25_inst : DFFR_X1 port map( D => n7118, CK => Clk, RN => n3890
                           , Q => net114589, QN => n1805);
   pc_lut_reg_13_23_inst : DFFR_X1 port map( D => n7117, CK => Clk, RN => n3890
                           , Q => net114588, QN => n1804);
   pc_lut_reg_13_21_inst : DFFR_X1 port map( D => n7116, CK => Clk, RN => n3890
                           , Q => net114587, QN => n1803);
   pc_lut_reg_13_19_inst : DFFR_X1 port map( D => n7115, CK => Clk, RN => n3890
                           , Q => net114586, QN => n1802);
   pc_lut_reg_13_17_inst : DFFR_X1 port map( D => n7114, CK => Clk, RN => n3890
                           , Q => net114585, QN => n1801);
   pc_lut_reg_13_15_inst : DFFR_X1 port map( D => n7113, CK => Clk, RN => n3890
                           , Q => net114584, QN => n1800);
   pc_lut_reg_13_13_inst : DFFR_X1 port map( D => n7112, CK => Clk, RN => n3891
                           , Q => net114583, QN => n1799);
   pc_lut_reg_13_11_inst : DFFR_X1 port map( D => n7111, CK => Clk, RN => n3891
                           , Q => net114582, QN => n1798);
   pc_lut_reg_13_9_inst : DFFR_X1 port map( D => n7110, CK => Clk, RN => n3891,
                           Q => net114581, QN => n1797);
   pc_lut_reg_13_7_inst : DFFR_X1 port map( D => n7109, CK => Clk, RN => n3891,
                           Q => net114580, QN => n1796);
   pc_lut_reg_13_5_inst : DFFR_X1 port map( D => n7108, CK => Clk, RN => n3859,
                           Q => net114579, QN => n1795);
   pc_lut_reg_13_3_inst : DFFR_X1 port map( D => n7107, CK => Clk, RN => n3891,
                           Q => net114578, QN => n1794);
   pc_lut_reg_13_0_inst : DFFR_X1 port map( D => n7105, CK => Clk, RN => n3891,
                           Q => net114577, QN => n1792);
   pc_lut_reg_13_2_inst : DFFR_X1 port map( D => n7104, CK => Clk, RN => n3891,
                           Q => net114576, QN => n1791);
   pc_lut_reg_13_6_inst : DFFR_X1 port map( D => n7102, CK => Clk, RN => n3891,
                           Q => net114575, QN => n1789);
   pc_lut_reg_13_8_inst : DFFR_X1 port map( D => n7101, CK => Clk, RN => n3891,
                           Q => net114574, QN => n1788);
   pc_lut_reg_13_10_inst : DFFR_X1 port map( D => n7100, CK => Clk, RN => n3891
                           , Q => net114573, QN => n1787);
   pc_lut_reg_13_12_inst : DFFR_X1 port map( D => n7099, CK => Clk, RN => n3891
                           , Q => net114572, QN => n1786);
   pc_lut_reg_13_14_inst : DFFR_X1 port map( D => n7098, CK => Clk, RN => n3891
                           , Q => net114571, QN => n1785);
   pc_lut_reg_13_16_inst : DFFR_X1 port map( D => n7097, CK => Clk, RN => n3891
                           , Q => net114570, QN => n1784);
   pc_lut_reg_13_18_inst : DFFR_X1 port map( D => n7096, CK => Clk, RN => n3862
                           , Q => net114569, QN => n1783);
   pc_lut_reg_13_20_inst : DFFR_X1 port map( D => n7095, CK => Clk, RN => n3891
                           , Q => net114568, QN => n1782);
   pc_lut_reg_13_22_inst : DFFR_X1 port map( D => n7094, CK => Clk, RN => n3891
                           , Q => net114567, QN => n1781);
   pc_lut_reg_13_24_inst : DFFR_X1 port map( D => n7093, CK => Clk, RN => n3892
                           , Q => net114566, QN => n1780);
   pc_lut_reg_13_26_inst : DFFR_X1 port map( D => n7092, CK => Clk, RN => n3892
                           , Q => net114565, QN => n1779);
   pc_lut_reg_13_28_inst : DFFR_X1 port map( D => n7091, CK => Clk, RN => n3892
                           , Q => net114564, QN => n1778);
   pc_lut_reg_13_30_inst : DFFR_X1 port map( D => n7090, CK => Clk, RN => n3892
                           , Q => net114563, QN => n1776);
   pc_lut_reg_14_31_inst : DFFR_X1 port map( D => n7089, CK => Clk, RN => n3892
                           , Q => pc_lut_14_31_port, QN => n1774);
   pc_lut_reg_14_29_inst : DFFR_X1 port map( D => n7088, CK => Clk, RN => n3892
                           , Q => pc_lut_14_29_port, QN => n1773);
   pc_lut_reg_14_27_inst : DFFR_X1 port map( D => n7087, CK => Clk, RN => n3892
                           , Q => pc_lut_14_27_port, QN => n1772);
   pc_lut_reg_14_25_inst : DFFR_X1 port map( D => n7086, CK => Clk, RN => n3892
                           , Q => pc_lut_14_25_port, QN => n1771);
   pc_lut_reg_14_23_inst : DFFR_X1 port map( D => n7085, CK => Clk, RN => n3892
                           , Q => pc_lut_14_23_port, QN => n1770);
   pc_lut_reg_14_21_inst : DFFR_X1 port map( D => n7084, CK => Clk, RN => n3892
                           , Q => pc_lut_14_21_port, QN => n1769);
   pc_lut_reg_14_19_inst : DFFR_X1 port map( D => n7083, CK => Clk, RN => n3892
                           , Q => pc_lut_14_19_port, QN => n1768);
   pc_lut_reg_14_17_inst : DFFR_X1 port map( D => n7082, CK => Clk, RN => n3892
                           , Q => pc_lut_14_17_port, QN => n1767);
   pc_lut_reg_14_15_inst : DFFR_X1 port map( D => n7081, CK => Clk, RN => n3892
                           , Q => pc_lut_14_15_port, QN => n1766);
   pc_lut_reg_14_13_inst : DFFR_X1 port map( D => n7080, CK => Clk, RN => n3892
                           , Q => pc_lut_14_13_port, QN => n1765);
   pc_lut_reg_14_11_inst : DFFR_X1 port map( D => n7079, CK => Clk, RN => n3893
                           , Q => pc_lut_14_11_port, QN => n1764);
   pc_lut_reg_14_9_inst : DFFR_X1 port map( D => n7078, CK => Clk, RN => n3893,
                           Q => pc_lut_14_9_port, QN => n1763);
   pc_lut_reg_14_7_inst : DFFR_X1 port map( D => n7077, CK => Clk, RN => n3893,
                           Q => pc_lut_14_7_port, QN => n1762);
   pc_lut_reg_14_5_inst : DFFR_X1 port map( D => n7076, CK => Clk, RN => n3859,
                           Q => pc_lut_14_5_port, QN => n1761);
   pc_lut_reg_14_6_inst : DFFR_X1 port map( D => n7070, CK => Clk, RN => n3893,
                           Q => pc_lut_14_6_port, QN => n1757);
   pc_lut_reg_14_8_inst : DFFR_X1 port map( D => n7069, CK => Clk, RN => n3893,
                           Q => pc_lut_14_8_port, QN => n1756);
   pc_lut_reg_14_10_inst : DFFR_X1 port map( D => n7068, CK => Clk, RN => n3893
                           , Q => pc_lut_14_10_port, QN => n1755);
   pc_lut_reg_14_12_inst : DFFR_X1 port map( D => n7067, CK => Clk, RN => n3893
                           , Q => pc_lut_14_12_port, QN => n1754);
   pc_lut_reg_14_14_inst : DFFR_X1 port map( D => n7066, CK => Clk, RN => n3893
                           , Q => pc_lut_14_14_port, QN => n1753);
   pc_lut_reg_14_16_inst : DFFR_X1 port map( D => n7065, CK => Clk, RN => n3893
                           , Q => pc_lut_14_16_port, QN => n1752);
   pc_lut_reg_14_18_inst : DFFR_X1 port map( D => n7064, CK => Clk, RN => n3862
                           , Q => pc_lut_14_18_port, QN => n1751);
   pc_lut_reg_14_20_inst : DFFR_X1 port map( D => n7063, CK => Clk, RN => n3893
                           , Q => pc_lut_14_20_port, QN => n1750);
   pc_lut_reg_14_22_inst : DFFR_X1 port map( D => n7062, CK => Clk, RN => n3893
                           , Q => pc_lut_14_22_port, QN => n1749);
   pc_lut_reg_14_24_inst : DFFR_X1 port map( D => n7061, CK => Clk, RN => n3893
                           , Q => pc_lut_14_24_port, QN => n1748);
   pc_lut_reg_14_26_inst : DFFR_X1 port map( D => n7060, CK => Clk, RN => n3893
                           , Q => pc_lut_14_26_port, QN => n1747);
   pc_lut_reg_14_28_inst : DFFR_X1 port map( D => n7059, CK => Clk, RN => n3893
                           , Q => pc_lut_14_28_port, QN => n1746);
   pc_lut_reg_14_30_inst : DFFR_X1 port map( D => n7058, CK => Clk, RN => n3893
                           , Q => pc_lut_14_30_port, QN => n1744);
   pc_lut_reg_15_31_inst : DFFR_X1 port map( D => n7057, CK => Clk, RN => n3894
                           , Q => pc_lut_15_31_port, QN => n1741);
   pc_lut_reg_15_29_inst : DFFR_X1 port map( D => n7056, CK => Clk, RN => n3894
                           , Q => pc_lut_15_29_port, QN => n1740);
   pc_lut_reg_15_27_inst : DFFR_X1 port map( D => n7055, CK => Clk, RN => n3894
                           , Q => pc_lut_15_27_port, QN => n1739);
   pc_lut_reg_15_25_inst : DFFR_X1 port map( D => n7054, CK => Clk, RN => n3894
                           , Q => pc_lut_15_25_port, QN => n1738);
   pc_lut_reg_15_23_inst : DFFR_X1 port map( D => n7053, CK => Clk, RN => n3894
                           , Q => pc_lut_15_23_port, QN => n1737);
   pc_lut_reg_15_21_inst : DFFR_X1 port map( D => n7052, CK => Clk, RN => n3894
                           , Q => pc_lut_15_21_port, QN => n1736);
   pc_lut_reg_15_19_inst : DFFR_X1 port map( D => n7051, CK => Clk, RN => n3894
                           , Q => pc_lut_15_19_port, QN => n1735);
   pc_lut_reg_15_17_inst : DFFR_X1 port map( D => n7050, CK => Clk, RN => n3894
                           , Q => pc_lut_15_17_port, QN => n1734);
   pc_lut_reg_15_15_inst : DFFR_X1 port map( D => n7049, CK => Clk, RN => n3894
                           , Q => pc_lut_15_15_port, QN => n1733);
   pc_lut_reg_15_13_inst : DFFR_X1 port map( D => n7048, CK => Clk, RN => n3894
                           , Q => pc_lut_15_13_port, QN => n1732);
   pc_lut_reg_15_11_inst : DFFR_X1 port map( D => n7047, CK => Clk, RN => n3894
                           , Q => pc_lut_15_11_port, QN => n1731);
   pc_lut_reg_15_9_inst : DFFR_X1 port map( D => n7046, CK => Clk, RN => n3894,
                           Q => pc_lut_15_9_port, QN => n1730);
   pc_lut_reg_15_7_inst : DFFR_X1 port map( D => n7045, CK => Clk, RN => n3894,
                           Q => pc_lut_15_7_port, QN => n1729);
   pc_lut_reg_15_5_inst : DFFR_X1 port map( D => n7044, CK => Clk, RN => n3859,
                           Q => pc_lut_15_5_port, QN => n1728);
   pc_lut_reg_15_6_inst : DFFR_X1 port map( D => n7038, CK => Clk, RN => n3947,
                           Q => pc_lut_15_6_port, QN => n1723);
   pc_lut_reg_15_8_inst : DFFR_X1 port map( D => n7037, CK => Clk, RN => n3947,
                           Q => pc_lut_15_8_port, QN => n1722);
   pc_lut_reg_15_10_inst : DFFR_X1 port map( D => n7036, CK => Clk, RN => n3947
                           , Q => pc_lut_15_10_port, QN => n1721);
   pc_lut_reg_15_12_inst : DFFR_X1 port map( D => n7035, CK => Clk, RN => n3947
                           , Q => pc_lut_15_12_port, QN => n1720);
   pc_lut_reg_15_14_inst : DFFR_X1 port map( D => n7034, CK => Clk, RN => n3947
                           , Q => pc_lut_15_14_port, QN => n1719);
   pc_lut_reg_15_16_inst : DFFR_X1 port map( D => n7033, CK => Clk, RN => n3948
                           , Q => pc_lut_15_16_port, QN => n1718);
   pc_lut_reg_15_18_inst : DFFR_X1 port map( D => n7032, CK => Clk, RN => n3863
                           , Q => pc_lut_15_18_port, QN => n1717);
   pc_lut_reg_15_20_inst : DFFR_X1 port map( D => n7031, CK => Clk, RN => n3948
                           , Q => pc_lut_15_20_port, QN => n1716);
   pc_lut_reg_15_22_inst : DFFR_X1 port map( D => n7030, CK => Clk, RN => n3948
                           , Q => pc_lut_15_22_port, QN => n1715);
   pc_lut_reg_15_24_inst : DFFR_X1 port map( D => n7029, CK => Clk, RN => n3948
                           , Q => pc_lut_15_24_port, QN => n1714);
   pc_lut_reg_15_26_inst : DFFR_X1 port map( D => n7028, CK => Clk, RN => n3948
                           , Q => pc_lut_15_26_port, QN => n1713);
   pc_lut_reg_15_28_inst : DFFR_X1 port map( D => n7027, CK => Clk, RN => n3948
                           , Q => pc_lut_15_28_port, QN => n1712);
   pc_lut_reg_15_30_inst : DFFR_X1 port map( D => n7026, CK => Clk, RN => n3949
                           , Q => pc_lut_15_30_port, QN => n1710);
   pc_lut_reg_16_31_inst : DFFR_X1 port map( D => n7025, CK => Clk, RN => n3948
                           , Q => net114508, QN => n1707);
   pc_lut_reg_16_29_inst : DFFR_X1 port map( D => n7024, CK => Clk, RN => n3948
                           , Q => net114507, QN => n1706);
   pc_lut_reg_16_27_inst : DFFR_X1 port map( D => n7023, CK => Clk, RN => n3948
                           , Q => net114506, QN => n1705);
   pc_lut_reg_16_25_inst : DFFR_X1 port map( D => n7022, CK => Clk, RN => n3948
                           , Q => net114505, QN => n1704);
   pc_lut_reg_16_23_inst : DFFR_X1 port map( D => n7021, CK => Clk, RN => n3948
                           , Q => net114504, QN => n1703);
   pc_lut_reg_16_21_inst : DFFR_X1 port map( D => n7020, CK => Clk, RN => n3948
                           , Q => net114503, QN => n1702);
   pc_lut_reg_16_19_inst : DFFR_X1 port map( D => n7019, CK => Clk, RN => n3948
                           , Q => net114502, QN => n1701);
   pc_lut_reg_16_17_inst : DFFR_X1 port map( D => n7018, CK => Clk, RN => n3948
                           , Q => net114501, QN => n1700);
   pc_lut_reg_16_15_inst : DFFR_X1 port map( D => n7017, CK => Clk, RN => n3948
                           , Q => net114500, QN => n1699);
   pc_lut_reg_16_13_inst : DFFR_X1 port map( D => n7016, CK => Clk, RN => n3949
                           , Q => net114499, QN => n1698);
   pc_lut_reg_16_11_inst : DFFR_X1 port map( D => n7015, CK => Clk, RN => n3949
                           , Q => net114498, QN => n1697);
   pc_lut_reg_16_9_inst : DFFR_X1 port map( D => n7014, CK => Clk, RN => n3949,
                           Q => net114497, QN => n1696);
   pc_lut_reg_16_7_inst : DFFR_X1 port map( D => n7013, CK => Clk, RN => n3949,
                           Q => net114496, QN => n1695);
   pc_lut_reg_16_5_inst : DFFR_X1 port map( D => n7012, CK => Clk, RN => n3859,
                           Q => net114495, QN => n1694);
   pc_lut_reg_16_4_inst : DFFR_X1 port map( D => n7007, CK => Clk, RN => n3949,
                           Q => net114494, QN => n1689);
   pc_lut_reg_16_6_inst : DFFR_X1 port map( D => n7006, CK => Clk, RN => n3949,
                           Q => net114493, QN => n1688);
   pc_lut_reg_16_8_inst : DFFR_X1 port map( D => n7005, CK => Clk, RN => n3949,
                           Q => net114492, QN => n1687);
   pc_lut_reg_16_10_inst : DFFR_X1 port map( D => n7004, CK => Clk, RN => n3949
                           , Q => net114491, QN => n1686);
   pc_lut_reg_16_12_inst : DFFR_X1 port map( D => n7003, CK => Clk, RN => n3949
                           , Q => net114490, QN => n1685);
   pc_lut_reg_16_14_inst : DFFR_X1 port map( D => n7002, CK => Clk, RN => n3949
                           , Q => net114489, QN => n1684);
   pc_lut_reg_16_16_inst : DFFR_X1 port map( D => n7001, CK => Clk, RN => n3949
                           , Q => net114488, QN => n1683);
   pc_lut_reg_16_18_inst : DFFR_X1 port map( D => n7000, CK => Clk, RN => n3862
                           , Q => net114487, QN => n1682);
   pc_lut_reg_16_20_inst : DFFR_X1 port map( D => n6999, CK => Clk, RN => n3949
                           , Q => net114486, QN => n1681);
   pc_lut_reg_16_22_inst : DFFR_X1 port map( D => n6998, CK => Clk, RN => n3950
                           , Q => net114485, QN => n1680);
   pc_lut_reg_16_24_inst : DFFR_X1 port map( D => n6997, CK => Clk, RN => n3950
                           , Q => net114484, QN => n1679);
   pc_lut_reg_16_26_inst : DFFR_X1 port map( D => n6996, CK => Clk, RN => n3950
                           , Q => net114483, QN => n1678);
   pc_lut_reg_16_28_inst : DFFR_X1 port map( D => n6995, CK => Clk, RN => n3950
                           , Q => net114482, QN => n1677);
   pc_lut_reg_16_30_inst : DFFR_X1 port map( D => n6994, CK => Clk, RN => n3950
                           , Q => net114481, QN => n1675);
   pc_lut_reg_17_31_inst : DFFR_X1 port map( D => n6993, CK => Clk, RN => n3950
                           , Q => net114480, QN => n1673);
   pc_lut_reg_17_29_inst : DFFR_X1 port map( D => n6992, CK => Clk, RN => n3950
                           , Q => net114479, QN => n1672);
   pc_lut_reg_17_27_inst : DFFR_X1 port map( D => n6991, CK => Clk, RN => n3950
                           , Q => net114478, QN => n1671);
   pc_lut_reg_17_25_inst : DFFR_X1 port map( D => n6990, CK => Clk, RN => n3950
                           , Q => net114477, QN => n1670);
   pc_lut_reg_17_23_inst : DFFR_X1 port map( D => n6989, CK => Clk, RN => n3950
                           , Q => net114476, QN => n1669);
   pc_lut_reg_17_21_inst : DFFR_X1 port map( D => n6988, CK => Clk, RN => n3950
                           , Q => net114475, QN => n1668);
   pc_lut_reg_17_19_inst : DFFR_X1 port map( D => n6987, CK => Clk, RN => n3950
                           , Q => net114474, QN => n1667);
   pc_lut_reg_17_17_inst : DFFR_X1 port map( D => n6986, CK => Clk, RN => n3950
                           , Q => net114473, QN => n1666);
   pc_lut_reg_17_15_inst : DFFR_X1 port map( D => n6985, CK => Clk, RN => n3950
                           , Q => net114472, QN => n1665);
   pc_lut_reg_17_13_inst : DFFR_X1 port map( D => n6984, CK => Clk, RN => n3951
                           , Q => net114471, QN => n1664);
   pc_lut_reg_17_11_inst : DFFR_X1 port map( D => n6983, CK => Clk, RN => n3951
                           , Q => net114470, QN => n1663);
   pc_lut_reg_17_9_inst : DFFR_X1 port map( D => n6982, CK => Clk, RN => n3951,
                           Q => net114469, QN => n1662);
   pc_lut_reg_17_7_inst : DFFR_X1 port map( D => n6981, CK => Clk, RN => n3950,
                           Q => net114468, QN => n1661);
   pc_lut_reg_17_5_inst : DFFR_X1 port map( D => n6980, CK => Clk, RN => n3859,
                           Q => net114467, QN => n1660);
   pc_lut_reg_17_0_inst : DFFR_X1 port map( D => n6977, CK => Clk, RN => n3951,
                           Q => net114466, QN => n1657);
   pc_lut_reg_17_4_inst : DFFR_X1 port map( D => n6975, CK => Clk, RN => n3951,
                           Q => net114465, QN => n1655);
   pc_lut_reg_17_6_inst : DFFR_X1 port map( D => n6974, CK => Clk, RN => n3951,
                           Q => net114464, QN => n1654);
   pc_lut_reg_17_8_inst : DFFR_X1 port map( D => n6973, CK => Clk, RN => n3951,
                           Q => net114463, QN => n1653);
   pc_lut_reg_17_10_inst : DFFR_X1 port map( D => n6972, CK => Clk, RN => n3951
                           , Q => net114462, QN => n1652);
   pc_lut_reg_17_12_inst : DFFR_X1 port map( D => n6971, CK => Clk, RN => n3951
                           , Q => net114461, QN => n1651);
   pc_lut_reg_17_14_inst : DFFR_X1 port map( D => n6970, CK => Clk, RN => n3949
                           , Q => net114460, QN => n1650);
   pc_lut_reg_17_16_inst : DFFR_X1 port map( D => n6969, CK => Clk, RN => n3951
                           , Q => net114459, QN => n1649);
   pc_lut_reg_17_18_inst : DFFR_X1 port map( D => n6968, CK => Clk, RN => n3862
                           , Q => net114458, QN => n1648);
   pc_lut_reg_17_20_inst : DFFR_X1 port map( D => n6967, CK => Clk, RN => n3952
                           , Q => net114457, QN => n1647);
   pc_lut_reg_17_22_inst : DFFR_X1 port map( D => n6966, CK => Clk, RN => n3952
                           , Q => net114456, QN => n1646);
   pc_lut_reg_17_24_inst : DFFR_X1 port map( D => n6965, CK => Clk, RN => n3951
                           , Q => net114455, QN => n1645);
   pc_lut_reg_17_26_inst : DFFR_X1 port map( D => n6964, CK => Clk, RN => n3952
                           , Q => net114454, QN => n1644);
   pc_lut_reg_17_28_inst : DFFR_X1 port map( D => n6963, CK => Clk, RN => n3951
                           , Q => net114453, QN => n1643);
   pc_lut_reg_17_30_inst : DFFR_X1 port map( D => n6962, CK => Clk, RN => n3952
                           , Q => net114452, QN => n1641);
   pc_lut_reg_18_31_inst : DFFR_X1 port map( D => n6961, CK => Clk, RN => n3951
                           , Q => pc_lut_18_31_port, QN => n1639);
   pc_lut_reg_18_29_inst : DFFR_X1 port map( D => n6960, CK => Clk, RN => n3951
                           , Q => pc_lut_18_29_port, QN => n1638);
   pc_lut_reg_18_27_inst : DFFR_X1 port map( D => n6959, CK => Clk, RN => n3952
                           , Q => pc_lut_18_27_port, QN => n1637);
   pc_lut_reg_18_25_inst : DFFR_X1 port map( D => n6958, CK => Clk, RN => n3952
                           , Q => pc_lut_18_25_port, QN => n1636);
   pc_lut_reg_18_23_inst : DFFR_X1 port map( D => n6957, CK => Clk, RN => n3952
                           , Q => pc_lut_18_23_port, QN => n1635);
   pc_lut_reg_18_21_inst : DFFR_X1 port map( D => n6956, CK => Clk, RN => n3952
                           , Q => pc_lut_18_21_port, QN => n1634);
   pc_lut_reg_18_19_inst : DFFR_X1 port map( D => n6955, CK => Clk, RN => n3953
                           , Q => pc_lut_18_19_port, QN => n1633);
   pc_lut_reg_18_17_inst : DFFR_X1 port map( D => n6954, CK => Clk, RN => n3952
                           , Q => pc_lut_18_17_port, QN => n1632);
   pc_lut_reg_18_15_inst : DFFR_X1 port map( D => n6953, CK => Clk, RN => n3953
                           , Q => pc_lut_18_15_port, QN => n1631);
   pc_lut_reg_18_13_inst : DFFR_X1 port map( D => n6952, CK => Clk, RN => n3952
                           , Q => pc_lut_18_13_port, QN => n1630);
   pc_lut_reg_18_11_inst : DFFR_X1 port map( D => n6951, CK => Clk, RN => n3953
                           , Q => pc_lut_18_11_port, QN => n1629);
   pc_lut_reg_18_9_inst : DFFR_X1 port map( D => n6950, CK => Clk, RN => n3952,
                           Q => pc_lut_18_9_port, QN => n1628);
   pc_lut_reg_18_7_inst : DFFR_X1 port map( D => n6949, CK => Clk, RN => n3951,
                           Q => pc_lut_18_7_port, QN => n1627);
   pc_lut_reg_18_5_inst : DFFR_X1 port map( D => n6948, CK => Clk, RN => n3860,
                           Q => pc_lut_18_5_port, QN => n1626);
   pc_lut_reg_18_1_inst : DFFR_X1 port map( D => n6946, CK => Clk, RN => n3952,
                           Q => pc_lut_18_1_port, QN => net114451);
   pc_lut_reg_18_4_inst : DFFR_X1 port map( D => n6943, CK => Clk, RN => n3952,
                           Q => pc_lut_18_4_port, QN => net114450);
   pc_lut_reg_18_6_inst : DFFR_X1 port map( D => n6942, CK => Clk, RN => n3952,
                           Q => pc_lut_18_6_port, QN => n1623);
   pc_lut_reg_18_8_inst : DFFR_X1 port map( D => n6941, CK => Clk, RN => n3952,
                           Q => pc_lut_18_8_port, QN => n1622);
   pc_lut_reg_18_10_inst : DFFR_X1 port map( D => n6940, CK => Clk, RN => n3941
                           , Q => pc_lut_18_10_port, QN => n1621);
   pc_lut_reg_18_12_inst : DFFR_X1 port map( D => n6939, CK => Clk, RN => n3937
                           , Q => pc_lut_18_12_port, QN => n1620);
   pc_lut_reg_18_14_inst : DFFR_X1 port map( D => n6938, CK => Clk, RN => n3937
                           , Q => pc_lut_18_14_port, QN => n1619);
   pc_lut_reg_18_16_inst : DFFR_X1 port map( D => n6937, CK => Clk, RN => n3937
                           , Q => pc_lut_18_16_port, QN => n1618);
   pc_lut_reg_18_18_inst : DFFR_X1 port map( D => n6936, CK => Clk, RN => n3862
                           , Q => pc_lut_18_18_port, QN => n1617);
   pc_lut_reg_18_20_inst : DFFR_X1 port map( D => n6935, CK => Clk, RN => n3937
                           , Q => pc_lut_18_20_port, QN => n1616);
   pc_lut_reg_18_22_inst : DFFR_X1 port map( D => n6934, CK => Clk, RN => n3937
                           , Q => pc_lut_18_22_port, QN => n1615);
   pc_lut_reg_18_24_inst : DFFR_X1 port map( D => n6933, CK => Clk, RN => n3937
                           , Q => pc_lut_18_24_port, QN => n1614);
   pc_lut_reg_18_26_inst : DFFR_X1 port map( D => n6932, CK => Clk, RN => n3938
                           , Q => pc_lut_18_26_port, QN => n1613);
   pc_lut_reg_18_28_inst : DFFR_X1 port map( D => n6931, CK => Clk, RN => n3937
                           , Q => pc_lut_18_28_port, QN => n1612);
   pc_lut_reg_18_30_inst : DFFR_X1 port map( D => n6930, CK => Clk, RN => n3938
                           , Q => pc_lut_18_30_port, QN => n1610);
   pc_lut_reg_19_31_inst : DFFR_X1 port map( D => n6929, CK => Clk, RN => n3937
                           , Q => pc_lut_19_31_port, QN => n1607);
   pc_lut_reg_19_29_inst : DFFR_X1 port map( D => n6928, CK => Clk, RN => n3937
                           , Q => pc_lut_19_29_port, QN => n1606);
   pc_lut_reg_19_27_inst : DFFR_X1 port map( D => n6927, CK => Clk, RN => n3937
                           , Q => pc_lut_19_27_port, QN => n1605);
   pc_lut_reg_19_25_inst : DFFR_X1 port map( D => n6926, CK => Clk, RN => n3938
                           , Q => pc_lut_19_25_port, QN => n1604);
   pc_lut_reg_19_23_inst : DFFR_X1 port map( D => n6925, CK => Clk, RN => n3938
                           , Q => pc_lut_19_23_port, QN => n1603);
   pc_lut_reg_19_21_inst : DFFR_X1 port map( D => n6924, CK => Clk, RN => n3938
                           , Q => pc_lut_19_21_port, QN => n1602);
   pc_lut_reg_19_19_inst : DFFR_X1 port map( D => n6923, CK => Clk, RN => n3938
                           , Q => pc_lut_19_19_port, QN => n1601);
   pc_lut_reg_19_17_inst : DFFR_X1 port map( D => n6922, CK => Clk, RN => n3938
                           , Q => pc_lut_19_17_port, QN => n1600);
   pc_lut_reg_19_15_inst : DFFR_X1 port map( D => n6921, CK => Clk, RN => n3938
                           , Q => pc_lut_19_15_port, QN => n1599);
   pc_lut_reg_19_13_inst : DFFR_X1 port map( D => n6920, CK => Clk, RN => n3938
                           , Q => pc_lut_19_13_port, QN => n1598);
   pc_lut_reg_19_11_inst : DFFR_X1 port map( D => n6919, CK => Clk, RN => n3938
                           , Q => pc_lut_19_11_port, QN => n1597);
   pc_lut_reg_19_9_inst : DFFR_X1 port map( D => n6918, CK => Clk, RN => n3938,
                           Q => pc_lut_19_9_port, QN => n1596);
   pc_lut_reg_19_7_inst : DFFR_X1 port map( D => n6917, CK => Clk, RN => n3938,
                           Q => pc_lut_19_7_port, QN => n1595);
   pc_lut_reg_19_5_inst : DFFR_X1 port map( D => n6916, CK => Clk, RN => n3860,
                           Q => pc_lut_19_5_port, QN => n1594);
   pc_lut_reg_19_1_inst : DFFR_X1 port map( D => n6914, CK => Clk, RN => n3938,
                           Q => pc_lut_19_1_port, QN => net114435);
   pc_lut_reg_19_0_inst : DFFR_X1 port map( D => n6913, CK => Clk, RN => n3938,
                           Q => pc_lut_19_0_port, QN => net114434);
   pc_lut_reg_19_4_inst : DFFR_X1 port map( D => n6911, CK => Clk, RN => n3938,
                           Q => pc_lut_19_4_port, QN => net114433);
   pc_lut_reg_19_6_inst : DFFR_X1 port map( D => n6910, CK => Clk, RN => n3939,
                           Q => pc_lut_19_6_port, QN => n1590);
   pc_lut_reg_19_8_inst : DFFR_X1 port map( D => n6909, CK => Clk, RN => n3939,
                           Q => pc_lut_19_8_port, QN => n1589);
   pc_lut_reg_19_10_inst : DFFR_X1 port map( D => n6908, CK => Clk, RN => n3939
                           , Q => pc_lut_19_10_port, QN => n1588);
   pc_lut_reg_19_12_inst : DFFR_X1 port map( D => n6907, CK => Clk, RN => n3939
                           , Q => pc_lut_19_12_port, QN => n1587);
   pc_lut_reg_19_14_inst : DFFR_X1 port map( D => n6906, CK => Clk, RN => n3939
                           , Q => pc_lut_19_14_port, QN => n1586);
   pc_lut_reg_19_16_inst : DFFR_X1 port map( D => n6905, CK => Clk, RN => n3939
                           , Q => pc_lut_19_16_port, QN => n1585);
   pc_lut_reg_19_18_inst : DFFR_X1 port map( D => n6904, CK => Clk, RN => n3862
                           , Q => pc_lut_19_18_port, QN => n1584);
   pc_lut_reg_19_20_inst : DFFR_X1 port map( D => n6903, CK => Clk, RN => n3939
                           , Q => pc_lut_19_20_port, QN => n1583);
   pc_lut_reg_19_22_inst : DFFR_X1 port map( D => n6902, CK => Clk, RN => n3939
                           , Q => pc_lut_19_22_port, QN => n1582);
   pc_lut_reg_19_24_inst : DFFR_X1 port map( D => n6901, CK => Clk, RN => n3939
                           , Q => pc_lut_19_24_port, QN => n1581);
   pc_lut_reg_19_26_inst : DFFR_X1 port map( D => n6900, CK => Clk, RN => n3939
                           , Q => pc_lut_19_26_port, QN => n1580);
   pc_lut_reg_19_28_inst : DFFR_X1 port map( D => n6899, CK => Clk, RN => n3939
                           , Q => pc_lut_19_28_port, QN => n1579);
   pc_lut_reg_19_30_inst : DFFR_X1 port map( D => n6898, CK => Clk, RN => n3939
                           , Q => pc_lut_19_30_port, QN => n1577);
   pc_lut_reg_20_31_inst : DFFR_X1 port map( D => n6897, CK => Clk, RN => n3939
                           , Q => pc_lut_20_31_port, QN => n1575);
   pc_lut_reg_20_29_inst : DFFR_X1 port map( D => n6896, CK => Clk, RN => n3939
                           , Q => pc_lut_20_29_port, QN => n1574);
   pc_lut_reg_20_27_inst : DFFR_X1 port map( D => n6895, CK => Clk, RN => n3939
                           , Q => pc_lut_20_27_port, QN => n1573);
   pc_lut_reg_20_25_inst : DFFR_X1 port map( D => n6894, CK => Clk, RN => n3940
                           , Q => pc_lut_20_25_port, QN => n1572);
   pc_lut_reg_20_23_inst : DFFR_X1 port map( D => n6893, CK => Clk, RN => n3940
                           , Q => pc_lut_20_23_port, QN => n1571);
   pc_lut_reg_20_21_inst : DFFR_X1 port map( D => n6892, CK => Clk, RN => n3940
                           , Q => pc_lut_20_21_port, QN => n1570);
   pc_lut_reg_20_19_inst : DFFR_X1 port map( D => n6891, CK => Clk, RN => n3940
                           , Q => pc_lut_20_19_port, QN => n1569);
   pc_lut_reg_20_17_inst : DFFR_X1 port map( D => n6890, CK => Clk, RN => n3940
                           , Q => pc_lut_20_17_port, QN => n1568);
   pc_lut_reg_20_15_inst : DFFR_X1 port map( D => n6889, CK => Clk, RN => n3940
                           , Q => pc_lut_20_15_port, QN => n1567);
   pc_lut_reg_20_13_inst : DFFR_X1 port map( D => n6888, CK => Clk, RN => n3940
                           , Q => pc_lut_20_13_port, QN => n1566);
   pc_lut_reg_20_11_inst : DFFR_X1 port map( D => n6887, CK => Clk, RN => n3940
                           , Q => pc_lut_20_11_port, QN => n1565);
   pc_lut_reg_20_9_inst : DFFR_X1 port map( D => n6886, CK => Clk, RN => n3940,
                           Q => pc_lut_20_9_port, QN => n1564);
   pc_lut_reg_20_7_inst : DFFR_X1 port map( D => n6885, CK => Clk, RN => n3940,
                           Q => pc_lut_20_7_port, QN => n1563);
   pc_lut_reg_20_5_inst : DFFR_X1 port map( D => n6884, CK => Clk, RN => n3860,
                           Q => pc_lut_20_5_port, QN => n1562);
   pc_lut_reg_20_2_inst : DFFR_X1 port map( D => n6880, CK => Clk, RN => n3940,
                           Q => pc_lut_20_2_port, QN => net114419);
   pc_lut_reg_20_4_inst : DFFR_X1 port map( D => n6879, CK => Clk, RN => n3940,
                           Q => pc_lut_20_4_port, QN => net114418);
   pc_lut_reg_20_6_inst : DFFR_X1 port map( D => n6878, CK => Clk, RN => n3940,
                           Q => pc_lut_20_6_port, QN => n1559);
   pc_lut_reg_20_8_inst : DFFR_X1 port map( D => n6877, CK => Clk, RN => n3940,
                           Q => pc_lut_20_8_port, QN => n1558);
   pc_lut_reg_20_10_inst : DFFR_X1 port map( D => n6876, CK => Clk, RN => n3940
                           , Q => pc_lut_20_10_port, QN => n1557);
   pc_lut_reg_20_12_inst : DFFR_X1 port map( D => n6875, CK => Clk, RN => n3941
                           , Q => pc_lut_20_12_port, QN => n1556);
   pc_lut_reg_20_14_inst : DFFR_X1 port map( D => n6874, CK => Clk, RN => n3941
                           , Q => pc_lut_20_14_port, QN => n1555);
   pc_lut_reg_20_16_inst : DFFR_X1 port map( D => n6873, CK => Clk, RN => n3941
                           , Q => pc_lut_20_16_port, QN => n1554);
   pc_lut_reg_20_18_inst : DFFR_X1 port map( D => n6872, CK => Clk, RN => n3863
                           , Q => pc_lut_20_18_port, QN => n1553);
   pc_lut_reg_20_20_inst : DFFR_X1 port map( D => n6871, CK => Clk, RN => n3941
                           , Q => pc_lut_20_20_port, QN => n1552);
   pc_lut_reg_20_22_inst : DFFR_X1 port map( D => n6870, CK => Clk, RN => n3941
                           , Q => pc_lut_20_22_port, QN => n1551);
   pc_lut_reg_20_24_inst : DFFR_X1 port map( D => n6869, CK => Clk, RN => n3941
                           , Q => pc_lut_20_24_port, QN => n1550);
   pc_lut_reg_20_26_inst : DFFR_X1 port map( D => n6868, CK => Clk, RN => n3941
                           , Q => pc_lut_20_26_port, QN => n1549);
   pc_lut_reg_20_28_inst : DFFR_X1 port map( D => n6867, CK => Clk, RN => n3941
                           , Q => pc_lut_20_28_port, QN => n1548);
   pc_lut_reg_20_30_inst : DFFR_X1 port map( D => n6866, CK => Clk, RN => n3941
                           , Q => pc_lut_20_30_port, QN => n1546);
   pc_lut_reg_21_31_inst : DFFR_X1 port map( D => n6865, CK => Clk, RN => n3941
                           , Q => pc_lut_21_31_port, QN => n1544);
   pc_lut_reg_21_29_inst : DFFR_X1 port map( D => n6864, CK => Clk, RN => n3941
                           , Q => pc_lut_21_29_port, QN => n1543);
   pc_lut_reg_21_27_inst : DFFR_X1 port map( D => n6863, CK => Clk, RN => n3941
                           , Q => pc_lut_21_27_port, QN => n1542);
   pc_lut_reg_21_25_inst : DFFR_X1 port map( D => n6862, CK => Clk, RN => n3941
                           , Q => pc_lut_21_25_port, QN => n1541);
   pc_lut_reg_21_23_inst : DFFR_X1 port map( D => n6861, CK => Clk, RN => n3941
                           , Q => pc_lut_21_23_port, QN => n1540);
   pc_lut_reg_21_21_inst : DFFR_X1 port map( D => n6860, CK => Clk, RN => n3942
                           , Q => pc_lut_21_21_port, QN => n1539);
   pc_lut_reg_21_19_inst : DFFR_X1 port map( D => n6859, CK => Clk, RN => n3942
                           , Q => pc_lut_21_19_port, QN => n1538);
   pc_lut_reg_21_17_inst : DFFR_X1 port map( D => n6858, CK => Clk, RN => n3942
                           , Q => pc_lut_21_17_port, QN => n1537);
   pc_lut_reg_21_15_inst : DFFR_X1 port map( D => n6857, CK => Clk, RN => n3942
                           , Q => pc_lut_21_15_port, QN => n1536);
   pc_lut_reg_21_13_inst : DFFR_X1 port map( D => n6856, CK => Clk, RN => n3942
                           , Q => pc_lut_21_13_port, QN => n1535);
   pc_lut_reg_21_11_inst : DFFR_X1 port map( D => n6855, CK => Clk, RN => n3942
                           , Q => pc_lut_21_11_port, QN => n1534);
   pc_lut_reg_21_9_inst : DFFR_X1 port map( D => n6854, CK => Clk, RN => n3942,
                           Q => pc_lut_21_9_port, QN => n1533);
   pc_lut_reg_21_7_inst : DFFR_X1 port map( D => n6853, CK => Clk, RN => n3942,
                           Q => pc_lut_21_7_port, QN => n1532);
   pc_lut_reg_21_5_inst : DFFR_X1 port map( D => n6852, CK => Clk, RN => n3860,
                           Q => pc_lut_21_5_port, QN => n1531);
   pc_lut_reg_21_0_inst : DFFR_X1 port map( D => n6849, CK => Clk, RN => n3942,
                           Q => pc_lut_21_0_port, QN => net114417);
   pc_lut_reg_21_2_inst : DFFR_X1 port map( D => n6848, CK => Clk, RN => n3942,
                           Q => pc_lut_21_2_port, QN => net114416);
   pc_lut_reg_21_4_inst : DFFR_X1 port map( D => n6847, CK => Clk, RN => n3942,
                           Q => pc_lut_21_4_port, QN => net114415);
   pc_lut_reg_21_6_inst : DFFR_X1 port map( D => n6846, CK => Clk, RN => n3942,
                           Q => pc_lut_21_6_port, QN => n1527);
   pc_lut_reg_21_8_inst : DFFR_X1 port map( D => n6845, CK => Clk, RN => n3942,
                           Q => pc_lut_21_8_port, QN => n1526);
   pc_lut_reg_21_10_inst : DFFR_X1 port map( D => n6844, CK => Clk, RN => n3942
                           , Q => pc_lut_21_10_port, QN => n1525);
   pc_lut_reg_21_12_inst : DFFR_X1 port map( D => n6843, CK => Clk, RN => n3942
                           , Q => pc_lut_21_12_port, QN => n1524);
   pc_lut_reg_21_14_inst : DFFR_X1 port map( D => n6842, CK => Clk, RN => n3943
                           , Q => pc_lut_21_14_port, QN => n1523);
   pc_lut_reg_21_16_inst : DFFR_X1 port map( D => n6841, CK => Clk, RN => n3943
                           , Q => pc_lut_21_16_port, QN => n1522);
   pc_lut_reg_21_18_inst : DFFR_X1 port map( D => n6840, CK => Clk, RN => n3863
                           , Q => pc_lut_21_18_port, QN => n1521);
   pc_lut_reg_21_20_inst : DFFR_X1 port map( D => n6839, CK => Clk, RN => n3943
                           , Q => pc_lut_21_20_port, QN => n1520);
   pc_lut_reg_21_22_inst : DFFR_X1 port map( D => n6838, CK => Clk, RN => n3943
                           , Q => pc_lut_21_22_port, QN => n1519);
   pc_lut_reg_21_24_inst : DFFR_X1 port map( D => n6837, CK => Clk, RN => n3943
                           , Q => pc_lut_21_24_port, QN => n1518);
   pc_lut_reg_21_26_inst : DFFR_X1 port map( D => n6836, CK => Clk, RN => n3943
                           , Q => pc_lut_21_26_port, QN => n1517);
   pc_lut_reg_21_28_inst : DFFR_X1 port map( D => n6835, CK => Clk, RN => n3943
                           , Q => pc_lut_21_28_port, QN => n1516);
   pc_lut_reg_21_30_inst : DFFR_X1 port map( D => n6834, CK => Clk, RN => n3943
                           , Q => pc_lut_21_30_port, QN => n1514);
   pc_lut_reg_22_31_inst : DFFR_X1 port map( D => n6833, CK => Clk, RN => n3943
                           , Q => net114414, QN => n1512);
   pc_lut_reg_22_29_inst : DFFR_X1 port map( D => n6832, CK => Clk, RN => n3943
                           , Q => net114413, QN => n1511);
   pc_lut_reg_22_27_inst : DFFR_X1 port map( D => n6831, CK => Clk, RN => n3943
                           , Q => net114412, QN => n1510);
   pc_lut_reg_22_25_inst : DFFR_X1 port map( D => n6830, CK => Clk, RN => n3943
                           , Q => net114411, QN => n1509);
   pc_lut_reg_22_23_inst : DFFR_X1 port map( D => n6829, CK => Clk, RN => n3943
                           , Q => net114410, QN => n1508);
   pc_lut_reg_22_21_inst : DFFR_X1 port map( D => n6828, CK => Clk, RN => n3943
                           , Q => net114409, QN => n1507);
   pc_lut_reg_22_19_inst : DFFR_X1 port map( D => n6827, CK => Clk, RN => n3943
                           , Q => net114408, QN => n1506);
   pc_lut_reg_22_17_inst : DFFR_X1 port map( D => n6826, CK => Clk, RN => n3944
                           , Q => net114407, QN => n1505);
   pc_lut_reg_22_15_inst : DFFR_X1 port map( D => n6825, CK => Clk, RN => n3944
                           , Q => net114406, QN => n1504);
   pc_lut_reg_22_13_inst : DFFR_X1 port map( D => n6824, CK => Clk, RN => n3944
                           , Q => net114405, QN => n1503);
   pc_lut_reg_22_11_inst : DFFR_X1 port map( D => n6823, CK => Clk, RN => n3944
                           , Q => net114404, QN => n1502);
   pc_lut_reg_22_9_inst : DFFR_X1 port map( D => n6822, CK => Clk, RN => n3944,
                           Q => net114403, QN => n1501);
   pc_lut_reg_22_7_inst : DFFR_X1 port map( D => n6821, CK => Clk, RN => n3944,
                           Q => net114402, QN => n1500);
   pc_lut_reg_22_5_inst : DFFR_X1 port map( D => n6820, CK => Clk, RN => n3860,
                           Q => net114401, QN => n1499);
   pc_lut_reg_22_1_inst : DFFR_X1 port map( D => n6818, CK => Clk, RN => n3944,
                           Q => net114400, QN => n1497);
   pc_lut_reg_22_2_inst : DFFR_X1 port map( D => n6816, CK => Clk, RN => n3944,
                           Q => net114399, QN => n1495);
   pc_lut_reg_22_4_inst : DFFR_X1 port map( D => n6815, CK => Clk, RN => n3944,
                           Q => net114398, QN => n1494);
   pc_lut_reg_22_6_inst : DFFR_X1 port map( D => n6814, CK => Clk, RN => n3944,
                           Q => net114397, QN => n1493);
   pc_lut_reg_22_8_inst : DFFR_X1 port map( D => n6813, CK => Clk, RN => n3944,
                           Q => net114396, QN => n1492);
   pc_lut_reg_22_10_inst : DFFR_X1 port map( D => n6812, CK => Clk, RN => n3944
                           , Q => net114395, QN => n1491);
   pc_lut_reg_22_12_inst : DFFR_X1 port map( D => n6811, CK => Clk, RN => n3944
                           , Q => net114394, QN => n1490);
   pc_lut_reg_22_14_inst : DFFR_X1 port map( D => n6810, CK => Clk, RN => n3944
                           , Q => net114393, QN => n1489);
   pc_lut_reg_22_16_inst : DFFR_X1 port map( D => n6809, CK => Clk, RN => n3945
                           , Q => net114392, QN => n1488);
   pc_lut_reg_22_18_inst : DFFR_X1 port map( D => n6808, CK => Clk, RN => n3863
                           , Q => net114391, QN => n1487);
   pc_lut_reg_22_20_inst : DFFR_X1 port map( D => n6807, CK => Clk, RN => n3945
                           , Q => net114390, QN => n1486);
   pc_lut_reg_22_22_inst : DFFR_X1 port map( D => n6806, CK => Clk, RN => n3944
                           , Q => net114389, QN => n1485);
   pc_lut_reg_22_24_inst : DFFR_X1 port map( D => n6805, CK => Clk, RN => n3945
                           , Q => net114388, QN => n1484);
   pc_lut_reg_22_26_inst : DFFR_X1 port map( D => n6804, CK => Clk, RN => n3945
                           , Q => net114387, QN => n1483);
   pc_lut_reg_22_28_inst : DFFR_X1 port map( D => n6803, CK => Clk, RN => n3945
                           , Q => net114386, QN => n1482);
   pc_lut_reg_22_30_inst : DFFR_X1 port map( D => n6802, CK => Clk, RN => n3945
                           , Q => net114385, QN => n1480);
   pc_lut_reg_23_31_inst : DFFR_X1 port map( D => n6801, CK => Clk, RN => n3904
                           , Q => net114384, QN => n1477);
   pc_lut_reg_23_29_inst : DFFR_X1 port map( D => n6800, CK => Clk, RN => n3900
                           , Q => net114383, QN => n1476);
   pc_lut_reg_23_27_inst : DFFR_X1 port map( D => n6799, CK => Clk, RN => n3896
                           , Q => net114382, QN => n1475);
   pc_lut_reg_23_25_inst : DFFR_X1 port map( D => n6798, CK => Clk, RN => n3896
                           , Q => net114381, QN => n1474);
   pc_lut_reg_23_23_inst : DFFR_X1 port map( D => n6797, CK => Clk, RN => n3896
                           , Q => net114380, QN => n1473);
   pc_lut_reg_23_21_inst : DFFR_X1 port map( D => n6796, CK => Clk, RN => n3896
                           , Q => net114379, QN => n1472);
   pc_lut_reg_23_19_inst : DFFR_X1 port map( D => n6795, CK => Clk, RN => n3896
                           , Q => net114378, QN => n1471);
   pc_lut_reg_23_17_inst : DFFR_X1 port map( D => n6794, CK => Clk, RN => n3896
                           , Q => net114377, QN => n1470);
   pc_lut_reg_23_15_inst : DFFR_X1 port map( D => n6793, CK => Clk, RN => n3896
                           , Q => net114376, QN => n1469);
   pc_lut_reg_23_13_inst : DFFR_X1 port map( D => n6792, CK => Clk, RN => n3896
                           , Q => net114375, QN => n1468);
   pc_lut_reg_23_11_inst : DFFR_X1 port map( D => n6791, CK => Clk, RN => n3897
                           , Q => net114374, QN => n1467);
   pc_lut_reg_23_9_inst : DFFR_X1 port map( D => n6790, CK => Clk, RN => n3897,
                           Q => net114373, QN => n1466);
   pc_lut_reg_23_7_inst : DFFR_X1 port map( D => n6789, CK => Clk, RN => n3934,
                           Q => net114372, QN => n1465);
   pc_lut_reg_23_5_inst : DFFR_X1 port map( D => n6788, CK => Clk, RN => n3860,
                           Q => net114371, QN => n1464);
   pc_lut_reg_23_1_inst : DFFR_X1 port map( D => n6786, CK => Clk, RN => n3934,
                           Q => net114370, QN => n1462);
   pc_lut_reg_23_0_inst : DFFR_X1 port map( D => n6785, CK => Clk, RN => n3934,
                           Q => net114369, QN => n1461);
   pc_lut_reg_23_2_inst : DFFR_X1 port map( D => n6784, CK => Clk, RN => n3934,
                           Q => net114368, QN => n1460);
   pc_lut_reg_23_4_inst : DFFR_X1 port map( D => n6783, CK => Clk, RN => n3934,
                           Q => net114367, QN => n1459);
   pc_lut_reg_23_6_inst : DFFR_X1 port map( D => n6782, CK => Clk, RN => n3934,
                           Q => net114366, QN => n1458);
   pc_lut_reg_23_8_inst : DFFR_X1 port map( D => n6781, CK => Clk, RN => n3934,
                           Q => net114365, QN => n1457);
   pc_lut_reg_23_10_inst : DFFR_X1 port map( D => n6780, CK => Clk, RN => n3934
                           , Q => net114364, QN => n1456);
   pc_lut_reg_23_12_inst : DFFR_X1 port map( D => n6779, CK => Clk, RN => n3934
                           , Q => net114363, QN => n1455);
   pc_lut_reg_23_14_inst : DFFR_X1 port map( D => n6778, CK => Clk, RN => n3934
                           , Q => net114362, QN => n1454);
   pc_lut_reg_23_16_inst : DFFR_X1 port map( D => n6777, CK => Clk, RN => n3934
                           , Q => net114361, QN => n1453);
   pc_lut_reg_23_18_inst : DFFR_X1 port map( D => n6776, CK => Clk, RN => n3863
                           , Q => net114360, QN => n1452);
   pc_lut_reg_23_20_inst : DFFR_X1 port map( D => n6775, CK => Clk, RN => n3934
                           , Q => net114359, QN => n1451);
   pc_lut_reg_23_22_inst : DFFR_X1 port map( D => n6774, CK => Clk, RN => n3934
                           , Q => net114358, QN => n1450);
   pc_lut_reg_23_24_inst : DFFR_X1 port map( D => n6773, CK => Clk, RN => n3934
                           , Q => net114357, QN => n1449);
   pc_lut_reg_23_26_inst : DFFR_X1 port map( D => n6772, CK => Clk, RN => n3934
                           , Q => net114356, QN => n1448);
   pc_lut_reg_23_28_inst : DFFR_X1 port map( D => n6771, CK => Clk, RN => n3935
                           , Q => net114355, QN => n1447);
   pc_lut_reg_23_30_inst : DFFR_X1 port map( D => n6770, CK => Clk, RN => n3935
                           , Q => net114354, QN => n1445);
   pc_lut_reg_24_31_inst : DFFR_X1 port map( D => n6769, CK => Clk, RN => n3935
                           , Q => net114353, QN => n1443);
   pc_lut_reg_24_29_inst : DFFR_X1 port map( D => n6768, CK => Clk, RN => n3935
                           , Q => net114352, QN => n1442);
   pc_lut_reg_24_27_inst : DFFR_X1 port map( D => n6767, CK => Clk, RN => n3935
                           , Q => net114351, QN => n1441);
   pc_lut_reg_24_25_inst : DFFR_X1 port map( D => n6766, CK => Clk, RN => n3935
                           , Q => net114350, QN => n1440);
   pc_lut_reg_24_23_inst : DFFR_X1 port map( D => n6765, CK => Clk, RN => n3935
                           , Q => net114349, QN => n1439);
   pc_lut_reg_24_21_inst : DFFR_X1 port map( D => n6764, CK => Clk, RN => n3935
                           , Q => net114348, QN => n1438);
   pc_lut_reg_24_19_inst : DFFR_X1 port map( D => n6763, CK => Clk, RN => n3935
                           , Q => net114347, QN => n1437);
   pc_lut_reg_24_17_inst : DFFR_X1 port map( D => n6762, CK => Clk, RN => n3935
                           , Q => net114346, QN => n1436);
   pc_lut_reg_24_15_inst : DFFR_X1 port map( D => n6761, CK => Clk, RN => n3935
                           , Q => net114345, QN => n1435);
   pc_lut_reg_24_13_inst : DFFR_X1 port map( D => n6760, CK => Clk, RN => n3935
                           , Q => net114344, QN => n1434);
   pc_lut_reg_24_11_inst : DFFR_X1 port map( D => n6759, CK => Clk, RN => n3935
                           , Q => net114343, QN => n1433);
   pc_lut_reg_24_9_inst : DFFR_X1 port map( D => n6758, CK => Clk, RN => n3935,
                           Q => net114342, QN => n1432);
   pc_lut_reg_24_7_inst : DFFR_X1 port map( D => n6757, CK => Clk, RN => n3935,
                           Q => net114341, QN => n1431);
   pc_lut_reg_24_5_inst : DFFR_X1 port map( D => n6756, CK => Clk, RN => n3860,
                           Q => net114340, QN => n1430);
   pc_lut_reg_24_3_inst : DFFR_X1 port map( D => n6755, CK => Clk, RN => n3936,
                           Q => net114339, QN => n1429);
   pc_lut_reg_24_4_inst : DFFR_X1 port map( D => n6751, CK => Clk, RN => n3936,
                           Q => net114338, QN => n1425);
   pc_lut_reg_24_6_inst : DFFR_X1 port map( D => n6750, CK => Clk, RN => n3936,
                           Q => net114337, QN => n1424);
   pc_lut_reg_24_8_inst : DFFR_X1 port map( D => n6749, CK => Clk, RN => n3936,
                           Q => net114336, QN => n1423);
   pc_lut_reg_24_10_inst : DFFR_X1 port map( D => n6748, CK => Clk, RN => n3936
                           , Q => net114335, QN => n1422);
   pc_lut_reg_24_12_inst : DFFR_X1 port map( D => n6747, CK => Clk, RN => n3936
                           , Q => net114334, QN => n1421);
   pc_lut_reg_24_14_inst : DFFR_X1 port map( D => n6746, CK => Clk, RN => n3936
                           , Q => net114333, QN => n1420);
   pc_lut_reg_24_16_inst : DFFR_X1 port map( D => n6745, CK => Clk, RN => n3936
                           , Q => net114332, QN => n1419);
   pc_lut_reg_24_18_inst : DFFR_X1 port map( D => n6744, CK => Clk, RN => n3863
                           , Q => net114331, QN => n1418);
   pc_lut_reg_24_20_inst : DFFR_X1 port map( D => n6743, CK => Clk, RN => n3936
                           , Q => net114330, QN => n1417);
   pc_lut_reg_24_22_inst : DFFR_X1 port map( D => n6742, CK => Clk, RN => n3936
                           , Q => net114329, QN => n1416);
   pc_lut_reg_24_24_inst : DFFR_X1 port map( D => n6741, CK => Clk, RN => n3936
                           , Q => net114328, QN => n1415);
   pc_lut_reg_24_26_inst : DFFR_X1 port map( D => n6740, CK => Clk, RN => n3936
                           , Q => net114327, QN => n1414);
   pc_lut_reg_24_28_inst : DFFR_X1 port map( D => n6739, CK => Clk, RN => n3936
                           , Q => net114326, QN => n1413);
   pc_lut_reg_24_30_inst : DFFR_X1 port map( D => n6738, CK => Clk, RN => n3936
                           , Q => net114325, QN => n1411);
   pc_lut_reg_25_31_inst : DFFR_X1 port map( D => n6737, CK => Clk, RN => n3936
                           , Q => net114324, QN => n1409);
   pc_lut_reg_25_29_inst : DFFR_X1 port map( D => n6736, CK => Clk, RN => n3937
                           , Q => net114323, QN => n1408);
   pc_lut_reg_25_27_inst : DFFR_X1 port map( D => n6735, CK => Clk, RN => n3937
                           , Q => net114322, QN => n1407);
   pc_lut_reg_25_25_inst : DFFR_X1 port map( D => n6734, CK => Clk, RN => n3937
                           , Q => net114321, QN => n1406);
   pc_lut_reg_25_23_inst : DFFR_X1 port map( D => n6733, CK => Clk, RN => n3937
                           , Q => net114320, QN => n1405);
   pc_lut_reg_25_21_inst : DFFR_X1 port map( D => n6732, CK => Clk, RN => n3925
                           , Q => net114319, QN => n1404);
   pc_lut_reg_25_19_inst : DFFR_X1 port map( D => n6731, CK => Clk, RN => n3921
                           , Q => net114318, QN => n1403);
   pc_lut_reg_25_17_inst : DFFR_X1 port map( D => n6730, CK => Clk, RN => n3921
                           , Q => net114317, QN => n1402);
   pc_lut_reg_25_15_inst : DFFR_X1 port map( D => n6729, CK => Clk, RN => n3921
                           , Q => net114316, QN => n1401);
   pc_lut_reg_25_13_inst : DFFR_X1 port map( D => n6728, CK => Clk, RN => n3921
                           , Q => net114315, QN => n1400);
   pc_lut_reg_25_11_inst : DFFR_X1 port map( D => n6727, CK => Clk, RN => n3921
                           , Q => net114314, QN => n1399);
   pc_lut_reg_25_9_inst : DFFR_X1 port map( D => n6726, CK => Clk, RN => n3921,
                           Q => net114313, QN => n1398);
   pc_lut_reg_25_7_inst : DFFR_X1 port map( D => n6725, CK => Clk, RN => n3921,
                           Q => net114312, QN => n1397);
   pc_lut_reg_25_5_inst : DFFR_X1 port map( D => n6724, CK => Clk, RN => n3860,
                           Q => net114311, QN => n1396);
   pc_lut_reg_25_3_inst : DFFR_X1 port map( D => n6723, CK => Clk, RN => n3921,
                           Q => net114310, QN => n1395);
   pc_lut_reg_25_0_inst : DFFR_X1 port map( D => n6721, CK => Clk, RN => n3921,
                           Q => net114309, QN => n1393);
   pc_lut_reg_25_4_inst : DFFR_X1 port map( D => n6719, CK => Clk, RN => n3921,
                           Q => net114308, QN => n1391);
   pc_lut_reg_25_6_inst : DFFR_X1 port map( D => n6718, CK => Clk, RN => n3921,
                           Q => net114307, QN => n1390);
   pc_lut_reg_25_8_inst : DFFR_X1 port map( D => n6717, CK => Clk, RN => n3921,
                           Q => net114306, QN => n1389);
   pc_lut_reg_25_10_inst : DFFR_X1 port map( D => n6716, CK => Clk, RN => n3921
                           , Q => net114305, QN => n1388);
   pc_lut_reg_25_12_inst : DFFR_X1 port map( D => n6715, CK => Clk, RN => n3921
                           , Q => net114304, QN => n1387);
   pc_lut_reg_25_14_inst : DFFR_X1 port map( D => n6714, CK => Clk, RN => n3922
                           , Q => net114303, QN => n1386);
   pc_lut_reg_25_16_inst : DFFR_X1 port map( D => n6713, CK => Clk, RN => n3922
                           , Q => net114302, QN => n1385);
   pc_lut_reg_25_18_inst : DFFR_X1 port map( D => n6712, CK => Clk, RN => n3863
                           , Q => net114301, QN => n1384);
   pc_lut_reg_25_20_inst : DFFR_X1 port map( D => n6711, CK => Clk, RN => n3922
                           , Q => net114300, QN => n1383);
   pc_lut_reg_25_22_inst : DFFR_X1 port map( D => n6710, CK => Clk, RN => n3922
                           , Q => net114299, QN => n1382);
   pc_lut_reg_25_24_inst : DFFR_X1 port map( D => n6709, CK => Clk, RN => n3922
                           , Q => net114298, QN => n1381);
   pc_lut_reg_25_26_inst : DFFR_X1 port map( D => n6708, CK => Clk, RN => n3922
                           , Q => net114297, QN => n1380);
   pc_lut_reg_25_28_inst : DFFR_X1 port map( D => n6707, CK => Clk, RN => n3922
                           , Q => net114296, QN => n1379);
   pc_lut_reg_25_30_inst : DFFR_X1 port map( D => n6706, CK => Clk, RN => n3922
                           , Q => net114295, QN => n1377);
   pc_lut_reg_26_31_inst : DFFR_X1 port map( D => n6705, CK => Clk, RN => n3922
                           , Q => pc_lut_26_31_port, QN => n1375);
   pc_lut_reg_26_29_inst : DFFR_X1 port map( D => n6704, CK => Clk, RN => n3922
                           , Q => pc_lut_26_29_port, QN => n1374);
   pc_lut_reg_26_27_inst : DFFR_X1 port map( D => n6703, CK => Clk, RN => n3922
                           , Q => pc_lut_26_27_port, QN => n1373);
   pc_lut_reg_26_25_inst : DFFR_X1 port map( D => n6702, CK => Clk, RN => n3922
                           , Q => pc_lut_26_25_port, QN => n1372);
   pc_lut_reg_26_23_inst : DFFR_X1 port map( D => n6701, CK => Clk, RN => n3922
                           , Q => pc_lut_26_23_port, QN => n1371);
   pc_lut_reg_26_21_inst : DFFR_X1 port map( D => n6700, CK => Clk, RN => n3922
                           , Q => pc_lut_26_21_port, QN => n1370);
   pc_lut_reg_26_19_inst : DFFR_X1 port map( D => n6699, CK => Clk, RN => n3922
                           , Q => pc_lut_26_19_port, QN => n1369);
   pc_lut_reg_26_17_inst : DFFR_X1 port map( D => n6698, CK => Clk, RN => n3923
                           , Q => pc_lut_26_17_port, QN => n1368);
   pc_lut_reg_26_15_inst : DFFR_X1 port map( D => n6697, CK => Clk, RN => n3923
                           , Q => pc_lut_26_15_port, QN => n1367);
   pc_lut_reg_26_13_inst : DFFR_X1 port map( D => n6696, CK => Clk, RN => n3923
                           , Q => pc_lut_26_13_port, QN => n1366);
   pc_lut_reg_26_11_inst : DFFR_X1 port map( D => n6695, CK => Clk, RN => n3923
                           , Q => pc_lut_26_11_port, QN => n1365);
   pc_lut_reg_26_9_inst : DFFR_X1 port map( D => n6694, CK => Clk, RN => n3923,
                           Q => pc_lut_26_9_port, QN => n1364);
   pc_lut_reg_26_7_inst : DFFR_X1 port map( D => n6693, CK => Clk, RN => n3923,
                           Q => pc_lut_26_7_port, QN => n1363);
   pc_lut_reg_26_5_inst : DFFR_X1 port map( D => n6692, CK => Clk, RN => n3860,
                           Q => pc_lut_26_5_port, QN => n1362);
   pc_lut_reg_26_6_inst : DFFR_X1 port map( D => n6686, CK => Clk, RN => n3923,
                           Q => pc_lut_26_6_port, QN => n1358);
   pc_lut_reg_26_8_inst : DFFR_X1 port map( D => n6685, CK => Clk, RN => n3923,
                           Q => pc_lut_26_8_port, QN => n1357);
   pc_lut_reg_26_10_inst : DFFR_X1 port map( D => n6684, CK => Clk, RN => n3923
                           , Q => pc_lut_26_10_port, QN => n1356);
   pc_lut_reg_26_12_inst : DFFR_X1 port map( D => n6683, CK => Clk, RN => n3923
                           , Q => pc_lut_26_12_port, QN => n1355);
   pc_lut_reg_26_14_inst : DFFR_X1 port map( D => n6682, CK => Clk, RN => n3923
                           , Q => pc_lut_26_14_port, QN => n1354);
   pc_lut_reg_26_16_inst : DFFR_X1 port map( D => n6681, CK => Clk, RN => n3923
                           , Q => pc_lut_26_16_port, QN => n1353);
   pc_lut_reg_26_18_inst : DFFR_X1 port map( D => n6680, CK => Clk, RN => n3863
                           , Q => pc_lut_26_18_port, QN => n1352);
   pc_lut_reg_26_20_inst : DFFR_X1 port map( D => n6679, CK => Clk, RN => n3923
                           , Q => pc_lut_26_20_port, QN => n1351);
   pc_lut_reg_26_22_inst : DFFR_X1 port map( D => n6678, CK => Clk, RN => n3923
                           , Q => pc_lut_26_22_port, QN => n1350);
   pc_lut_reg_26_24_inst : DFFR_X1 port map( D => n6677, CK => Clk, RN => n3923
                           , Q => pc_lut_26_24_port, QN => n1349);
   pc_lut_reg_26_26_inst : DFFR_X1 port map( D => n6676, CK => Clk, RN => n3924
                           , Q => pc_lut_26_26_port, QN => n1348);
   pc_lut_reg_26_28_inst : DFFR_X1 port map( D => n6675, CK => Clk, RN => n3924
                           , Q => pc_lut_26_28_port, QN => n1347);
   pc_lut_reg_26_30_inst : DFFR_X1 port map( D => n6674, CK => Clk, RN => n3924
                           , Q => pc_lut_26_30_port, QN => n1345);
   pc_lut_reg_27_31_inst : DFFR_X1 port map( D => n6673, CK => Clk, RN => n3924
                           , Q => pc_lut_27_31_port, QN => n1342);
   pc_lut_reg_27_29_inst : DFFR_X1 port map( D => n6672, CK => Clk, RN => n3924
                           , Q => pc_lut_27_29_port, QN => n1341);
   pc_lut_reg_27_27_inst : DFFR_X1 port map( D => n6671, CK => Clk, RN => n3924
                           , Q => pc_lut_27_27_port, QN => n1340);
   pc_lut_reg_27_25_inst : DFFR_X1 port map( D => n6670, CK => Clk, RN => n3924
                           , Q => pc_lut_27_25_port, QN => n1339);
   pc_lut_reg_27_23_inst : DFFR_X1 port map( D => n6669, CK => Clk, RN => n3924
                           , Q => pc_lut_27_23_port, QN => n1338);
   pc_lut_reg_27_21_inst : DFFR_X1 port map( D => n6668, CK => Clk, RN => n3924
                           , Q => pc_lut_27_21_port, QN => n1337);
   pc_lut_reg_27_19_inst : DFFR_X1 port map( D => n6667, CK => Clk, RN => n3924
                           , Q => pc_lut_27_19_port, QN => n1336);
   pc_lut_reg_27_17_inst : DFFR_X1 port map( D => n6666, CK => Clk, RN => n3924
                           , Q => pc_lut_27_17_port, QN => n1335);
   pc_lut_reg_27_15_inst : DFFR_X1 port map( D => n6665, CK => Clk, RN => n3924
                           , Q => pc_lut_27_15_port, QN => n1334);
   pc_lut_reg_27_13_inst : DFFR_X1 port map( D => n6664, CK => Clk, RN => n3924
                           , Q => pc_lut_27_13_port, QN => n1333);
   pc_lut_reg_27_11_inst : DFFR_X1 port map( D => n6663, CK => Clk, RN => n3924
                           , Q => pc_lut_27_11_port, QN => n1332);
   pc_lut_reg_27_9_inst : DFFR_X1 port map( D => n6662, CK => Clk, RN => n3924,
                           Q => pc_lut_27_9_port, QN => n1331);
   pc_lut_reg_27_7_inst : DFFR_X1 port map( D => n6661, CK => Clk, RN => n3925,
                           Q => pc_lut_27_7_port, QN => n1330);
   pc_lut_reg_27_5_inst : DFFR_X1 port map( D => n6660, CK => Clk, RN => n3860,
                           Q => pc_lut_27_5_port, QN => n1329);
   pc_lut_reg_27_6_inst : DFFR_X1 port map( D => n6654, CK => Clk, RN => n3925,
                           Q => pc_lut_27_6_port, QN => n1324);
   pc_lut_reg_27_8_inst : DFFR_X1 port map( D => n6653, CK => Clk, RN => n3925,
                           Q => pc_lut_27_8_port, QN => n1323);
   pc_lut_reg_27_10_inst : DFFR_X1 port map( D => n6652, CK => Clk, RN => n3925
                           , Q => pc_lut_27_10_port, QN => n1322);
   pc_lut_reg_27_12_inst : DFFR_X1 port map( D => n6651, CK => Clk, RN => n3925
                           , Q => pc_lut_27_12_port, QN => n1321);
   pc_lut_reg_27_14_inst : DFFR_X1 port map( D => n6650, CK => Clk, RN => n3925
                           , Q => pc_lut_27_14_port, QN => n1320);
   pc_lut_reg_27_16_inst : DFFR_X1 port map( D => n6649, CK => Clk, RN => n3925
                           , Q => pc_lut_27_16_port, QN => n1319);
   pc_lut_reg_27_18_inst : DFFR_X1 port map( D => n6648, CK => Clk, RN => n3863
                           , Q => pc_lut_27_18_port, QN => n1318);
   pc_lut_reg_27_20_inst : DFFR_X1 port map( D => n6647, CK => Clk, RN => n3925
                           , Q => pc_lut_27_20_port, QN => n1317);
   pc_lut_reg_27_22_inst : DFFR_X1 port map( D => n6646, CK => Clk, RN => n3925
                           , Q => pc_lut_27_22_port, QN => n1316);
   pc_lut_reg_27_24_inst : DFFR_X1 port map( D => n6645, CK => Clk, RN => n3925
                           , Q => pc_lut_27_24_port, QN => n1315);
   pc_lut_reg_27_26_inst : DFFR_X1 port map( D => n6644, CK => Clk, RN => n3926
                           , Q => pc_lut_27_26_port, QN => n1314);
   pc_lut_reg_27_28_inst : DFFR_X1 port map( D => n6643, CK => Clk, RN => n3926
                           , Q => pc_lut_27_28_port, QN => n1313);
   pc_lut_reg_27_30_inst : DFFR_X1 port map( D => n6642, CK => Clk, RN => n3926
                           , Q => pc_lut_27_30_port, QN => n1311);
   pc_lut_reg_28_31_inst : DFFR_X1 port map( D => n6641, CK => Clk, RN => n3926
                           , Q => n_1006, QN => n1308);
   pc_lut_reg_28_29_inst : DFFR_X1 port map( D => n6640, CK => Clk, RN => n3926
                           , Q => n_1007, QN => n1307);
   pc_lut_reg_28_27_inst : DFFR_X1 port map( D => n6639, CK => Clk, RN => n3926
                           , Q => n_1008, QN => n1306);
   pc_lut_reg_28_25_inst : DFFR_X1 port map( D => n6638, CK => Clk, RN => n3926
                           , Q => n_1009, QN => n1305);
   pc_lut_reg_28_23_inst : DFFR_X1 port map( D => n6637, CK => Clk, RN => n3926
                           , Q => n_1010, QN => n1304);
   pc_lut_reg_28_21_inst : DFFR_X1 port map( D => n6636, CK => Clk, RN => n3926
                           , Q => n_1011, QN => n1303);
   pc_lut_reg_28_19_inst : DFFR_X1 port map( D => n6635, CK => Clk, RN => n3926
                           , Q => n_1012, QN => n1302);
   pc_lut_reg_28_17_inst : DFFR_X1 port map( D => n6634, CK => Clk, RN => n3926
                           , Q => n_1013, QN => n1301);
   pc_lut_reg_28_15_inst : DFFR_X1 port map( D => n6633, CK => Clk, RN => n3926
                           , Q => n_1014, QN => n1300);
   pc_lut_reg_28_13_inst : DFFR_X1 port map( D => n6632, CK => Clk, RN => n3926
                           , Q => n_1015, QN => n1299);
   pc_lut_reg_28_11_inst : DFFR_X1 port map( D => n6631, CK => Clk, RN => n3926
                           , Q => n_1016, QN => n1298);
   pc_lut_reg_28_9_inst : DFFR_X1 port map( D => n6630, CK => Clk, RN => n3926,
                           Q => n_1017, QN => n1297);
   pc_lut_reg_28_7_inst : DFFR_X1 port map( D => n6629, CK => Clk, RN => n3927,
                           Q => n_1018, QN => n1296);
   pc_lut_reg_28_5_inst : DFFR_X1 port map( D => n6628, CK => Clk, RN => n3860,
                           Q => n_1019, QN => n1295);
   pc_lut_reg_28_6_inst : DFFR_X1 port map( D => n6622, CK => Clk, RN => n3927,
                           Q => n_1020, QN => n1289);
   pc_lut_reg_28_8_inst : DFFR_X1 port map( D => n6621, CK => Clk, RN => n3927,
                           Q => n_1021, QN => n1288);
   pc_lut_reg_28_10_inst : DFFR_X1 port map( D => n6620, CK => Clk, RN => n3927
                           , Q => n_1022, QN => n1287);
   pc_lut_reg_28_12_inst : DFFR_X1 port map( D => n6619, CK => Clk, RN => n3927
                           , Q => n_1023, QN => n1286);
   pc_lut_reg_28_14_inst : DFFR_X1 port map( D => n6618, CK => Clk, RN => n3927
                           , Q => n_1024, QN => n1285);
   pc_lut_reg_28_16_inst : DFFR_X1 port map( D => n6617, CK => Clk, RN => n3927
                           , Q => n_1025, QN => n1284);
   pc_lut_reg_28_18_inst : DFFR_X1 port map( D => n6616, CK => Clk, RN => n3863
                           , Q => n_1026, QN => n1283);
   pc_lut_reg_28_20_inst : DFFR_X1 port map( D => n6615, CK => Clk, RN => n3927
                           , Q => n_1027, QN => n1282);
   pc_lut_reg_28_22_inst : DFFR_X1 port map( D => n6614, CK => Clk, RN => n3927
                           , Q => n_1028, QN => n1281);
   pc_lut_reg_28_24_inst : DFFR_X1 port map( D => n6613, CK => Clk, RN => n3927
                           , Q => n_1029, QN => n1280);
   pc_lut_reg_28_26_inst : DFFR_X1 port map( D => n6612, CK => Clk, RN => n3927
                           , Q => n_1030, QN => n1279);
   pc_lut_reg_28_28_inst : DFFR_X1 port map( D => n6611, CK => Clk, RN => n3927
                           , Q => n_1031, QN => n1278);
   pc_lut_reg_28_30_inst : DFFR_X1 port map( D => n6610, CK => Clk, RN => n3927
                           , Q => n_1032, QN => n1276);
   pc_lut_reg_29_31_inst : DFFR_X1 port map( D => n6609, CK => Clk, RN => n3927
                           , Q => n_1033, QN => n1274);
   pc_lut_reg_29_29_inst : DFFR_X1 port map( D => n6608, CK => Clk, RN => n3927
                           , Q => n_1034, QN => n1273);
   pc_lut_reg_29_27_inst : DFFR_X1 port map( D => n6607, CK => Clk, RN => n3928
                           , Q => n_1035, QN => n1272);
   pc_lut_reg_29_25_inst : DFFR_X1 port map( D => n6606, CK => Clk, RN => n3928
                           , Q => n_1036, QN => n1271);
   pc_lut_reg_29_23_inst : DFFR_X1 port map( D => n6605, CK => Clk, RN => n3928
                           , Q => n_1037, QN => n1270);
   pc_lut_reg_29_21_inst : DFFR_X1 port map( D => n6604, CK => Clk, RN => n3928
                           , Q => n_1038, QN => n1269);
   pc_lut_reg_29_19_inst : DFFR_X1 port map( D => n6603, CK => Clk, RN => n3928
                           , Q => n_1039, QN => n1268);
   pc_lut_reg_29_17_inst : DFFR_X1 port map( D => n6602, CK => Clk, RN => n3928
                           , Q => n_1040, QN => n1267);
   pc_lut_reg_29_15_inst : DFFR_X1 port map( D => n6601, CK => Clk, RN => n3928
                           , Q => n_1041, QN => n1266);
   pc_lut_reg_29_13_inst : DFFR_X1 port map( D => n6600, CK => Clk, RN => n3928
                           , Q => n_1042, QN => n1265);
   pc_lut_reg_29_11_inst : DFFR_X1 port map( D => n6599, CK => Clk, RN => n3928
                           , Q => n_1043, QN => n1264);
   pc_lut_reg_29_9_inst : DFFR_X1 port map( D => n6598, CK => Clk, RN => n3928,
                           Q => n_1044, QN => n1263);
   pc_lut_reg_29_7_inst : DFFR_X1 port map( D => n6597, CK => Clk, RN => n3928,
                           Q => n_1045, QN => n1262);
   pc_lut_reg_29_5_inst : DFFR_X1 port map( D => n6596, CK => Clk, RN => n3860,
                           Q => n_1046, QN => n1261);
   pc_lut_reg_29_6_inst : DFFR_X1 port map( D => n6590, CK => Clk, RN => n3928,
                           Q => n_1047, QN => n1254);
   pc_lut_reg_29_8_inst : DFFR_X1 port map( D => n6589, CK => Clk, RN => n3928,
                           Q => n_1048, QN => n1253);
   pc_lut_reg_29_10_inst : DFFR_X1 port map( D => n6588, CK => Clk, RN => n3928
                           , Q => n_1049, QN => n1252);
   pc_lut_reg_29_12_inst : DFFR_X1 port map( D => n6587, CK => Clk, RN => n3928
                           , Q => n_1050, QN => n1251);
   pc_lut_reg_29_14_inst : DFFR_X1 port map( D => n6586, CK => Clk, RN => n3929
                           , Q => n_1051, QN => n1250);
   pc_lut_reg_29_16_inst : DFFR_X1 port map( D => n6585, CK => Clk, RN => n3929
                           , Q => n_1052, QN => n1249);
   pc_lut_reg_29_18_inst : DFFR_X1 port map( D => n6584, CK => Clk, RN => n3884
                           , Q => n_1053, QN => n1248);
   pc_lut_reg_29_20_inst : DFFR_X1 port map( D => n6583, CK => Clk, RN => n3929
                           , Q => n_1054, QN => n1247);
   pc_lut_reg_29_22_inst : DFFR_X1 port map( D => n6582, CK => Clk, RN => n3949
                           , Q => n_1055, QN => n1246);
   pc_lut_reg_29_24_inst : DFFR_X1 port map( D => n6581, CK => Clk, RN => n3945
                           , Q => n_1056, QN => n1245);
   pc_lut_reg_29_26_inst : DFFR_X1 port map( D => n6580, CK => Clk, RN => n3945
                           , Q => n_1057, QN => n1244);
   pc_lut_reg_29_28_inst : DFFR_X1 port map( D => n6579, CK => Clk, RN => n3945
                           , Q => n_1058, QN => n1243);
   pc_lut_reg_29_30_inst : DFFR_X1 port map( D => n6578, CK => Clk, RN => n3945
                           , Q => n_1059, QN => n1241);
   pc_lut_reg_30_31_inst : DFFR_X1 port map( D => n6577, CK => Clk, RN => n3945
                           , Q => pc_lut_30_31_port, QN => n1239);
   pc_lut_reg_30_29_inst : DFFR_X1 port map( D => n6576, CK => Clk, RN => n3945
                           , Q => pc_lut_30_29_port, QN => n1238);
   pc_lut_reg_30_27_inst : DFFR_X1 port map( D => n6575, CK => Clk, RN => n3945
                           , Q => pc_lut_30_27_port, QN => n1237);
   pc_lut_reg_30_25_inst : DFFR_X1 port map( D => n6574, CK => Clk, RN => n3945
                           , Q => pc_lut_30_25_port, QN => n1236);
   pc_lut_reg_30_23_inst : DFFR_X1 port map( D => n6573, CK => Clk, RN => n3945
                           , Q => pc_lut_30_23_port, QN => n1235);
   pc_lut_reg_30_21_inst : DFFR_X1 port map( D => n6572, CK => Clk, RN => n3946
                           , Q => pc_lut_30_21_port, QN => n1234);
   pc_lut_reg_30_19_inst : DFFR_X1 port map( D => n6571, CK => Clk, RN => n3946
                           , Q => pc_lut_30_19_port, QN => n1233);
   pc_lut_reg_30_17_inst : DFFR_X1 port map( D => n6570, CK => Clk, RN => n3946
                           , Q => pc_lut_30_17_port, QN => n1232);
   pc_lut_reg_30_15_inst : DFFR_X1 port map( D => n6569, CK => Clk, RN => n3946
                           , Q => pc_lut_30_15_port, QN => n1231);
   pc_lut_reg_30_13_inst : DFFR_X1 port map( D => n6568, CK => Clk, RN => n3946
                           , Q => pc_lut_30_13_port, QN => n1230);
   pc_lut_reg_30_11_inst : DFFR_X1 port map( D => n6567, CK => Clk, RN => n3946
                           , Q => pc_lut_30_11_port, QN => n1229);
   pc_lut_reg_30_9_inst : DFFR_X1 port map( D => n6566, CK => Clk, RN => n3946,
                           Q => pc_lut_30_9_port, QN => n1228);
   pc_lut_reg_30_7_inst : DFFR_X1 port map( D => n6565, CK => Clk, RN => n3946,
                           Q => pc_lut_30_7_port, QN => n1227);
   pc_lut_reg_30_5_inst : DFFR_X1 port map( D => n6564, CK => Clk, RN => n3861,
                           Q => pc_lut_30_5_port, QN => n1226);
   pc_lut_reg_30_3_inst : DFFR_X1 port map( D => n6563, CK => Clk, RN => n3946,
                           Q => pc_lut_30_3_port, QN => net114209);
   pc_lut_reg_30_1_inst : DFFR_X1 port map( D => n6562, CK => Clk, RN => n3946,
                           Q => pc_lut_30_1_port, QN => net114208);
   pc_lut_reg_30_2_inst : DFFR_X1 port map( D => n6560, CK => Clk, RN => n3946,
                           Q => pc_lut_30_2_port, QN => net114207);
   pc_lut_reg_30_4_inst : DFFR_X1 port map( D => n6559, CK => Clk, RN => n3946,
                           Q => pc_lut_30_4_port, QN => net114206);
   pc_lut_reg_30_6_inst : DFFR_X1 port map( D => n6558, CK => Clk, RN => n3946,
                           Q => pc_lut_30_6_port, QN => n1221);
   pc_lut_reg_30_8_inst : DFFR_X1 port map( D => n6557, CK => Clk, RN => n3946,
                           Q => pc_lut_30_8_port, QN => n1220);
   pc_lut_reg_30_10_inst : DFFR_X1 port map( D => n6556, CK => Clk, RN => n3946
                           , Q => pc_lut_30_10_port, QN => n1219);
   pc_lut_reg_30_12_inst : DFFR_X1 port map( D => n6555, CK => Clk, RN => n3947
                           , Q => pc_lut_30_12_port, QN => n1218);
   pc_lut_reg_30_14_inst : DFFR_X1 port map( D => n6554, CK => Clk, RN => n3947
                           , Q => pc_lut_30_14_port, QN => n1217);
   pc_lut_reg_30_16_inst : DFFR_X1 port map( D => n6553, CK => Clk, RN => n3947
                           , Q => pc_lut_30_16_port, QN => n1216);
   pc_lut_reg_30_18_inst : DFFR_X1 port map( D => n6552, CK => Clk, RN => n3880
                           , Q => pc_lut_30_18_port, QN => n1215);
   pc_lut_reg_30_20_inst : DFFR_X1 port map( D => n6551, CK => Clk, RN => n3947
                           , Q => pc_lut_30_20_port, QN => n1214);
   pc_lut_reg_30_22_inst : DFFR_X1 port map( D => n6550, CK => Clk, RN => n3947
                           , Q => pc_lut_30_22_port, QN => n1213);
   pc_lut_reg_30_24_inst : DFFR_X1 port map( D => n6549, CK => Clk, RN => n3947
                           , Q => pc_lut_30_24_port, QN => n1212);
   pc_lut_reg_30_26_inst : DFFR_X1 port map( D => n6548, CK => Clk, RN => n3947
                           , Q => pc_lut_30_26_port, QN => n1211);
   pc_lut_reg_30_28_inst : DFFR_X1 port map( D => n6547, CK => Clk, RN => n3947
                           , Q => pc_lut_30_28_port, QN => n1210);
   pc_lut_reg_30_30_inst : DFFR_X1 port map( D => n6546, CK => Clk, RN => n3947
                           , Q => pc_lut_30_30_port, QN => n1208);
   pc_lut_reg_31_31_inst : DFFR_X1 port map( D => n6545, CK => Clk, RN => n3947
                           , Q => pc_lut_31_31_port, QN => n1204);
   pc_lut_reg_31_29_inst : DFFR_X1 port map( D => n6544, CK => Clk, RN => n3841
                           , Q => pc_lut_31_29_port, QN => n1202);
   pc_lut_reg_31_27_inst : DFFR_X1 port map( D => n6543, CK => Clk, RN => n3841
                           , Q => pc_lut_31_27_port, QN => n1200);
   pc_lut_reg_31_25_inst : DFFR_X1 port map( D => n6542, CK => Clk, RN => n3894
                           , Q => pc_lut_31_25_port, QN => n1198);
   pc_lut_reg_31_23_inst : DFFR_X1 port map( D => n6541, CK => Clk, RN => n3841
                           , Q => pc_lut_31_23_port, QN => n1196);
   pc_lut_reg_31_21_inst : DFFR_X1 port map( D => n6540, CK => Clk, RN => n3841
                           , Q => pc_lut_31_21_port, QN => n1194);
   pc_lut_reg_31_19_inst : DFFR_X1 port map( D => n6539, CK => Clk, RN => n3841
                           , Q => pc_lut_31_19_port, QN => n1192);
   pc_lut_reg_31_17_inst : DFFR_X1 port map( D => n6538, CK => Clk, RN => n3841
                           , Q => pc_lut_31_17_port, QN => n1190);
   pc_lut_reg_31_15_inst : DFFR_X1 port map( D => n6537, CK => Clk, RN => n3842
                           , Q => pc_lut_31_15_port, QN => n1188);
   pc_lut_reg_31_13_inst : DFFR_X1 port map( D => n6536, CK => Clk, RN => n3842
                           , Q => pc_lut_31_13_port, QN => n1186);
   pc_lut_reg_31_11_inst : DFFR_X1 port map( D => n6535, CK => Clk, RN => n3842
                           , Q => pc_lut_31_11_port, QN => n1184);
   pc_lut_reg_31_9_inst : DFFR_X1 port map( D => n6534, CK => Clk, RN => n3842,
                           Q => pc_lut_31_9_port, QN => n1182);
   pc_lut_reg_31_7_inst : DFFR_X1 port map( D => n6533, CK => Clk, RN => n3842,
                           Q => pc_lut_31_7_port, QN => n1180);
   pc_lut_reg_31_5_inst : DFFR_X1 port map( D => n6532, CK => Clk, RN => n3861,
                           Q => pc_lut_31_5_port, QN => n1178);
   pc_lut_reg_31_6_inst : DFFR_X1 port map( D => n6526, CK => Clk, RN => n3842,
                           Q => pc_lut_31_6_port, QN => n1171);
   pc_lut_reg_31_8_inst : DFFR_X1 port map( D => n6525, CK => Clk, RN => n3842,
                           Q => pc_lut_31_8_port, QN => n1169);
   pc_lut_reg_31_10_inst : DFFR_X1 port map( D => n6524, CK => Clk, RN => n3842
                           , Q => pc_lut_31_10_port, QN => n1167);
   pc_lut_reg_31_12_inst : DFFR_X1 port map( D => n6523, CK => Clk, RN => n3842
                           , Q => pc_lut_31_12_port, QN => n1165);
   pc_lut_reg_31_14_inst : DFFR_X1 port map( D => n6522, CK => Clk, RN => n3842
                           , Q => pc_lut_31_14_port, QN => n1163);
   pc_lut_reg_31_16_inst : DFFR_X1 port map( D => n6521, CK => Clk, RN => n3843
                           , Q => pc_lut_31_16_port, QN => n1161);
   pc_lut_reg_31_18_inst : DFFR_X1 port map( D => n6520, CK => Clk, RN => n3880
                           , Q => pc_lut_31_18_port, QN => n1159);
   pc_lut_reg_31_20_inst : DFFR_X1 port map( D => n6519, CK => Clk, RN => n3843
                           , Q => pc_lut_31_20_port, QN => n1157);
   pc_lut_reg_31_22_inst : DFFR_X1 port map( D => n6518, CK => Clk, RN => n3843
                           , Q => pc_lut_31_22_port, QN => n1155);
   pc_lut_reg_31_24_inst : DFFR_X1 port map( D => n6517, CK => Clk, RN => n3843
                           , Q => pc_lut_31_24_port, QN => n1153);
   pc_lut_reg_31_26_inst : DFFR_X1 port map( D => n6516, CK => Clk, RN => n3843
                           , Q => pc_lut_31_26_port, QN => n1151);
   pc_lut_reg_31_28_inst : DFFR_X1 port map( D => n6515, CK => Clk, RN => n3843
                           , Q => pc_lut_31_28_port, QN => n1149);
   pc_lut_reg_31_30_inst : DFFR_X1 port map( D => n6514, CK => Clk, RN => n3844
                           , Q => pc_lut_31_30_port, QN => n1146);
   OUTT_NTs_reg : DLH_X1 port map( G => Enable, D => N220, Q => OUTT_NT_port);
   pc_target_reg_0_31_inst : DFFR_X1 port map( D => n6513, CK => Clk, RN => 
                           n3864, Q => net114200, QN => n1142);
   pc_target_reg_0_29_inst : DFFR_X1 port map( D => n6512, CK => Clk, RN => 
                           n3843, Q => net114199, QN => n1141);
   pc_target_reg_0_27_inst : DFFR_X1 port map( D => n6511, CK => Clk, RN => 
                           n3843, Q => net114198, QN => n1140);
   pc_target_reg_0_25_inst : DFFR_X1 port map( D => n6510, CK => Clk, RN => 
                           n3843, Q => net114197, QN => n1139);
   pc_target_reg_0_23_inst : DFFR_X1 port map( D => n6509, CK => Clk, RN => 
                           n3843, Q => net114196, QN => n1138);
   pc_target_reg_0_21_inst : DFFR_X1 port map( D => n6508, CK => Clk, RN => 
                           n3843, Q => net114195, QN => n1137);
   pc_target_reg_0_19_inst : DFFR_X1 port map( D => n6507, CK => Clk, RN => 
                           n3843, Q => net114194, QN => n1136);
   pc_target_reg_0_17_inst : DFFR_X1 port map( D => n6506, CK => Clk, RN => 
                           n3843, Q => net114193, QN => n1135);
   pc_target_reg_0_15_inst : DFFR_X1 port map( D => n6505, CK => Clk, RN => 
                           n3843, Q => net114192, QN => n1134);
   pc_target_reg_0_13_inst : DFFR_X1 port map( D => n6504, CK => Clk, RN => 
                           n3844, Q => net114191, QN => n1133);
   pc_target_reg_0_11_inst : DFFR_X1 port map( D => n6503, CK => Clk, RN => 
                           n3844, Q => net114190, QN => n1132);
   pc_target_reg_0_9_inst : DFFR_X1 port map( D => n6502, CK => Clk, RN => 
                           n3844, Q => net114189, QN => n1131);
   pc_target_reg_0_7_inst : DFFR_X1 port map( D => n6501, CK => Clk, RN => 
                           n3844, Q => net114188, QN => n1130);
   pc_target_reg_0_5_inst : DFFR_X1 port map( D => n6500, CK => Clk, RN => 
                           n3844, Q => n_1060, QN => n1129);
   pc_target_reg_0_3_inst : DFFR_X1 port map( D => n6499, CK => Clk, RN => 
                           n3844, Q => net114186, QN => n1128);
   pc_target_reg_0_1_inst : DFFR_X1 port map( D => n6498, CK => Clk, RN => 
                           n3844, Q => n_1061, QN => n1127);
   pc_target_reg_0_0_inst : DFFR_X1 port map( D => n6497, CK => Clk, RN => 
                           n3844, Q => n_1062, QN => n1126);
   pc_target_reg_0_2_inst : DFFR_X1 port map( D => n6496, CK => Clk, RN => 
                           n3844, Q => net114183, QN => n1125);
   pc_target_reg_0_4_inst : DFFR_X1 port map( D => n6495, CK => Clk, RN => 
                           n3844, Q => n_1063, QN => n1124);
   pc_target_reg_0_6_inst : DFFR_X1 port map( D => n6494, CK => Clk, RN => 
                           n3844, Q => n_1064, QN => n1123);
   pc_target_reg_0_8_inst : DFFR_X1 port map( D => n6493, CK => Clk, RN => 
                           n3844, Q => net114180, QN => n1122);
   pc_target_reg_0_10_inst : DFFR_X1 port map( D => n6492, CK => Clk, RN => 
                           n3844, Q => net114179, QN => n1121);
   pc_target_reg_0_12_inst : DFFR_X1 port map( D => n6491, CK => Clk, RN => 
                           n3844, Q => net114178, QN => n1120);
   pc_target_reg_0_14_inst : DFFR_X1 port map( D => n6490, CK => Clk, RN => 
                           n3845, Q => net114177, QN => n1119);
   pc_target_reg_0_16_inst : DFFR_X1 port map( D => n6489, CK => Clk, RN => 
                           n3845, Q => net114176, QN => n1118);
   pc_target_reg_0_18_inst : DFFR_X1 port map( D => n6488, CK => Clk, RN => 
                           n3845, Q => net114175, QN => n1117);
   pc_target_reg_0_20_inst : DFFR_X1 port map( D => n6487, CK => Clk, RN => 
                           n3845, Q => net114174, QN => n1116);
   pc_target_reg_0_22_inst : DFFR_X1 port map( D => n6486, CK => Clk, RN => 
                           n3845, Q => net114173, QN => n1115);
   pc_target_reg_0_24_inst : DFFR_X1 port map( D => n6485, CK => Clk, RN => 
                           n3845, Q => net114172, QN => n1114);
   pc_target_reg_0_26_inst : DFFR_X1 port map( D => n6484, CK => Clk, RN => 
                           n3845, Q => net114171, QN => n1113);
   pc_target_reg_0_28_inst : DFFR_X1 port map( D => n6483, CK => Clk, RN => 
                           n3845, Q => net114170, QN => n1112);
   pc_target_reg_1_31_inst : DFFR_X1 port map( D => n6481, CK => Clk, RN => 
                           n3865, Q => net114169, QN => n1108);
   pc_target_reg_1_29_inst : DFFR_X1 port map( D => n6480, CK => Clk, RN => 
                           n3845, Q => net114168, QN => n1107);
   pc_target_reg_1_27_inst : DFFR_X1 port map( D => n6479, CK => Clk, RN => 
                           n3845, Q => net114167, QN => n1106);
   pc_target_reg_1_25_inst : DFFR_X1 port map( D => n6478, CK => Clk, RN => 
                           n3845, Q => net114166, QN => n1105);
   pc_target_reg_1_23_inst : DFFR_X1 port map( D => n6477, CK => Clk, RN => 
                           n3845, Q => net114165, QN => n1104);
   pc_target_reg_1_21_inst : DFFR_X1 port map( D => n6476, CK => Clk, RN => 
                           n3845, Q => net114164, QN => n1103);
   pc_target_reg_1_19_inst : DFFR_X1 port map( D => n6475, CK => Clk, RN => 
                           n3845, Q => net114163, QN => n1102);
   pc_target_reg_1_17_inst : DFFR_X1 port map( D => n6474, CK => Clk, RN => 
                           n3845, Q => net114162, QN => n1101);
   pc_target_reg_1_15_inst : DFFR_X1 port map( D => n6473, CK => Clk, RN => 
                           n3846, Q => net114161, QN => n1100);
   pc_target_reg_1_13_inst : DFFR_X1 port map( D => n6472, CK => Clk, RN => 
                           n3846, Q => net114160, QN => n1099);
   pc_target_reg_1_11_inst : DFFR_X1 port map( D => n6471, CK => Clk, RN => 
                           n3846, Q => net114159, QN => n1098);
   pc_target_reg_1_9_inst : DFFR_X1 port map( D => n6470, CK => Clk, RN => 
                           n3846, Q => net114158, QN => n1097);
   pc_target_reg_1_7_inst : DFFR_X1 port map( D => n6469, CK => Clk, RN => 
                           n3846, Q => net114157, QN => n1096);
   pc_target_reg_1_5_inst : DFFR_X1 port map( D => n6468, CK => Clk, RN => 
                           n3846, Q => n_1065, QN => n1095);
   pc_target_reg_1_3_inst : DFFR_X1 port map( D => n6467, CK => Clk, RN => 
                           n3846, Q => net114155, QN => n1094);
   pc_target_reg_1_1_inst : DFFR_X1 port map( D => n6466, CK => Clk, RN => 
                           n3846, Q => n_1066, QN => n1093);
   pc_target_reg_1_0_inst : DFFR_X1 port map( D => n6465, CK => Clk, RN => 
                           n3847, Q => n_1067, QN => n1092);
   pc_target_reg_1_2_inst : DFFR_X1 port map( D => n6464, CK => Clk, RN => 
                           n3846, Q => net114152, QN => n1091);
   pc_target_reg_1_4_inst : DFFR_X1 port map( D => n6463, CK => Clk, RN => 
                           n3846, Q => n_1068, QN => n1090);
   pc_target_reg_1_6_inst : DFFR_X1 port map( D => n6462, CK => Clk, RN => 
                           n3846, Q => n_1069, QN => n1089);
   pc_target_reg_1_8_inst : DFFR_X1 port map( D => n6461, CK => Clk, RN => 
                           n3846, Q => net114149, QN => n1088);
   pc_target_reg_1_10_inst : DFFR_X1 port map( D => n6460, CK => Clk, RN => 
                           n3846, Q => net114148, QN => n1087);
   pc_target_reg_1_12_inst : DFFR_X1 port map( D => n6459, CK => Clk, RN => 
                           n3846, Q => net114147, QN => n1086);
   pc_target_reg_1_14_inst : DFFR_X1 port map( D => n6458, CK => Clk, RN => 
                           n3846, Q => net114146, QN => n1085);
   pc_target_reg_1_16_inst : DFFR_X1 port map( D => n6457, CK => Clk, RN => 
                           n3847, Q => net114145, QN => n1084);
   pc_target_reg_1_18_inst : DFFR_X1 port map( D => n6456, CK => Clk, RN => 
                           n3847, Q => net114144, QN => n1083);
   pc_target_reg_1_20_inst : DFFR_X1 port map( D => n6455, CK => Clk, RN => 
                           n3847, Q => net114143, QN => n1082);
   pc_target_reg_1_22_inst : DFFR_X1 port map( D => n6454, CK => Clk, RN => 
                           n3847, Q => net114142, QN => n1081);
   pc_target_reg_1_24_inst : DFFR_X1 port map( D => n6453, CK => Clk, RN => 
                           n3847, Q => net114141, QN => n1080);
   pc_target_reg_1_26_inst : DFFR_X1 port map( D => n6452, CK => Clk, RN => 
                           n3847, Q => net114140, QN => n1079);
   pc_target_reg_1_28_inst : DFFR_X1 port map( D => n6451, CK => Clk, RN => 
                           n3847, Q => net114139, QN => n1078);
   pc_target_reg_3_31_inst : DFFR_X1 port map( D => n6417, CK => Clk, RN => 
                           n3864, Q => pc_target_3_31_port, QN => net114138);
   pc_target_reg_3_29_inst : DFFR_X1 port map( D => n6416, CK => Clk, RN => 
                           n3847, Q => pc_target_3_29_port, QN => net114137);
   pc_target_reg_3_27_inst : DFFR_X1 port map( D => n6415, CK => Clk, RN => 
                           n3847, Q => pc_target_3_27_port, QN => net114136);
   pc_target_reg_3_25_inst : DFFR_X1 port map( D => n6414, CK => Clk, RN => 
                           n3847, Q => pc_target_3_25_port, QN => net114135);
   pc_target_reg_3_23_inst : DFFR_X1 port map( D => n6413, CK => Clk, RN => 
                           n3847, Q => pc_target_3_23_port, QN => net114134);
   pc_target_reg_3_21_inst : DFFR_X1 port map( D => n6412, CK => Clk, RN => 
                           n3847, Q => pc_target_3_21_port, QN => net114133);
   pc_target_reg_3_19_inst : DFFR_X1 port map( D => n6411, CK => Clk, RN => 
                           n3855, Q => pc_target_3_19_port, QN => net114132);
   pc_target_reg_3_17_inst : DFFR_X1 port map( D => n6410, CK => Clk, RN => 
                           n3937, Q => pc_target_3_17_port, QN => net114131);
   pc_target_reg_3_15_inst : DFFR_X1 port map( D => n6409, CK => Clk, RN => 
                           n3933, Q => pc_target_3_15_port, QN => net114130);
   pc_target_reg_3_13_inst : DFFR_X1 port map( D => n6408, CK => Clk, RN => 
                           n3929, Q => pc_target_3_13_port, QN => net114129);
   pc_target_reg_3_11_inst : DFFR_X1 port map( D => n6407, CK => Clk, RN => 
                           n3929, Q => pc_target_3_11_port, QN => net114128);
   pc_target_reg_3_7_inst : DFFR_X1 port map( D => n6405, CK => Clk, RN => 
                           n3929, Q => pc_target_3_7_port, QN => net114127);
   pc_target_reg_3_12_inst : DFFR_X1 port map( D => n6395, CK => Clk, RN => 
                           n3929, Q => pc_target_3_12_port, QN => net114126);
   pc_target_reg_3_14_inst : DFFR_X1 port map( D => n6394, CK => Clk, RN => 
                           n3929, Q => pc_target_3_14_port, QN => net114125);
   pc_target_reg_3_16_inst : DFFR_X1 port map( D => n6393, CK => Clk, RN => 
                           n3929, Q => pc_target_3_16_port, QN => net114124);
   pc_target_reg_3_18_inst : DFFR_X1 port map( D => n6392, CK => Clk, RN => 
                           n3929, Q => pc_target_3_18_port, QN => net114123);
   pc_target_reg_3_20_inst : DFFR_X1 port map( D => n6391, CK => Clk, RN => 
                           n3929, Q => pc_target_3_20_port, QN => net114122);
   pc_target_reg_3_22_inst : DFFR_X1 port map( D => n6390, CK => Clk, RN => 
                           n3930, Q => pc_target_3_22_port, QN => net114121);
   pc_target_reg_3_24_inst : DFFR_X1 port map( D => n6389, CK => Clk, RN => 
                           n3930, Q => pc_target_3_24_port, QN => net114120);
   pc_target_reg_3_26_inst : DFFR_X1 port map( D => n6388, CK => Clk, RN => 
                           n3930, Q => pc_target_3_26_port, QN => net114119);
   pc_target_reg_3_28_inst : DFFR_X1 port map( D => n6387, CK => Clk, RN => 
                           n3930, Q => pc_target_3_28_port, QN => net114118);
   pc_target_reg_3_30_inst : DFFR_X1 port map( D => n6386, CK => Clk, RN => 
                           n3930, Q => pc_target_3_30_port, QN => net114117);
   pc_target_reg_4_31_inst : DFFR_X1 port map( D => n6385, CK => Clk, RN => 
                           n3864, Q => net114116, QN => n1005);
   pc_target_reg_4_29_inst : DFFR_X1 port map( D => n6384, CK => Clk, RN => 
                           n3929, Q => net114115, QN => n1004);
   pc_target_reg_4_27_inst : DFFR_X1 port map( D => n6383, CK => Clk, RN => 
                           n3929, Q => net114114, QN => n1003);
   pc_target_reg_4_25_inst : DFFR_X1 port map( D => n6382, CK => Clk, RN => 
                           n3929, Q => net114113, QN => n1002);
   pc_target_reg_4_23_inst : DFFR_X1 port map( D => n6381, CK => Clk, RN => 
                           n3929, Q => net114112, QN => n1001);
   pc_target_reg_4_21_inst : DFFR_X1 port map( D => n6380, CK => Clk, RN => 
                           n3930, Q => net114111, QN => n1000);
   pc_target_reg_4_19_inst : DFFR_X1 port map( D => n6379, CK => Clk, RN => 
                           n3930, Q => net114110, QN => n999);
   pc_target_reg_4_17_inst : DFFR_X1 port map( D => n6378, CK => Clk, RN => 
                           n3930, Q => net114109, QN => n998);
   pc_target_reg_4_15_inst : DFFR_X1 port map( D => n6377, CK => Clk, RN => 
                           n3930, Q => net114108, QN => n997);
   pc_target_reg_4_13_inst : DFFR_X1 port map( D => n6376, CK => Clk, RN => 
                           n3930, Q => net114107, QN => n996);
   pc_target_reg_4_11_inst : DFFR_X1 port map( D => n6375, CK => Clk, RN => 
                           n3930, Q => net114106, QN => n995);
   pc_target_reg_4_9_inst : DFFR_X1 port map( D => n6374, CK => Clk, RN => 
                           n3930, Q => net114105, QN => n994);
   pc_target_reg_4_7_inst : DFFR_X1 port map( D => n6373, CK => Clk, RN => 
                           n3930, Q => net114104, QN => n993);
   pc_target_reg_4_3_inst : DFFR_X1 port map( D => n6371, CK => Clk, RN => 
                           n3930, Q => net114103, QN => n991);
   pc_target_reg_4_1_inst : DFFR_X1 port map( D => n6370, CK => Clk, RN => 
                           n3930, Q => n_1070, QN => n990);
   pc_target_reg_4_0_inst : DFFR_X1 port map( D => n6369, CK => Clk, RN => 
                           n3931, Q => n_1071, QN => n989);
   pc_target_reg_4_2_inst : DFFR_X1 port map( D => n6368, CK => Clk, RN => 
                           n3931, Q => net114100, QN => n988);
   pc_target_reg_4_6_inst : DFFR_X1 port map( D => n6366, CK => Clk, RN => 
                           n3931, Q => n_1072, QN => n986);
   pc_target_reg_4_8_inst : DFFR_X1 port map( D => n6365, CK => Clk, RN => 
                           n3931, Q => net114098, QN => n985);
   pc_target_reg_4_10_inst : DFFR_X1 port map( D => n6364, CK => Clk, RN => 
                           n3931, Q => net114097, QN => n984);
   pc_target_reg_4_12_inst : DFFR_X1 port map( D => n6363, CK => Clk, RN => 
                           n3931, Q => net114096, QN => n983);
   pc_target_reg_4_14_inst : DFFR_X1 port map( D => n6362, CK => Clk, RN => 
                           n3931, Q => net114095, QN => n982);
   pc_target_reg_4_16_inst : DFFR_X1 port map( D => n6361, CK => Clk, RN => 
                           n3931, Q => net114094, QN => n981);
   pc_target_reg_4_18_inst : DFFR_X1 port map( D => n6360, CK => Clk, RN => 
                           n3931, Q => net114093, QN => n980);
   pc_target_reg_4_20_inst : DFFR_X1 port map( D => n6359, CK => Clk, RN => 
                           n3931, Q => net114092, QN => n979);
   pc_target_reg_4_22_inst : DFFR_X1 port map( D => n6358, CK => Clk, RN => 
                           n3931, Q => net114091, QN => n978);
   pc_target_reg_4_24_inst : DFFR_X1 port map( D => n6357, CK => Clk, RN => 
                           n3931, Q => net114090, QN => n977);
   pc_target_reg_4_26_inst : DFFR_X1 port map( D => n6356, CK => Clk, RN => 
                           n3932, Q => net114089, QN => n976);
   pc_target_reg_4_28_inst : DFFR_X1 port map( D => n6355, CK => Clk, RN => 
                           n3932, Q => net114088, QN => n975);
   pc_target_reg_5_31_inst : DFFR_X1 port map( D => n6353, CK => Clk, RN => 
                           n3864, Q => net114087, QN => n971);
   pc_target_reg_5_29_inst : DFFR_X1 port map( D => n6352, CK => Clk, RN => 
                           n3931, Q => net114086, QN => n970);
   pc_target_reg_5_27_inst : DFFR_X1 port map( D => n6351, CK => Clk, RN => 
                           n3931, Q => net114085, QN => n969);
   pc_target_reg_5_25_inst : DFFR_X1 port map( D => n6350, CK => Clk, RN => 
                           n3931, Q => net114084, QN => n968);
   pc_target_reg_5_23_inst : DFFR_X1 port map( D => n6349, CK => Clk, RN => 
                           n3932, Q => net114083, QN => n967);
   pc_target_reg_5_21_inst : DFFR_X1 port map( D => n6348, CK => Clk, RN => 
                           n3932, Q => net114082, QN => n966);
   pc_target_reg_5_19_inst : DFFR_X1 port map( D => n6347, CK => Clk, RN => 
                           n3932, Q => net114081, QN => n965);
   pc_target_reg_5_17_inst : DFFR_X1 port map( D => n6346, CK => Clk, RN => 
                           n3932, Q => net114080, QN => n964);
   pc_target_reg_5_15_inst : DFFR_X1 port map( D => n6345, CK => Clk, RN => 
                           n3932, Q => net114079, QN => n963);
   pc_target_reg_5_13_inst : DFFR_X1 port map( D => n6344, CK => Clk, RN => 
                           n3932, Q => net114078, QN => n962);
   pc_target_reg_5_11_inst : DFFR_X1 port map( D => n6343, CK => Clk, RN => 
                           n3932, Q => net114077, QN => n961);
   pc_target_reg_5_9_inst : DFFR_X1 port map( D => n6342, CK => Clk, RN => 
                           n3932, Q => net114076, QN => n960);
   pc_target_reg_5_7_inst : DFFR_X1 port map( D => n6341, CK => Clk, RN => 
                           n3932, Q => net114075, QN => n959);
   pc_target_reg_5_5_inst : DFFR_X1 port map( D => n6340, CK => Clk, RN => 
                           n3932, Q => net114074, QN => n958);
   pc_target_reg_5_3_inst : DFFR_X1 port map( D => n6339, CK => Clk, RN => 
                           n3932, Q => net114073, QN => n957);
   pc_target_reg_5_1_inst : DFFR_X1 port map( D => n6338, CK => Clk, RN => 
                           n3932, Q => net114072, QN => n956);
   pc_target_reg_5_0_inst : DFFR_X1 port map( D => n6337, CK => Clk, RN => 
                           n3933, Q => net114071, QN => n955);
   pc_target_reg_5_2_inst : DFFR_X1 port map( D => n6336, CK => Clk, RN => 
                           n3932, Q => net114070, QN => n954);
   pc_target_reg_5_4_inst : DFFR_X1 port map( D => n6335, CK => Clk, RN => 
                           n3933, Q => net114069, QN => n953);
   pc_target_reg_5_6_inst : DFFR_X1 port map( D => n6334, CK => Clk, RN => 
                           n3933, Q => net114068, QN => n952);
   pc_target_reg_5_8_inst : DFFR_X1 port map( D => n6333, CK => Clk, RN => 
                           n3933, Q => net114067, QN => n951);
   pc_target_reg_5_10_inst : DFFR_X1 port map( D => n6332, CK => Clk, RN => 
                           n3933, Q => net114066, QN => n950);
   pc_target_reg_5_12_inst : DFFR_X1 port map( D => n6331, CK => Clk, RN => 
                           n3933, Q => net114065, QN => n949);
   pc_target_reg_5_14_inst : DFFR_X1 port map( D => n6330, CK => Clk, RN => 
                           n3933, Q => net114064, QN => n948);
   pc_target_reg_5_16_inst : DFFR_X1 port map( D => n6329, CK => Clk, RN => 
                           n3933, Q => net114063, QN => n947);
   pc_target_reg_5_18_inst : DFFR_X1 port map( D => n6328, CK => Clk, RN => 
                           n3933, Q => net114062, QN => n946);
   pc_target_reg_5_20_inst : DFFR_X1 port map( D => n6327, CK => Clk, RN => 
                           n3933, Q => net114061, QN => n945);
   pc_target_reg_5_22_inst : DFFR_X1 port map( D => n6326, CK => Clk, RN => 
                           n3933, Q => net114060, QN => n944);
   pc_target_reg_5_24_inst : DFFR_X1 port map( D => n6325, CK => Clk, RN => 
                           n3933, Q => net114059, QN => n943);
   pc_target_reg_5_26_inst : DFFR_X1 port map( D => n6324, CK => Clk, RN => 
                           n3933, Q => net114058, QN => n942);
   pc_target_reg_5_28_inst : DFFR_X1 port map( D => n6323, CK => Clk, RN => 
                           n3933, Q => net114057, QN => n941);
   pc_target_reg_7_5_inst : DFFR_X1 port map( D => n6276, CK => Clk, RN => 
                           n3830, Q => pc_target_7_5_port, QN => net114043);
   pc_target_reg_7_3_inst : DFFR_X1 port map( D => n6275, CK => Clk, RN => 
                           n3830, Q => pc_target_7_3_port, QN => net114042);
   pc_target_reg_7_1_inst : DFFR_X1 port map( D => n6274, CK => Clk, RN => 
                           n3830, Q => pc_target_7_1_port, QN => net114041);
   pc_target_reg_7_0_inst : DFFR_X1 port map( D => n6273, CK => Clk, RN => 
                           n3831, Q => pc_target_7_0_port, QN => net114040);
   pc_target_reg_7_2_inst : DFFR_X1 port map( D => n6272, CK => Clk, RN => 
                           n3830, Q => pc_target_7_2_port, QN => net114039);
   pc_target_reg_7_4_inst : DFFR_X1 port map( D => n6271, CK => Clk, RN => 
                           n3830, Q => pc_target_7_4_port, QN => net114038);
   pc_target_reg_7_6_inst : DFFR_X1 port map( D => n6270, CK => Clk, RN => 
                           n3830, Q => pc_target_7_6_port, QN => net114037);
   pc_target_reg_8_31_inst : DFFR_X1 port map( D => n6257, CK => Clk, RN => 
                           n3865, Q => net114024, QN => n868);
   pc_target_reg_8_29_inst : DFFR_X1 port map( D => n6256, CK => Clk, RN => 
                           n3831, Q => net114023, QN => n867);
   pc_target_reg_8_27_inst : DFFR_X1 port map( D => n6255, CK => Clk, RN => 
                           n3831, Q => net114022, QN => n866);
   pc_target_reg_8_25_inst : DFFR_X1 port map( D => n6254, CK => Clk, RN => 
                           n3832, Q => net114021, QN => n865);
   pc_target_reg_8_23_inst : DFFR_X1 port map( D => n6253, CK => Clk, RN => 
                           n3832, Q => net114020, QN => n864);
   pc_target_reg_8_21_inst : DFFR_X1 port map( D => n6252, CK => Clk, RN => 
                           n3832, Q => net114019, QN => n863);
   pc_target_reg_8_19_inst : DFFR_X1 port map( D => n6251, CK => Clk, RN => 
                           n3832, Q => net114018, QN => n862);
   pc_target_reg_8_17_inst : DFFR_X1 port map( D => n6250, CK => Clk, RN => 
                           n3832, Q => net114017, QN => n861);
   pc_target_reg_8_15_inst : DFFR_X1 port map( D => n6249, CK => Clk, RN => 
                           n3832, Q => net114016, QN => n860);
   pc_target_reg_8_13_inst : DFFR_X1 port map( D => n6248, CK => Clk, RN => 
                           n3851, Q => net114015, QN => n859);
   pc_target_reg_8_11_inst : DFFR_X1 port map( D => n6247, CK => Clk, RN => 
                           n3847, Q => net114014, QN => n858);
   pc_target_reg_8_9_inst : DFFR_X1 port map( D => n6246, CK => Clk, RN => 
                           n3847, Q => net114013, QN => n857);
   pc_target_reg_8_7_inst : DFFR_X1 port map( D => n6245, CK => Clk, RN => 
                           n3848, Q => net114012, QN => n856);
   pc_target_reg_8_5_inst : DFFR_X1 port map( D => n6244, CK => Clk, RN => 
                           n3848, Q => net114011, QN => n855);
   pc_target_reg_8_3_inst : DFFR_X1 port map( D => n6243, CK => Clk, RN => 
                           n3848, Q => net114010, QN => n854);
   pc_target_reg_8_1_inst : DFFR_X1 port map( D => n6242, CK => Clk, RN => 
                           n3848, Q => net114009, QN => n853);
   pc_target_reg_8_0_inst : DFFR_X1 port map( D => n6241, CK => Clk, RN => 
                           n3848, Q => net114008, QN => n852);
   pc_target_reg_8_2_inst : DFFR_X1 port map( D => n6240, CK => Clk, RN => 
                           n3848, Q => net114007, QN => n851);
   pc_target_reg_8_4_inst : DFFR_X1 port map( D => n6239, CK => Clk, RN => 
                           n3848, Q => net114006, QN => n850);
   pc_target_reg_8_6_inst : DFFR_X1 port map( D => n6238, CK => Clk, RN => 
                           n3848, Q => net114005, QN => n849);
   pc_target_reg_8_8_inst : DFFR_X1 port map( D => n6237, CK => Clk, RN => 
                           n3848, Q => net114004, QN => n848);
   pc_target_reg_8_10_inst : DFFR_X1 port map( D => n6236, CK => Clk, RN => 
                           n3848, Q => net114003, QN => n847);
   pc_target_reg_8_12_inst : DFFR_X1 port map( D => n6235, CK => Clk, RN => 
                           n3848, Q => net114002, QN => n846);
   pc_target_reg_8_14_inst : DFFR_X1 port map( D => n6234, CK => Clk, RN => 
                           n3848, Q => net114001, QN => n845);
   pc_target_reg_8_16_inst : DFFR_X1 port map( D => n6233, CK => Clk, RN => 
                           n3848, Q => net114000, QN => n844);
   pc_target_reg_8_18_inst : DFFR_X1 port map( D => n6232, CK => Clk, RN => 
                           n3848, Q => net113999, QN => n843);
   pc_target_reg_8_20_inst : DFFR_X1 port map( D => n6231, CK => Clk, RN => 
                           n3848, Q => net113998, QN => n842);
   pc_target_reg_8_22_inst : DFFR_X1 port map( D => n6230, CK => Clk, RN => 
                           n3849, Q => net113997, QN => n841);
   pc_target_reg_8_24_inst : DFFR_X1 port map( D => n6229, CK => Clk, RN => 
                           n3849, Q => net113996, QN => n840);
   pc_target_reg_8_26_inst : DFFR_X1 port map( D => n6228, CK => Clk, RN => 
                           n3849, Q => net113995, QN => n839);
   pc_target_reg_8_28_inst : DFFR_X1 port map( D => n6227, CK => Clk, RN => 
                           n3849, Q => net113994, QN => n838);
   pc_target_reg_9_31_inst : DFFR_X1 port map( D => n6225, CK => Clk, RN => 
                           n3865, Q => net113993, QN => n834);
   pc_target_reg_9_29_inst : DFFR_X1 port map( D => n6224, CK => Clk, RN => 
                           n3849, Q => net113992, QN => n833);
   pc_target_reg_9_27_inst : DFFR_X1 port map( D => n6223, CK => Clk, RN => 
                           n3849, Q => net113991, QN => n832);
   pc_target_reg_9_25_inst : DFFR_X1 port map( D => n6222, CK => Clk, RN => 
                           n3849, Q => net113990, QN => n831);
   pc_target_reg_9_23_inst : DFFR_X1 port map( D => n6221, CK => Clk, RN => 
                           n3849, Q => net113989, QN => n830);
   pc_target_reg_9_21_inst : DFFR_X1 port map( D => n6220, CK => Clk, RN => 
                           n3849, Q => net113988, QN => n829);
   pc_target_reg_9_19_inst : DFFR_X1 port map( D => n6219, CK => Clk, RN => 
                           n3849, Q => net113987, QN => n828);
   pc_target_reg_9_17_inst : DFFR_X1 port map( D => n6218, CK => Clk, RN => 
                           n3849, Q => net113986, QN => n827);
   pc_target_reg_9_15_inst : DFFR_X1 port map( D => n6217, CK => Clk, RN => 
                           n3849, Q => net113985, QN => n826);
   pc_target_reg_9_13_inst : DFFR_X1 port map( D => n6216, CK => Clk, RN => 
                           n3849, Q => net113984, QN => n825);
   pc_target_reg_9_11_inst : DFFR_X1 port map( D => n6215, CK => Clk, RN => 
                           n3849, Q => net113983, QN => n824);
   pc_target_reg_9_9_inst : DFFR_X1 port map( D => n6214, CK => Clk, RN => 
                           n3849, Q => net113982, QN => n823);
   pc_target_reg_9_7_inst : DFFR_X1 port map( D => n6213, CK => Clk, RN => 
                           n3850, Q => net113981, QN => n822);
   pc_target_reg_9_3_inst : DFFR_X1 port map( D => n6211, CK => Clk, RN => 
                           n3850, Q => net113980, QN => n820);
   pc_target_reg_9_1_inst : DFFR_X1 port map( D => n6210, CK => Clk, RN => 
                           n3850, Q => n_1073, QN => n819);
   pc_target_reg_9_0_inst : DFFR_X1 port map( D => n6209, CK => Clk, RN => 
                           n3850, Q => n_1074, QN => n818);
   pc_target_reg_9_2_inst : DFFR_X1 port map( D => n6208, CK => Clk, RN => 
                           n3850, Q => net113977, QN => n817);
   pc_target_reg_9_6_inst : DFFR_X1 port map( D => n6206, CK => Clk, RN => 
                           n3850, Q => n_1075, QN => n815);
   pc_target_reg_9_8_inst : DFFR_X1 port map( D => n6205, CK => Clk, RN => 
                           n3850, Q => net113975, QN => n814);
   pc_target_reg_9_10_inst : DFFR_X1 port map( D => n6204, CK => Clk, RN => 
                           n3850, Q => net113974, QN => n813);
   pc_target_reg_9_12_inst : DFFR_X1 port map( D => n6203, CK => Clk, RN => 
                           n3850, Q => net113973, QN => n812);
   pc_target_reg_9_14_inst : DFFR_X1 port map( D => n6202, CK => Clk, RN => 
                           n3850, Q => net113972, QN => n811);
   pc_target_reg_9_16_inst : DFFR_X1 port map( D => n6201, CK => Clk, RN => 
                           n3850, Q => net113971, QN => n810);
   pc_target_reg_9_18_inst : DFFR_X1 port map( D => n6200, CK => Clk, RN => 
                           n3850, Q => net113970, QN => n809);
   pc_target_reg_9_20_inst : DFFR_X1 port map( D => n6199, CK => Clk, RN => 
                           n3850, Q => net113969, QN => n808);
   pc_target_reg_9_22_inst : DFFR_X1 port map( D => n6198, CK => Clk, RN => 
                           n3850, Q => net113968, QN => n807);
   pc_target_reg_9_24_inst : DFFR_X1 port map( D => n6197, CK => Clk, RN => 
                           n3850, Q => net113967, QN => n806);
   pc_target_reg_9_26_inst : DFFR_X1 port map( D => n6196, CK => Clk, RN => 
                           n3851, Q => net113966, QN => n805);
   pc_target_reg_9_28_inst : DFFR_X1 port map( D => n6195, CK => Clk, RN => 
                           n3851, Q => net113965, QN => n804);
   pc_target_reg_10_31_inst : DFFR_X1 port map( D => n6193, CK => Clk, RN => 
                           n3864, Q => pc_target_10_31_port, QN => net113964);
   pc_target_reg_10_29_inst : DFFR_X1 port map( D => n6192, CK => Clk, RN => 
                           n3851, Q => pc_target_10_29_port, QN => net113963);
   pc_target_reg_10_27_inst : DFFR_X1 port map( D => n6191, CK => Clk, RN => 
                           n3851, Q => pc_target_10_27_port, QN => net113962);
   pc_target_reg_10_25_inst : DFFR_X1 port map( D => n6190, CK => Clk, RN => 
                           n3851, Q => pc_target_10_25_port, QN => net113961);
   pc_target_reg_10_23_inst : DFFR_X1 port map( D => n6189, CK => Clk, RN => 
                           n3851, Q => pc_target_10_23_port, QN => net113960);
   pc_target_reg_10_21_inst : DFFR_X1 port map( D => n6188, CK => Clk, RN => 
                           n3851, Q => pc_target_10_21_port, QN => net113959);
   pc_target_reg_10_19_inst : DFFR_X1 port map( D => n6187, CK => Clk, RN => 
                           n3851, Q => pc_target_10_19_port, QN => net113958);
   pc_target_reg_10_17_inst : DFFR_X1 port map( D => n6186, CK => Clk, RN => 
                           n3851, Q => pc_target_10_17_port, QN => net113957);
   pc_target_reg_10_15_inst : DFFR_X1 port map( D => n6185, CK => Clk, RN => 
                           n3851, Q => pc_target_10_15_port, QN => net113956);
   pc_target_reg_10_13_inst : DFFR_X1 port map( D => n6184, CK => Clk, RN => 
                           n3851, Q => pc_target_10_13_port, QN => net113955);
   pc_target_reg_10_11_inst : DFFR_X1 port map( D => n6183, CK => Clk, RN => 
                           n3851, Q => pc_target_10_11_port, QN => net113954);
   pc_target_reg_10_7_inst : DFFR_X1 port map( D => n6181, CK => Clk, RN => 
                           n3851, Q => pc_target_10_7_port, QN => net113953);
   pc_target_reg_10_5_inst : DFFR_X1 port map( D => n6180, CK => Clk, RN => 
                           n3851, Q => pc_target_10_5_port, QN => net113952);
   pc_target_reg_10_1_inst : DFFR_X1 port map( D => n6178, CK => Clk, RN => 
                           n3852, Q => pc_target_10_1_port, QN => net113951);
   pc_target_reg_10_0_inst : DFFR_X1 port map( D => n6177, CK => Clk, RN => 
                           n3852, Q => pc_target_10_0_port, QN => net113950);
   pc_target_reg_10_2_inst : DFFR_X1 port map( D => n6176, CK => Clk, RN => 
                           n3852, Q => pc_target_10_2_port, QN => net113949);
   pc_target_reg_10_4_inst : DFFR_X1 port map( D => n6175, CK => Clk, RN => 
                           n3852, Q => pc_target_10_4_port, QN => net113948);
   pc_target_reg_10_6_inst : DFFR_X1 port map( D => n6174, CK => Clk, RN => 
                           n3852, Q => pc_target_10_6_port, QN => net113947);
   pc_target_reg_10_12_inst : DFFR_X1 port map( D => n6171, CK => Clk, RN => 
                           n3852, Q => pc_target_10_12_port, QN => net113946);
   pc_target_reg_10_14_inst : DFFR_X1 port map( D => n6170, CK => Clk, RN => 
                           n3852, Q => pc_target_10_14_port, QN => net113945);
   pc_target_reg_10_16_inst : DFFR_X1 port map( D => n6169, CK => Clk, RN => 
                           n3852, Q => pc_target_10_16_port, QN => net113944);
   pc_target_reg_10_18_inst : DFFR_X1 port map( D => n6168, CK => Clk, RN => 
                           n3852, Q => pc_target_10_18_port, QN => net113943);
   pc_target_reg_10_20_inst : DFFR_X1 port map( D => n6167, CK => Clk, RN => 
                           n3852, Q => pc_target_10_20_port, QN => net113942);
   pc_target_reg_10_22_inst : DFFR_X1 port map( D => n6166, CK => Clk, RN => 
                           n3852, Q => pc_target_10_22_port, QN => net113941);
   pc_target_reg_10_24_inst : DFFR_X1 port map( D => n6165, CK => Clk, RN => 
                           n3853, Q => pc_target_10_24_port, QN => net113940);
   pc_target_reg_10_26_inst : DFFR_X1 port map( D => n6164, CK => Clk, RN => 
                           n3853, Q => pc_target_10_26_port, QN => net113939);
   pc_target_reg_10_28_inst : DFFR_X1 port map( D => n6163, CK => Clk, RN => 
                           n3853, Q => pc_target_10_28_port, QN => net113938);
   pc_target_reg_10_30_inst : DFFR_X1 port map( D => n6162, CK => Clk, RN => 
                           n3852, Q => pc_target_10_30_port, QN => net113937);
   pc_target_reg_11_31_inst : DFFR_X1 port map( D => n6161, CK => Clk, RN => 
                           n3864, Q => pc_target_11_31_port, QN => net113936);
   pc_target_reg_11_29_inst : DFFR_X1 port map( D => n6160, CK => Clk, RN => 
                           n3852, Q => pc_target_11_29_port, QN => net113935);
   pc_target_reg_11_27_inst : DFFR_X1 port map( D => n6159, CK => Clk, RN => 
                           n3852, Q => pc_target_11_27_port, QN => net113934);
   pc_target_reg_11_25_inst : DFFR_X1 port map( D => n6158, CK => Clk, RN => 
                           n3852, Q => pc_target_11_25_port, QN => net113933);
   pc_target_reg_11_23_inst : DFFR_X1 port map( D => n6157, CK => Clk, RN => 
                           n3853, Q => pc_target_11_23_port, QN => net113932);
   pc_target_reg_11_21_inst : DFFR_X1 port map( D => n6156, CK => Clk, RN => 
                           n3853, Q => pc_target_11_21_port, QN => net113931);
   pc_target_reg_11_19_inst : DFFR_X1 port map( D => n6155, CK => Clk, RN => 
                           n3853, Q => pc_target_11_19_port, QN => net113930);
   pc_target_reg_11_17_inst : DFFR_X1 port map( D => n6154, CK => Clk, RN => 
                           n3853, Q => pc_target_11_17_port, QN => net113929);
   pc_target_reg_11_15_inst : DFFR_X1 port map( D => n6153, CK => Clk, RN => 
                           n3853, Q => pc_target_11_15_port, QN => net113928);
   pc_target_reg_11_13_inst : DFFR_X1 port map( D => n6152, CK => Clk, RN => 
                           n3853, Q => pc_target_11_13_port, QN => net113927);
   pc_target_reg_11_11_inst : DFFR_X1 port map( D => n6151, CK => Clk, RN => 
                           n3853, Q => pc_target_11_11_port, QN => net113926);
   pc_target_reg_11_9_inst : DFFR_X1 port map( D => n6150, CK => Clk, RN => 
                           n3853, Q => pc_target_11_9_port, QN => net113925);
   pc_target_reg_11_7_inst : DFFR_X1 port map( D => n6149, CK => Clk, RN => 
                           n3853, Q => pc_target_11_7_port, QN => net113924);
   pc_target_reg_11_5_inst : DFFR_X1 port map( D => n6148, CK => Clk, RN => 
                           n3853, Q => pc_target_11_5_port, QN => net113923);
   pc_target_reg_11_3_inst : DFFR_X1 port map( D => n6147, CK => Clk, RN => 
                           n3853, Q => pc_target_11_3_port, QN => net113922);
   pc_target_reg_11_1_inst : DFFR_X1 port map( D => n6146, CK => Clk, RN => 
                           n3853, Q => pc_target_11_1_port, QN => net113921);
   pc_target_reg_11_0_inst : DFFR_X1 port map( D => n6145, CK => Clk, RN => 
                           n3854, Q => pc_target_11_0_port, QN => net113920);
   pc_target_reg_11_2_inst : DFFR_X1 port map( D => n6144, CK => Clk, RN => 
                           n3854, Q => pc_target_11_2_port, QN => net113919);
   pc_target_reg_11_4_inst : DFFR_X1 port map( D => n6143, CK => Clk, RN => 
                           n3854, Q => pc_target_11_4_port, QN => net113918);
   pc_target_reg_11_6_inst : DFFR_X1 port map( D => n6142, CK => Clk, RN => 
                           n3854, Q => pc_target_11_6_port, QN => net113917);
   pc_target_reg_11_8_inst : DFFR_X1 port map( D => n6141, CK => Clk, RN => 
                           n3854, Q => pc_target_11_8_port, QN => net113916);
   pc_target_reg_11_10_inst : DFFR_X1 port map( D => n6140, CK => Clk, RN => 
                           n3854, Q => pc_target_11_10_port, QN => net113915);
   pc_target_reg_11_12_inst : DFFR_X1 port map( D => n6139, CK => Clk, RN => 
                           n3854, Q => pc_target_11_12_port, QN => net113914);
   pc_target_reg_11_14_inst : DFFR_X1 port map( D => n6138, CK => Clk, RN => 
                           n3854, Q => pc_target_11_14_port, QN => net113913);
   pc_target_reg_11_16_inst : DFFR_X1 port map( D => n6137, CK => Clk, RN => 
                           n3854, Q => pc_target_11_16_port, QN => net113912);
   pc_target_reg_11_18_inst : DFFR_X1 port map( D => n6136, CK => Clk, RN => 
                           n3854, Q => pc_target_11_18_port, QN => net113911);
   pc_target_reg_11_20_inst : DFFR_X1 port map( D => n6135, CK => Clk, RN => 
                           n3854, Q => pc_target_11_20_port, QN => net113910);
   pc_target_reg_11_22_inst : DFFR_X1 port map( D => n6134, CK => Clk, RN => 
                           n3854, Q => pc_target_11_22_port, QN => net113909);
   pc_target_reg_11_24_inst : DFFR_X1 port map( D => n6133, CK => Clk, RN => 
                           n3854, Q => pc_target_11_24_port, QN => net113908);
   pc_target_reg_11_26_inst : DFFR_X1 port map( D => n6132, CK => Clk, RN => 
                           n3854, Q => pc_target_11_26_port, QN => net113907);
   pc_target_reg_11_28_inst : DFFR_X1 port map( D => n6131, CK => Clk, RN => 
                           n3854, Q => pc_target_11_28_port, QN => net113906);
   pc_target_reg_11_30_inst : DFFR_X1 port map( D => n6130, CK => Clk, RN => 
                           n3855, Q => pc_target_11_30_port, QN => net113905);
   pc_target_reg_12_31_inst : DFFR_X1 port map( D => n6129, CK => Clk, RN => 
                           n3865, Q => net113904, QN => n730);
   pc_target_reg_12_29_inst : DFFR_X1 port map( D => n6128, CK => Clk, RN => 
                           n3855, Q => net113903, QN => n729);
   pc_target_reg_12_27_inst : DFFR_X1 port map( D => n6127, CK => Clk, RN => 
                           n3855, Q => net113902, QN => n728);
   pc_target_reg_12_25_inst : DFFR_X1 port map( D => n6126, CK => Clk, RN => 
                           n3855, Q => net113901, QN => n727);
   pc_target_reg_12_23_inst : DFFR_X1 port map( D => n6125, CK => Clk, RN => 
                           n3855, Q => net113900, QN => n726);
   pc_target_reg_12_21_inst : DFFR_X1 port map( D => n6124, CK => Clk, RN => 
                           n3855, Q => net113899, QN => n725);
   pc_target_reg_12_19_inst : DFFR_X1 port map( D => n6123, CK => Clk, RN => 
                           n3855, Q => net113898, QN => n724);
   pc_target_reg_12_17_inst : DFFR_X1 port map( D => n6122, CK => Clk, RN => 
                           n3855, Q => net113897, QN => n723);
   pc_target_reg_12_15_inst : DFFR_X1 port map( D => n6121, CK => Clk, RN => 
                           n3855, Q => net113896, QN => n722);
   pc_target_reg_12_13_inst : DFFR_X1 port map( D => n6120, CK => Clk, RN => 
                           n3843, Q => net113895, QN => n721);
   pc_target_reg_12_11_inst : DFFR_X1 port map( D => n6119, CK => Clk, RN => 
                           n3840, Q => net113894, QN => n720);
   pc_target_reg_12_9_inst : DFFR_X1 port map( D => n6118, CK => Clk, RN => 
                           n3840, Q => net113893, QN => n719);
   pc_target_reg_12_7_inst : DFFR_X1 port map( D => n6117, CK => Clk, RN => 
                           n3840, Q => net113892, QN => n718);
   pc_target_reg_12_5_inst : DFFR_X1 port map( D => n6116, CK => Clk, RN => 
                           n3840, Q => n_1076, QN => n717);
   pc_target_reg_12_3_inst : DFFR_X1 port map( D => n6115, CK => Clk, RN => 
                           n3840, Q => net113890, QN => n716);
   pc_target_reg_12_1_inst : DFFR_X1 port map( D => n6114, CK => Clk, RN => 
                           n3840, Q => n_1077, QN => n715);
   pc_target_reg_12_0_inst : DFFR_X1 port map( D => n6113, CK => Clk, RN => 
                           n3840, Q => n_1078, QN => n714);
   pc_target_reg_12_2_inst : DFFR_X1 port map( D => n6112, CK => Clk, RN => 
                           n3840, Q => net113887, QN => n713);
   pc_target_reg_12_4_inst : DFFR_X1 port map( D => n6111, CK => Clk, RN => 
                           n3840, Q => n_1079, QN => n712);
   pc_target_reg_12_6_inst : DFFR_X1 port map( D => n6110, CK => Clk, RN => 
                           n3840, Q => n_1080, QN => n711);
   pc_target_reg_12_8_inst : DFFR_X1 port map( D => n6109, CK => Clk, RN => 
                           n3840, Q => net113884, QN => n710);
   pc_target_reg_12_10_inst : DFFR_X1 port map( D => n6108, CK => Clk, RN => 
                           n3840, Q => net113883, QN => n709);
   pc_target_reg_12_12_inst : DFFR_X1 port map( D => n6107, CK => Clk, RN => 
                           n3840, Q => net113882, QN => n708);
   pc_target_reg_12_14_inst : DFFR_X1 port map( D => n6106, CK => Clk, RN => 
                           n3841, Q => net113881, QN => n707);
   pc_target_reg_12_16_inst : DFFR_X1 port map( D => n6105, CK => Clk, RN => 
                           n3841, Q => net113880, QN => n706);
   pc_target_reg_12_18_inst : DFFR_X1 port map( D => n6104, CK => Clk, RN => 
                           n3841, Q => net113879, QN => n705);
   pc_target_reg_12_20_inst : DFFR_X1 port map( D => n6103, CK => Clk, RN => 
                           n3841, Q => net113878, QN => n704);
   pc_target_reg_12_22_inst : DFFR_X1 port map( D => n6102, CK => Clk, RN => 
                           n3841, Q => net113877, QN => n703);
   pc_target_reg_12_24_inst : DFFR_X1 port map( D => n6101, CK => Clk, RN => 
                           n3841, Q => net113876, QN => n702);
   pc_target_reg_12_26_inst : DFFR_X1 port map( D => n6100, CK => Clk, RN => 
                           n3841, Q => net113875, QN => n701);
   pc_target_reg_12_28_inst : DFFR_X1 port map( D => n6099, CK => Clk, RN => 
                           n3841, Q => net113874, QN => n700);
   pc_target_reg_13_31_inst : DFFR_X1 port map( D => n6097, CK => Clk, RN => 
                           n3865, Q => net113873, QN => n696);
   pc_target_reg_13_29_inst : DFFR_X1 port map( D => n6096, CK => Clk, RN => 
                           n3841, Q => net113872, QN => n695);
   pc_target_reg_13_27_inst : DFFR_X1 port map( D => n6095, CK => Clk, RN => 
                           n3877, Q => net113871, QN => n694);
   pc_target_reg_13_25_inst : DFFR_X1 port map( D => n6094, CK => Clk, RN => 
                           n3877, Q => net113870, QN => n693);
   pc_target_reg_13_23_inst : DFFR_X1 port map( D => n6093, CK => Clk, RN => 
                           n3877, Q => net113869, QN => n692);
   pc_target_reg_13_21_inst : DFFR_X1 port map( D => n6092, CK => Clk, RN => 
                           n3877, Q => net113868, QN => n691);
   pc_target_reg_13_19_inst : DFFR_X1 port map( D => n6091, CK => Clk, RN => 
                           n3877, Q => net113867, QN => n690);
   pc_target_reg_13_17_inst : DFFR_X1 port map( D => n6090, CK => Clk, RN => 
                           n3877, Q => net113866, QN => n689);
   pc_target_reg_13_15_inst : DFFR_X1 port map( D => n6089, CK => Clk, RN => 
                           n3878, Q => net113865, QN => n688);
   pc_target_reg_13_13_inst : DFFR_X1 port map( D => n6088, CK => Clk, RN => 
                           n3878, Q => net113864, QN => n687);
   pc_target_reg_13_11_inst : DFFR_X1 port map( D => n6087, CK => Clk, RN => 
                           n3878, Q => net113863, QN => n686);
   pc_target_reg_13_9_inst : DFFR_X1 port map( D => n6086, CK => Clk, RN => 
                           n3878, Q => net113862, QN => n685);
   pc_target_reg_13_7_inst : DFFR_X1 port map( D => n6085, CK => Clk, RN => 
                           n3878, Q => net113861, QN => n684);
   pc_target_reg_13_5_inst : DFFR_X1 port map( D => n6084, CK => Clk, RN => 
                           n3878, Q => n_1081, QN => n683);
   pc_target_reg_13_3_inst : DFFR_X1 port map( D => n6083, CK => Clk, RN => 
                           n3878, Q => net113859, QN => n682);
   pc_target_reg_13_1_inst : DFFR_X1 port map( D => n6082, CK => Clk, RN => 
                           n3878, Q => n_1082, QN => n681);
   pc_target_reg_13_0_inst : DFFR_X1 port map( D => n6081, CK => Clk, RN => 
                           n3879, Q => n_1083, QN => n680);
   pc_target_reg_13_2_inst : DFFR_X1 port map( D => n6080, CK => Clk, RN => 
                           n3878, Q => net113856, QN => n679);
   pc_target_reg_13_4_inst : DFFR_X1 port map( D => n6079, CK => Clk, RN => 
                           n3878, Q => n_1084, QN => n678);
   pc_target_reg_13_6_inst : DFFR_X1 port map( D => n6078, CK => Clk, RN => 
                           n3878, Q => n_1085, QN => n677);
   pc_target_reg_13_8_inst : DFFR_X1 port map( D => n6077, CK => Clk, RN => 
                           n3878, Q => net113853, QN => n676);
   pc_target_reg_13_10_inst : DFFR_X1 port map( D => n6076, CK => Clk, RN => 
                           n3878, Q => net113852, QN => n675);
   pc_target_reg_13_12_inst : DFFR_X1 port map( D => n6075, CK => Clk, RN => 
                           n3878, Q => net113851, QN => n674);
   pc_target_reg_13_14_inst : DFFR_X1 port map( D => n6074, CK => Clk, RN => 
                           n3878, Q => net113850, QN => n673);
   pc_target_reg_13_16_inst : DFFR_X1 port map( D => n6073, CK => Clk, RN => 
                           n3879, Q => net113849, QN => n672);
   pc_target_reg_13_18_inst : DFFR_X1 port map( D => n6072, CK => Clk, RN => 
                           n3879, Q => net113848, QN => n671);
   pc_target_reg_13_20_inst : DFFR_X1 port map( D => n6071, CK => Clk, RN => 
                           n3879, Q => net113847, QN => n670);
   pc_target_reg_13_22_inst : DFFR_X1 port map( D => n6070, CK => Clk, RN => 
                           n3879, Q => net113846, QN => n669);
   pc_target_reg_13_24_inst : DFFR_X1 port map( D => n6069, CK => Clk, RN => 
                           n3879, Q => net113845, QN => n668);
   pc_target_reg_13_26_inst : DFFR_X1 port map( D => n6068, CK => Clk, RN => 
                           n3879, Q => net113844, QN => n667);
   pc_target_reg_13_28_inst : DFFR_X1 port map( D => n6067, CK => Clk, RN => 
                           n3879, Q => net113843, QN => n666);
   pc_target_reg_14_31_inst : DFFR_X1 port map( D => n6065, CK => Clk, RN => 
                           n3864, Q => pc_target_14_31_port, QN => net113842);
   pc_target_reg_14_29_inst : DFFR_X1 port map( D => n6064, CK => Clk, RN => 
                           n3879, Q => pc_target_14_29_port, QN => net113841);
   pc_target_reg_14_27_inst : DFFR_X1 port map( D => n6063, CK => Clk, RN => 
                           n3879, Q => pc_target_14_27_port, QN => net113840);
   pc_target_reg_14_25_inst : DFFR_X1 port map( D => n6062, CK => Clk, RN => 
                           n3879, Q => pc_target_14_25_port, QN => net113839);
   pc_target_reg_14_23_inst : DFFR_X1 port map( D => n6061, CK => Clk, RN => 
                           n3879, Q => pc_target_14_23_port, QN => net113838);
   pc_target_reg_14_21_inst : DFFR_X1 port map( D => n6060, CK => Clk, RN => 
                           n3879, Q => pc_target_14_21_port, QN => net113837);
   pc_target_reg_14_19_inst : DFFR_X1 port map( D => n6059, CK => Clk, RN => 
                           n3879, Q => pc_target_14_19_port, QN => net113836);
   pc_target_reg_14_17_inst : DFFR_X1 port map( D => n6058, CK => Clk, RN => 
                           n3879, Q => pc_target_14_17_port, QN => net113835);
   pc_target_reg_14_15_inst : DFFR_X1 port map( D => n6057, CK => Clk, RN => 
                           n3880, Q => pc_target_14_15_port, QN => net113834);
   pc_target_reg_14_13_inst : DFFR_X1 port map( D => n6056, CK => Clk, RN => 
                           n3840, Q => pc_target_14_13_port, QN => net113833);
   pc_target_reg_14_11_inst : DFFR_X1 port map( D => n6055, CK => Clk, RN => 
                           n3836, Q => pc_target_14_11_port, QN => net113832);
   pc_target_reg_14_9_inst : DFFR_X1 port map( D => n6054, CK => Clk, RN => 
                           n3832, Q => pc_target_14_9_port, QN => net113831);
   pc_target_reg_14_7_inst : DFFR_X1 port map( D => n6053, CK => Clk, RN => 
                           n3832, Q => pc_target_14_7_port, QN => net113830);
   pc_target_reg_14_5_inst : DFFR_X1 port map( D => n6052, CK => Clk, RN => 
                           n3832, Q => pc_target_14_5_port, QN => net113829);
   pc_target_reg_14_3_inst : DFFR_X1 port map( D => n6051, CK => Clk, RN => 
                           n3832, Q => pc_target_14_3_port, QN => net113828);
   pc_target_reg_14_1_inst : DFFR_X1 port map( D => n6050, CK => Clk, RN => 
                           n3832, Q => pc_target_14_1_port, QN => net113827);
   pc_target_reg_14_0_inst : DFFR_X1 port map( D => n6049, CK => Clk, RN => 
                           n3832, Q => pc_target_14_0_port, QN => net113826);
   pc_target_reg_14_2_inst : DFFR_X1 port map( D => n6048, CK => Clk, RN => 
                           n3832, Q => pc_target_14_2_port, QN => net113825);
   pc_target_reg_14_4_inst : DFFR_X1 port map( D => n6047, CK => Clk, RN => 
                           n3832, Q => pc_target_14_4_port, QN => net113824);
   pc_target_reg_14_6_inst : DFFR_X1 port map( D => n6046, CK => Clk, RN => 
                           n3832, Q => pc_target_14_6_port, QN => net113823);
   pc_target_reg_14_8_inst : DFFR_X1 port map( D => n6045, CK => Clk, RN => 
                           n3833, Q => pc_target_14_8_port, QN => net113822);
   pc_target_reg_14_10_inst : DFFR_X1 port map( D => n6044, CK => Clk, RN => 
                           n3833, Q => pc_target_14_10_port, QN => net113821);
   pc_target_reg_14_12_inst : DFFR_X1 port map( D => n6043, CK => Clk, RN => 
                           n3833, Q => pc_target_14_12_port, QN => net113820);
   pc_target_reg_14_14_inst : DFFR_X1 port map( D => n6042, CK => Clk, RN => 
                           n3833, Q => pc_target_14_14_port, QN => net113819);
   pc_target_reg_14_16_inst : DFFR_X1 port map( D => n6041, CK => Clk, RN => 
                           n3833, Q => pc_target_14_16_port, QN => net113818);
   pc_target_reg_14_18_inst : DFFR_X1 port map( D => n6040, CK => Clk, RN => 
                           n3833, Q => pc_target_14_18_port, QN => net113817);
   pc_target_reg_14_20_inst : DFFR_X1 port map( D => n6039, CK => Clk, RN => 
                           n3833, Q => pc_target_14_20_port, QN => net113816);
   pc_target_reg_14_22_inst : DFFR_X1 port map( D => n6038, CK => Clk, RN => 
                           n3833, Q => pc_target_14_22_port, QN => net113815);
   pc_target_reg_14_24_inst : DFFR_X1 port map( D => n6037, CK => Clk, RN => 
                           n3833, Q => pc_target_14_24_port, QN => net113814);
   pc_target_reg_14_26_inst : DFFR_X1 port map( D => n6036, CK => Clk, RN => 
                           n3833, Q => pc_target_14_26_port, QN => net113813);
   pc_target_reg_14_28_inst : DFFR_X1 port map( D => n6035, CK => Clk, RN => 
                           n3833, Q => pc_target_14_28_port, QN => net113812);
   pc_target_reg_14_30_inst : DFFR_X1 port map( D => n6034, CK => Clk, RN => 
                           n3834, Q => pc_target_14_30_port, QN => net113811);
   pc_target_reg_15_31_inst : DFFR_X1 port map( D => n6033, CK => Clk, RN => 
                           n3864, Q => pc_target_15_31_port, QN => net113810);
   pc_target_reg_15_29_inst : DFFR_X1 port map( D => n6032, CK => Clk, RN => 
                           n3833, Q => pc_target_15_29_port, QN => net113809);
   pc_target_reg_15_27_inst : DFFR_X1 port map( D => n6031, CK => Clk, RN => 
                           n3833, Q => pc_target_15_27_port, QN => net113808);
   pc_target_reg_15_25_inst : DFFR_X1 port map( D => n6030, CK => Clk, RN => 
                           n3833, Q => pc_target_15_25_port, QN => net113807);
   pc_target_reg_15_23_inst : DFFR_X1 port map( D => n6029, CK => Clk, RN => 
                           n3833, Q => pc_target_15_23_port, QN => net113806);
   pc_target_reg_15_21_inst : DFFR_X1 port map( D => n6028, CK => Clk, RN => 
                           n3834, Q => pc_target_15_21_port, QN => net113805);
   pc_target_reg_15_19_inst : DFFR_X1 port map( D => n6027, CK => Clk, RN => 
                           n3834, Q => pc_target_15_19_port, QN => net113804);
   pc_target_reg_15_17_inst : DFFR_X1 port map( D => n6026, CK => Clk, RN => 
                           n3834, Q => pc_target_15_17_port, QN => net113803);
   pc_target_reg_15_15_inst : DFFR_X1 port map( D => n6025, CK => Clk, RN => 
                           n3834, Q => pc_target_15_15_port, QN => net113802);
   pc_target_reg_15_13_inst : DFFR_X1 port map( D => n6024, CK => Clk, RN => 
                           n3834, Q => pc_target_15_13_port, QN => net113801);
   pc_target_reg_15_11_inst : DFFR_X1 port map( D => n6023, CK => Clk, RN => 
                           n3834, Q => pc_target_15_11_port, QN => net113800);
   pc_target_reg_15_7_inst : DFFR_X1 port map( D => n6021, CK => Clk, RN => 
                           n3838, Q => pc_target_15_7_port, QN => net113799);
   pc_target_reg_15_12_inst : DFFR_X1 port map( D => n6011, CK => Clk, RN => 
                           n3838, Q => pc_target_15_12_port, QN => net113798);
   pc_target_reg_15_14_inst : DFFR_X1 port map( D => n6010, CK => Clk, RN => 
                           n3838, Q => pc_target_15_14_port, QN => net113797);
   pc_target_reg_15_16_inst : DFFR_X1 port map( D => n6009, CK => Clk, RN => 
                           n3834, Q => pc_target_15_16_port, QN => net113796);
   pc_target_reg_15_18_inst : DFFR_X1 port map( D => n6008, CK => Clk, RN => 
                           n3834, Q => pc_target_15_18_port, QN => net113795);
   pc_target_reg_15_20_inst : DFFR_X1 port map( D => n6007, CK => Clk, RN => 
                           n3834, Q => pc_target_15_20_port, QN => net113794);
   pc_target_reg_15_22_inst : DFFR_X1 port map( D => n6006, CK => Clk, RN => 
                           n3834, Q => pc_target_15_22_port, QN => net113793);
   pc_target_reg_15_24_inst : DFFR_X1 port map( D => n6005, CK => Clk, RN => 
                           n3834, Q => pc_target_15_24_port, QN => net113792);
   pc_target_reg_15_26_inst : DFFR_X1 port map( D => n6004, CK => Clk, RN => 
                           n3834, Q => pc_target_15_26_port, QN => net113791);
   pc_target_reg_15_28_inst : DFFR_X1 port map( D => n6003, CK => Clk, RN => 
                           n3834, Q => pc_target_15_28_port, QN => net113790);
   pc_target_reg_15_30_inst : DFFR_X1 port map( D => n6002, CK => Clk, RN => 
                           n3834, Q => pc_target_15_30_port, QN => net113789);
   pc_target_reg_16_31_inst : DFFR_X1 port map( D => n6001, CK => Clk, RN => 
                           n3865, Q => net113788, QN => n591);
   pc_target_reg_16_29_inst : DFFR_X1 port map( D => n6000, CK => Clk, RN => 
                           n3835, Q => net113787, QN => n590);
   pc_target_reg_16_27_inst : DFFR_X1 port map( D => n5999, CK => Clk, RN => 
                           n3835, Q => net113786, QN => n589);
   pc_target_reg_16_25_inst : DFFR_X1 port map( D => n5998, CK => Clk, RN => 
                           n3835, Q => net113785, QN => n588);
   pc_target_reg_16_23_inst : DFFR_X1 port map( D => n5997, CK => Clk, RN => 
                           n3835, Q => net113784, QN => n587);
   pc_target_reg_16_21_inst : DFFR_X1 port map( D => n5996, CK => Clk, RN => 
                           n3835, Q => net113783, QN => n586);
   pc_target_reg_16_19_inst : DFFR_X1 port map( D => n5995, CK => Clk, RN => 
                           n3835, Q => net113782, QN => n585);
   pc_target_reg_16_17_inst : DFFR_X1 port map( D => n5994, CK => Clk, RN => 
                           n3835, Q => net113781, QN => n584);
   pc_target_reg_16_15_inst : DFFR_X1 port map( D => n5993, CK => Clk, RN => 
                           n3835, Q => net113780, QN => n583);
   pc_target_reg_16_13_inst : DFFR_X1 port map( D => n5992, CK => Clk, RN => 
                           n3835, Q => net113779, QN => n582);
   pc_target_reg_16_11_inst : DFFR_X1 port map( D => n5991, CK => Clk, RN => 
                           n3835, Q => net113778, QN => n581);
   pc_target_reg_16_9_inst : DFFR_X1 port map( D => n5990, CK => Clk, RN => 
                           n3835, Q => net113777, QN => n580);
   pc_target_reg_16_7_inst : DFFR_X1 port map( D => n5989, CK => Clk, RN => 
                           n3835, Q => net113776, QN => n579);
   pc_target_reg_16_5_inst : DFFR_X1 port map( D => n5988, CK => Clk, RN => 
                           n3835, Q => net113775, QN => n578);
   pc_target_reg_16_3_inst : DFFR_X1 port map( D => n5987, CK => Clk, RN => 
                           n3835, Q => net113774, QN => n577);
   pc_target_reg_16_1_inst : DFFR_X1 port map( D => n5986, CK => Clk, RN => 
                           n3835, Q => net113773, QN => n576);
   pc_target_reg_16_0_inst : DFFR_X1 port map( D => n5985, CK => Clk, RN => 
                           n3836, Q => net113772, QN => n575);
   pc_target_reg_16_2_inst : DFFR_X1 port map( D => n5984, CK => Clk, RN => 
                           n3836, Q => net113771, QN => n574);
   pc_target_reg_16_4_inst : DFFR_X1 port map( D => n5983, CK => Clk, RN => 
                           n3836, Q => net113770, QN => n573);
   pc_target_reg_16_6_inst : DFFR_X1 port map( D => n5982, CK => Clk, RN => 
                           n3836, Q => net113769, QN => n572);
   pc_target_reg_16_8_inst : DFFR_X1 port map( D => n5981, CK => Clk, RN => 
                           n3836, Q => net113768, QN => n571);
   pc_target_reg_16_10_inst : DFFR_X1 port map( D => n5980, CK => Clk, RN => 
                           n3836, Q => net113767, QN => n570);
   pc_target_reg_16_12_inst : DFFR_X1 port map( D => n5979, CK => Clk, RN => 
                           n3836, Q => net113766, QN => n569);
   pc_target_reg_16_14_inst : DFFR_X1 port map( D => n5978, CK => Clk, RN => 
                           n3836, Q => net113765, QN => n568);
   pc_target_reg_16_16_inst : DFFR_X1 port map( D => n5977, CK => Clk, RN => 
                           n3836, Q => net113764, QN => n567);
   pc_target_reg_16_18_inst : DFFR_X1 port map( D => n5976, CK => Clk, RN => 
                           n3836, Q => net113763, QN => n566);
   pc_target_reg_16_20_inst : DFFR_X1 port map( D => n5975, CK => Clk, RN => 
                           n3836, Q => net113762, QN => n565);
   pc_target_reg_16_24_inst : DFFR_X1 port map( D => n5973, CK => Clk, RN => 
                           n3836, Q => net113760, QN => n563);
   pc_target_reg_16_26_inst : DFFR_X1 port map( D => n5972, CK => Clk, RN => 
                           n3836, Q => net113759, QN => n562);
   pc_target_reg_16_28_inst : DFFR_X1 port map( D => n5971, CK => Clk, RN => 
                           n3837, Q => net113758, QN => n561);
   pc_target_reg_17_31_inst : DFFR_X1 port map( D => n5969, CK => Clk, RN => 
                           n3865, Q => net113757, QN => n557);
   pc_target_reg_17_29_inst : DFFR_X1 port map( D => n5968, CK => Clk, RN => 
                           n3837, Q => net113756, QN => n556);
   pc_target_reg_17_27_inst : DFFR_X1 port map( D => n5967, CK => Clk, RN => 
                           n3837, Q => net113755, QN => n555);
   pc_target_reg_17_25_inst : DFFR_X1 port map( D => n5966, CK => Clk, RN => 
                           n3837, Q => net113754, QN => n554);
   pc_target_reg_17_23_inst : DFFR_X1 port map( D => n5965, CK => Clk, RN => 
                           n3837, Q => net113753, QN => n553);
   pc_target_reg_17_21_inst : DFFR_X1 port map( D => n5964, CK => Clk, RN => 
                           n3837, Q => net113752, QN => n552);
   pc_target_reg_17_19_inst : DFFR_X1 port map( D => n5963, CK => Clk, RN => 
                           n3837, Q => net113751, QN => n551);
   pc_target_reg_17_17_inst : DFFR_X1 port map( D => n5962, CK => Clk, RN => 
                           n3837, Q => net113750, QN => n550);
   pc_target_reg_17_15_inst : DFFR_X1 port map( D => n5961, CK => Clk, RN => 
                           n3837, Q => net113749, QN => n549);
   pc_target_reg_17_13_inst : DFFR_X1 port map( D => n5960, CK => Clk, RN => 
                           n3837, Q => net113748, QN => n548);
   pc_target_reg_17_11_inst : DFFR_X1 port map( D => n5959, CK => Clk, RN => 
                           n3837, Q => net113747, QN => n547);
   pc_target_reg_17_9_inst : DFFR_X1 port map( D => n5958, CK => Clk, RN => 
                           n3837, Q => net113746, QN => n546);
   pc_target_reg_17_7_inst : DFFR_X1 port map( D => n5957, CK => Clk, RN => 
                           n3837, Q => net113745, QN => n545);
   pc_target_reg_17_3_inst : DFFR_X1 port map( D => n5955, CK => Clk, RN => 
                           n3837, Q => net113744, QN => n543);
   pc_target_reg_17_1_inst : DFFR_X1 port map( D => n5954, CK => Clk, RN => 
                           n3837, Q => n_1086, QN => n542);
   pc_target_reg_17_0_inst : DFFR_X1 port map( D => n5953, CK => Clk, RN => 
                           n3838, Q => n_1087, QN => n541);
   pc_target_reg_17_2_inst : DFFR_X1 port map( D => n5952, CK => Clk, RN => 
                           n3838, Q => net113741, QN => n540);
   pc_target_reg_17_6_inst : DFFR_X1 port map( D => n5950, CK => Clk, RN => 
                           n3838, Q => n_1088, QN => n538);
   pc_target_reg_17_8_inst : DFFR_X1 port map( D => n5949, CK => Clk, RN => 
                           n3838, Q => net113739, QN => n537);
   pc_target_reg_17_10_inst : DFFR_X1 port map( D => n5948, CK => Clk, RN => 
                           n3838, Q => net113738, QN => n536);
   pc_target_reg_17_12_inst : DFFR_X1 port map( D => n5947, CK => Clk, RN => 
                           n3838, Q => net113737, QN => n535);
   pc_target_reg_17_14_inst : DFFR_X1 port map( D => n5946, CK => Clk, RN => 
                           n3838, Q => net113736, QN => n534);
   pc_target_reg_17_16_inst : DFFR_X1 port map( D => n5945, CK => Clk, RN => 
                           n3838, Q => net113735, QN => n533);
   pc_target_reg_17_18_inst : DFFR_X1 port map( D => n5944, CK => Clk, RN => 
                           n3838, Q => net113734, QN => n532);
   pc_target_reg_17_20_inst : DFFR_X1 port map( D => n5943, CK => Clk, RN => 
                           n3838, Q => net113733, QN => n531);
   pc_target_reg_17_22_inst : DFFR_X1 port map( D => n5942, CK => Clk, RN => 
                           n3838, Q => net113732, QN => n530);
   pc_target_reg_17_24_inst : DFFR_X1 port map( D => n5941, CK => Clk, RN => 
                           n3838, Q => net113731, QN => n529);
   pc_target_reg_17_26_inst : DFFR_X1 port map( D => n5940, CK => Clk, RN => 
                           n3839, Q => net113730, QN => n528);
   pc_target_reg_17_28_inst : DFFR_X1 port map( D => n5939, CK => Clk, RN => 
                           n3839, Q => net113729, QN => n527);
   pc_target_reg_18_31_inst : DFFR_X1 port map( D => n5937, CK => Clk, RN => 
                           n3864, Q => pc_target_18_31_port, QN => net113728);
   pc_target_reg_18_29_inst : DFFR_X1 port map( D => n5936, CK => Clk, RN => 
                           n3839, Q => pc_target_18_29_port, QN => net113727);
   pc_target_reg_18_27_inst : DFFR_X1 port map( D => n5935, CK => Clk, RN => 
                           n3839, Q => pc_target_18_27_port, QN => net113726);
   pc_target_reg_18_25_inst : DFFR_X1 port map( D => n5934, CK => Clk, RN => 
                           n3839, Q => pc_target_18_25_port, QN => net113725);
   pc_target_reg_18_23_inst : DFFR_X1 port map( D => n5933, CK => Clk, RN => 
                           n3839, Q => pc_target_18_23_port, QN => net113724);
   pc_target_reg_18_21_inst : DFFR_X1 port map( D => n5932, CK => Clk, RN => 
                           n3839, Q => pc_target_18_21_port, QN => net113723);
   pc_target_reg_18_19_inst : DFFR_X1 port map( D => n5931, CK => Clk, RN => 
                           n3839, Q => pc_target_18_19_port, QN => net113722);
   pc_target_reg_18_17_inst : DFFR_X1 port map( D => n5930, CK => Clk, RN => 
                           n3839, Q => pc_target_18_17_port, QN => net113721);
   pc_target_reg_18_15_inst : DFFR_X1 port map( D => n5929, CK => Clk, RN => 
                           n3839, Q => pc_target_18_15_port, QN => net113720);
   pc_target_reg_18_13_inst : DFFR_X1 port map( D => n5928, CK => Clk, RN => 
                           n3839, Q => pc_target_18_13_port, QN => net113719);
   pc_target_reg_18_11_inst : DFFR_X1 port map( D => n5927, CK => Clk, RN => 
                           n3839, Q => pc_target_18_11_port, QN => net113718);
   pc_target_reg_18_9_inst : DFFR_X1 port map( D => n5926, CK => Clk, RN => 
                           n3839, Q => pc_target_18_9_port, QN => net113717);
   pc_target_reg_18_7_inst : DFFR_X1 port map( D => n5925, CK => Clk, RN => 
                           n3839, Q => pc_target_18_7_port, QN => net113716);
   pc_target_reg_18_5_inst : DFFR_X1 port map( D => n5924, CK => Clk, RN => 
                           n3839, Q => pc_target_18_5_port, QN => net113715);
   pc_target_reg_18_3_inst : DFFR_X1 port map( D => n5923, CK => Clk, RN => 
                           n3840, Q => pc_target_18_3_port, QN => net113714);
   pc_target_reg_18_1_inst : DFFR_X1 port map( D => n5922, CK => Clk, RN => 
                           n3829, Q => pc_target_18_1_port, QN => net113713);
   pc_target_reg_18_0_inst : DFFR_X1 port map( D => n5921, CK => Clk, RN => 
                           n3826, Q => pc_target_18_0_port, QN => net113712);
   pc_target_reg_18_2_inst : DFFR_X1 port map( D => n5920, CK => Clk, RN => 
                           n3828, Q => pc_target_18_2_port, QN => net113711);
   pc_target_reg_18_4_inst : DFFR_X1 port map( D => n5919, CK => Clk, RN => 
                           n3826, Q => pc_target_18_4_port, QN => net113710);
   pc_target_reg_18_6_inst : DFFR_X1 port map( D => n5918, CK => Clk, RN => 
                           n3826, Q => pc_target_18_6_port, QN => net113709);
   pc_target_reg_18_8_inst : DFFR_X1 port map( D => n5917, CK => Clk, RN => 
                           n3826, Q => pc_target_18_8_port, QN => net113708);
   pc_target_reg_18_10_inst : DFFR_X1 port map( D => n5916, CK => Clk, RN => 
                           n3827, Q => pc_target_18_10_port, QN => net113707);
   pc_target_reg_18_12_inst : DFFR_X1 port map( D => n5915, CK => Clk, RN => 
                           n3826, Q => pc_target_18_12_port, QN => net113706);
   pc_target_reg_18_14_inst : DFFR_X1 port map( D => n5914, CK => Clk, RN => 
                           n3828, Q => pc_target_18_14_port, QN => net113705);
   pc_target_reg_18_16_inst : DFFR_X1 port map( D => n5913, CK => Clk, RN => 
                           n3826, Q => pc_target_18_16_port, QN => net113704);
   pc_target_reg_18_18_inst : DFFR_X1 port map( D => n5912, CK => Clk, RN => 
                           n3828, Q => pc_target_18_18_port, QN => net113703);
   pc_target_reg_18_20_inst : DFFR_X1 port map( D => n5911, CK => Clk, RN => 
                           n3828, Q => pc_target_18_20_port, QN => net113702);
   pc_target_reg_18_22_inst : DFFR_X1 port map( D => n5910, CK => Clk, RN => 
                           n3828, Q => pc_target_18_22_port, QN => net113701);
   pc_target_reg_18_24_inst : DFFR_X1 port map( D => n5909, CK => Clk, RN => 
                           n3827, Q => pc_target_18_24_port, QN => net113700);
   pc_target_reg_18_26_inst : DFFR_X1 port map( D => n5908, CK => Clk, RN => 
                           n3827, Q => pc_target_18_26_port, QN => net113699);
   pc_target_reg_18_28_inst : DFFR_X1 port map( D => n5907, CK => Clk, RN => 
                           n3828, Q => pc_target_18_28_port, QN => net113698);
   pc_target_reg_18_30_inst : DFFR_X1 port map( D => n5906, CK => Clk, RN => 
                           n3827, Q => pc_target_18_30_port, QN => net113697);
   pc_target_reg_19_31_inst : DFFR_X1 port map( D => n5905, CK => Clk, RN => 
                           n3864, Q => pc_target_19_31_port, QN => net113696);
   pc_target_reg_19_29_inst : DFFR_X1 port map( D => n5904, CK => Clk, RN => 
                           n3826, Q => pc_target_19_29_port, QN => net113695);
   pc_target_reg_19_27_inst : DFFR_X1 port map( D => n5903, CK => Clk, RN => 
                           n3828, Q => pc_target_19_27_port, QN => net113694);
   pc_target_reg_19_25_inst : DFFR_X1 port map( D => n5902, CK => Clk, RN => 
                           n3827, Q => pc_target_19_25_port, QN => net113693);
   pc_target_reg_19_23_inst : DFFR_X1 port map( D => n5901, CK => Clk, RN => 
                           n3827, Q => pc_target_19_23_port, QN => net113692);
   pc_target_reg_19_21_inst : DFFR_X1 port map( D => n5900, CK => Clk, RN => 
                           n3827, Q => pc_target_19_21_port, QN => net113691);
   pc_target_reg_19_19_inst : DFFR_X1 port map( D => n5899, CK => Clk, RN => 
                           n3829, Q => pc_target_19_19_port, QN => net113690);
   pc_target_reg_19_17_inst : DFFR_X1 port map( D => n5898, CK => Clk, RN => 
                           n3827, Q => pc_target_19_17_port, QN => net113689);
   pc_target_reg_19_15_inst : DFFR_X1 port map( D => n5897, CK => Clk, RN => 
                           n3827, Q => pc_target_19_15_port, QN => net113688);
   pc_target_reg_19_13_inst : DFFR_X1 port map( D => n5896, CK => Clk, RN => 
                           n3828, Q => pc_target_19_13_port, QN => net113687);
   pc_target_reg_19_11_inst : DFFR_X1 port map( D => n5895, CK => Clk, RN => 
                           n3827, Q => pc_target_19_11_port, QN => net113686);
   pc_target_reg_19_9_inst : DFFR_X1 port map( D => n5894, CK => Clk, RN => 
                           n3827, Q => pc_target_19_9_port, QN => net113685);
   pc_target_reg_19_7_inst : DFFR_X1 port map( D => n5893, CK => Clk, RN => 
                           n3828, Q => pc_target_19_7_port, QN => net113684);
   pc_target_reg_19_5_inst : DFFR_X1 port map( D => n5892, CK => Clk, RN => 
                           n3827, Q => pc_target_19_5_port, QN => net113683);
   pc_target_reg_19_3_inst : DFFR_X1 port map( D => n5891, CK => Clk, RN => 
                           n3827, Q => pc_target_19_3_port, QN => net113682);
   pc_target_reg_19_1_inst : DFFR_X1 port map( D => n5890, CK => Clk, RN => 
                           n3828, Q => pc_target_19_1_port, QN => net113681);
   pc_target_reg_19_0_inst : DFFR_X1 port map( D => n5889, CK => Clk, RN => 
                           n3828, Q => pc_target_19_0_port, QN => net113680);
   pc_target_reg_19_2_inst : DFFR_X1 port map( D => n5888, CK => Clk, RN => 
                           n3827, Q => pc_target_19_2_port, QN => net113679);
   pc_target_reg_19_4_inst : DFFR_X1 port map( D => n5887, CK => Clk, RN => 
                           n3829, Q => pc_target_19_4_port, QN => net113678);
   pc_target_reg_19_6_inst : DFFR_X1 port map( D => n5886, CK => Clk, RN => 
                           n3828, Q => pc_target_19_6_port, QN => net113677);
   pc_target_reg_19_8_inst : DFFR_X1 port map( D => n5885, CK => Clk, RN => 
                           n3828, Q => pc_target_19_8_port, QN => net113676);
   pc_target_reg_19_10_inst : DFFR_X1 port map( D => n5884, CK => Clk, RN => 
                           n3828, Q => pc_target_19_10_port, QN => net113675);
   pc_target_reg_19_12_inst : DFFR_X1 port map( D => n5883, CK => Clk, RN => 
                           n3828, Q => pc_target_19_12_port, QN => net113674);
   pc_target_reg_19_14_inst : DFFR_X1 port map( D => n5882, CK => Clk, RN => 
                           n3829, Q => pc_target_19_14_port, QN => net113673);
   pc_target_reg_19_16_inst : DFFR_X1 port map( D => n5881, CK => Clk, RN => 
                           n3829, Q => pc_target_19_16_port, QN => net113672);
   pc_target_reg_19_18_inst : DFFR_X1 port map( D => n5880, CK => Clk, RN => 
                           n3829, Q => pc_target_19_18_port, QN => net113671);
   pc_target_reg_19_20_inst : DFFR_X1 port map( D => n5879, CK => Clk, RN => 
                           n3829, Q => pc_target_19_20_port, QN => net113670);
   pc_target_reg_19_22_inst : DFFR_X1 port map( D => n5878, CK => Clk, RN => 
                           n3829, Q => pc_target_19_22_port, QN => net113669);
   pc_target_reg_19_24_inst : DFFR_X1 port map( D => n5877, CK => Clk, RN => 
                           n3829, Q => pc_target_19_24_port, QN => net113668);
   pc_target_reg_19_26_inst : DFFR_X1 port map( D => n5876, CK => Clk, RN => 
                           n3829, Q => pc_target_19_26_port, QN => net113667);
   pc_target_reg_19_28_inst : DFFR_X1 port map( D => n5875, CK => Clk, RN => 
                           n3829, Q => pc_target_19_28_port, QN => net113666);
   pc_target_reg_19_30_inst : DFFR_X1 port map( D => n5874, CK => Clk, RN => 
                           n3829, Q => pc_target_19_30_port, QN => net113665);
   pc_target_reg_20_31_inst : DFFR_X1 port map( D => n5873, CK => Clk, RN => 
                           n3864, Q => pc_target_20_31_port, QN => net113664);
   pc_target_reg_20_29_inst : DFFR_X1 port map( D => n5872, CK => Clk, RN => 
                           n3880, Q => pc_target_20_29_port, QN => net113663);
   pc_target_reg_20_27_inst : DFFR_X1 port map( D => n5871, CK => Clk, RN => 
                           n3880, Q => pc_target_20_27_port, QN => net113662);
   pc_target_reg_20_25_inst : DFFR_X1 port map( D => n5870, CK => Clk, RN => 
                           n3880, Q => pc_target_20_25_port, QN => net113661);
   pc_target_reg_20_23_inst : DFFR_X1 port map( D => n5869, CK => Clk, RN => 
                           n3880, Q => pc_target_20_23_port, QN => net113660);
   pc_target_reg_20_21_inst : DFFR_X1 port map( D => n5868, CK => Clk, RN => 
                           n3880, Q => pc_target_20_21_port, QN => net113659);
   pc_target_reg_20_19_inst : DFFR_X1 port map( D => n5867, CK => Clk, RN => 
                           n3880, Q => pc_target_20_19_port, QN => net113658);
   pc_target_reg_20_17_inst : DFFR_X1 port map( D => n5866, CK => Clk, RN => 
                           n3880, Q => pc_target_20_17_port, QN => net113657);
   pc_target_reg_20_15_inst : DFFR_X1 port map( D => n5865, CK => Clk, RN => 
                           n3880, Q => pc_target_20_15_port, QN => net113656);
   pc_target_reg_20_13_inst : DFFR_X1 port map( D => n5864, CK => Clk, RN => 
                           n3880, Q => pc_target_20_13_port, QN => net113655);
   pc_target_reg_20_11_inst : DFFR_X1 port map( D => n5863, CK => Clk, RN => 
                           n3880, Q => pc_target_20_11_port, QN => net113654);
   pc_target_reg_20_9_inst : DFFR_X1 port map( D => n5862, CK => Clk, RN => 
                           n3880, Q => pc_target_20_9_port, QN => net113653);
   pc_target_reg_20_7_inst : DFFR_X1 port map( D => n5861, CK => Clk, RN => 
                           n3880, Q => pc_target_20_7_port, QN => net113652);
   pc_target_reg_20_5_inst : DFFR_X1 port map( D => n5860, CK => Clk, RN => 
                           n3881, Q => pc_target_20_5_port, QN => net113651);
   pc_target_reg_20_3_inst : DFFR_X1 port map( D => n5859, CK => Clk, RN => 
                           n3881, Q => pc_target_20_3_port, QN => net113650);
   pc_target_reg_20_1_inst : DFFR_X1 port map( D => n5858, CK => Clk, RN => 
                           n3881, Q => pc_target_20_1_port, QN => net113649);
   pc_target_reg_20_0_inst : DFFR_X1 port map( D => n5857, CK => Clk, RN => 
                           n3881, Q => pc_target_20_0_port, QN => net113648);
   pc_target_reg_20_2_inst : DFFR_X1 port map( D => n5856, CK => Clk, RN => 
                           n3881, Q => pc_target_20_2_port, QN => net113647);
   pc_target_reg_20_4_inst : DFFR_X1 port map( D => n5855, CK => Clk, RN => 
                           n3881, Q => pc_target_20_4_port, QN => net113646);
   pc_target_reg_20_6_inst : DFFR_X1 port map( D => n5854, CK => Clk, RN => 
                           n3881, Q => pc_target_20_6_port, QN => net113645);
   pc_target_reg_20_8_inst : DFFR_X1 port map( D => n5853, CK => Clk, RN => 
                           n3881, Q => pc_target_20_8_port, QN => net113644);
   pc_target_reg_20_10_inst : DFFR_X1 port map( D => n5852, CK => Clk, RN => 
                           n3881, Q => pc_target_20_10_port, QN => net113643);
   pc_target_reg_20_12_inst : DFFR_X1 port map( D => n5851, CK => Clk, RN => 
                           n3881, Q => pc_target_20_12_port, QN => net113642);
   pc_target_reg_20_14_inst : DFFR_X1 port map( D => n5850, CK => Clk, RN => 
                           n3881, Q => pc_target_20_14_port, QN => net113641);
   pc_target_reg_20_16_inst : DFFR_X1 port map( D => n5849, CK => Clk, RN => 
                           n3881, Q => pc_target_20_16_port, QN => net113640);
   pc_target_reg_20_18_inst : DFFR_X1 port map( D => n5848, CK => Clk, RN => 
                           n3881, Q => pc_target_20_18_port, QN => net113639);
   pc_target_reg_20_20_inst : DFFR_X1 port map( D => n5847, CK => Clk, RN => 
                           n3881, Q => pc_target_20_20_port, QN => net113638);
   pc_target_reg_20_22_inst : DFFR_X1 port map( D => n5846, CK => Clk, RN => 
                           n3881, Q => pc_target_20_22_port, QN => net113637);
   pc_target_reg_20_24_inst : DFFR_X1 port map( D => n5845, CK => Clk, RN => 
                           n3882, Q => pc_target_20_24_port, QN => net113636);
   pc_target_reg_20_26_inst : DFFR_X1 port map( D => n5844, CK => Clk, RN => 
                           n3882, Q => pc_target_20_26_port, QN => net113635);
   pc_target_reg_20_28_inst : DFFR_X1 port map( D => n5843, CK => Clk, RN => 
                           n3882, Q => pc_target_20_28_port, QN => net113634);
   pc_target_reg_20_30_inst : DFFR_X1 port map( D => n5842, CK => Clk, RN => 
                           n3882, Q => pc_target_20_30_port, QN => net113633);
   pc_target_reg_21_31_inst : DFFR_X1 port map( D => n5841, CK => Clk, RN => 
                           n3864, Q => pc_target_21_31_port, QN => net113632);
   pc_target_reg_21_29_inst : DFFR_X1 port map( D => n5840, CK => Clk, RN => 
                           n3882, Q => pc_target_21_29_port, QN => net113631);
   pc_target_reg_21_27_inst : DFFR_X1 port map( D => n5839, CK => Clk, RN => 
                           n3882, Q => pc_target_21_27_port, QN => net113630);
   pc_target_reg_21_25_inst : DFFR_X1 port map( D => n5838, CK => Clk, RN => 
                           n3882, Q => pc_target_21_25_port, QN => net113629);
   pc_target_reg_21_23_inst : DFFR_X1 port map( D => n5837, CK => Clk, RN => 
                           n3882, Q => pc_target_21_23_port, QN => net113628);
   pc_target_reg_21_21_inst : DFFR_X1 port map( D => n5836, CK => Clk, RN => 
                           n3882, Q => pc_target_21_21_port, QN => net113627);
   pc_target_reg_21_19_inst : DFFR_X1 port map( D => n5835, CK => Clk, RN => 
                           n3882, Q => pc_target_21_19_port, QN => net113626);
   pc_target_reg_21_17_inst : DFFR_X1 port map( D => n5834, CK => Clk, RN => 
                           n3882, Q => pc_target_21_17_port, QN => net113625);
   pc_target_reg_21_15_inst : DFFR_X1 port map( D => n5833, CK => Clk, RN => 
                           n3882, Q => pc_target_21_15_port, QN => net113624);
   pc_target_reg_21_13_inst : DFFR_X1 port map( D => n5832, CK => Clk, RN => 
                           n3882, Q => pc_target_21_13_port, QN => net113623);
   pc_target_reg_21_11_inst : DFFR_X1 port map( D => n5831, CK => Clk, RN => 
                           n3882, Q => pc_target_21_11_port, QN => net113622);
   pc_target_reg_21_7_inst : DFFR_X1 port map( D => n5829, CK => Clk, RN => 
                           n3882, Q => pc_target_21_7_port, QN => net113621);
   pc_target_reg_21_3_inst : DFFR_X1 port map( D => n5827, CK => Clk, RN => 
                           n3883, Q => pc_target_21_3_port, QN => net113620);
   pc_target_reg_21_1_inst : DFFR_X1 port map( D => n5826, CK => Clk, RN => 
                           n3883, Q => pc_target_21_1_port, QN => net113619);
   pc_target_reg_21_0_inst : DFFR_X1 port map( D => n5825, CK => Clk, RN => 
                           n3883, Q => pc_target_21_0_port, QN => net113618);
   pc_target_reg_21_2_inst : DFFR_X1 port map( D => n5824, CK => Clk, RN => 
                           n3883, Q => pc_target_21_2_port, QN => net113617);
   pc_target_reg_21_12_inst : DFFR_X1 port map( D => n5819, CK => Clk, RN => 
                           n3883, Q => pc_target_21_12_port, QN => net113616);
   pc_target_reg_21_14_inst : DFFR_X1 port map( D => n5818, CK => Clk, RN => 
                           n3883, Q => pc_target_21_14_port, QN => net113615);
   pc_target_reg_21_16_inst : DFFR_X1 port map( D => n5817, CK => Clk, RN => 
                           n3883, Q => pc_target_21_16_port, QN => net113614);
   pc_target_reg_21_18_inst : DFFR_X1 port map( D => n5816, CK => Clk, RN => 
                           n3883, Q => pc_target_21_18_port, QN => net113613);
   pc_target_reg_21_20_inst : DFFR_X1 port map( D => n5815, CK => Clk, RN => 
                           n3883, Q => pc_target_21_20_port, QN => net113612);
   pc_target_reg_21_22_inst : DFFR_X1 port map( D => n5814, CK => Clk, RN => 
                           n3883, Q => pc_target_21_22_port, QN => net113611);
   pc_target_reg_21_24_inst : DFFR_X1 port map( D => n5813, CK => Clk, RN => 
                           n3883, Q => pc_target_21_24_port, QN => net113610);
   pc_target_reg_21_26_inst : DFFR_X1 port map( D => n5812, CK => Clk, RN => 
                           n3883, Q => pc_target_21_26_port, QN => net113609);
   pc_target_reg_21_28_inst : DFFR_X1 port map( D => n5811, CK => Clk, RN => 
                           n3883, Q => pc_target_21_28_port, QN => net113608);
   pc_target_reg_21_30_inst : DFFR_X1 port map( D => n5810, CK => Clk, RN => 
                           n3883, Q => pc_target_21_30_port, QN => net113607);
   pc_target_reg_22_31_inst : DFFR_X1 port map( D => n5809, CK => Clk, RN => 
                           n3865, Q => net113606, QN => n385);
   pc_target_reg_22_29_inst : DFFR_X1 port map( D => n5808, CK => Clk, RN => 
                           n3883, Q => net113605, QN => n384);
   pc_target_reg_22_27_inst : DFFR_X1 port map( D => n5807, CK => Clk, RN => 
                           n3884, Q => net113604, QN => n383);
   pc_target_reg_22_25_inst : DFFR_X1 port map( D => n5806, CK => Clk, RN => 
                           n3884, Q => net113603, QN => n382);
   pc_target_reg_22_23_inst : DFFR_X1 port map( D => n5805, CK => Clk, RN => 
                           n3884, Q => net113602, QN => n381);
   pc_target_reg_22_21_inst : DFFR_X1 port map( D => n5804, CK => Clk, RN => 
                           n3884, Q => net113601, QN => n380);
   pc_target_reg_22_19_inst : DFFR_X1 port map( D => n5803, CK => Clk, RN => 
                           n3884, Q => net113600, QN => n379);
   pc_target_reg_22_17_inst : DFFR_X1 port map( D => n5802, CK => Clk, RN => 
                           n3884, Q => net113599, QN => n378);
   pc_target_reg_22_15_inst : DFFR_X1 port map( D => n5801, CK => Clk, RN => 
                           n3884, Q => net113598, QN => n377);
   pc_target_reg_22_13_inst : DFFR_X1 port map( D => n5800, CK => Clk, RN => 
                           n3884, Q => net113597, QN => n376);
   pc_target_reg_22_11_inst : DFFR_X1 port map( D => n5799, CK => Clk, RN => 
                           n3884, Q => net113596, QN => n375);
   pc_target_reg_22_9_inst : DFFR_X1 port map( D => n5798, CK => Clk, RN => 
                           n3884, Q => net113595, QN => n374);
   pc_target_reg_22_7_inst : DFFR_X1 port map( D => n5797, CK => Clk, RN => 
                           n3884, Q => net113594, QN => n373);
   pc_target_reg_22_5_inst : DFFR_X1 port map( D => n5796, CK => Clk, RN => 
                           n3884, Q => n_1089, QN => n372);
   pc_target_reg_22_3_inst : DFFR_X1 port map( D => n5795, CK => Clk, RN => 
                           n3884, Q => net113592, QN => n371);
   pc_target_reg_22_1_inst : DFFR_X1 port map( D => n5794, CK => Clk, RN => 
                           n3884, Q => n_1090, QN => n370);
   pc_target_reg_22_0_inst : DFFR_X1 port map( D => n5793, CK => Clk, RN => 
                           n3885, Q => n_1091, QN => n369);
   pc_target_reg_22_2_inst : DFFR_X1 port map( D => n5792, CK => Clk, RN => 
                           n3885, Q => net113589, QN => n368);
   pc_target_reg_22_4_inst : DFFR_X1 port map( D => n5791, CK => Clk, RN => 
                           n3885, Q => n_1092, QN => n367);
   pc_target_reg_22_6_inst : DFFR_X1 port map( D => n5790, CK => Clk, RN => 
                           n3885, Q => n_1093, QN => n366);
   pc_target_reg_22_8_inst : DFFR_X1 port map( D => n5789, CK => Clk, RN => 
                           n3885, Q => net113586, QN => n365);
   pc_target_reg_22_10_inst : DFFR_X1 port map( D => n5788, CK => Clk, RN => 
                           n3885, Q => net113585, QN => n364);
   pc_target_reg_22_12_inst : DFFR_X1 port map( D => n5787, CK => Clk, RN => 
                           n3885, Q => net113584, QN => n363);
   pc_target_reg_22_14_inst : DFFR_X1 port map( D => n5786, CK => Clk, RN => 
                           n3885, Q => net113583, QN => n362);
   pc_target_reg_22_16_inst : DFFR_X1 port map( D => n5785, CK => Clk, RN => 
                           n3885, Q => net113582, QN => n361);
   pc_target_reg_22_18_inst : DFFR_X1 port map( D => n5784, CK => Clk, RN => 
                           n3885, Q => net113581, QN => n360);
   pc_target_reg_22_20_inst : DFFR_X1 port map( D => n5783, CK => Clk, RN => 
                           n3885, Q => net113580, QN => n359);
   pc_target_reg_22_22_inst : DFFR_X1 port map( D => n5782, CK => Clk, RN => 
                           n3885, Q => net113579, QN => n358);
   pc_target_reg_22_24_inst : DFFR_X1 port map( D => n5781, CK => Clk, RN => 
                           n3886, Q => net113578, QN => n357);
   pc_target_reg_22_26_inst : DFFR_X1 port map( D => n5780, CK => Clk, RN => 
                           n3886, Q => net113577, QN => n356);
   pc_target_reg_22_28_inst : DFFR_X1 port map( D => n5779, CK => Clk, RN => 
                           n3886, Q => net113576, QN => n355);
   pc_target_reg_23_31_inst : DFFR_X1 port map( D => n5777, CK => Clk, RN => 
                           n3865, Q => net113575, QN => n350);
   pc_target_reg_23_29_inst : DFFR_X1 port map( D => n5776, CK => Clk, RN => 
                           n3885, Q => net113574, QN => n349);
   pc_target_reg_23_27_inst : DFFR_X1 port map( D => n5775, CK => Clk, RN => 
                           n3885, Q => net113573, QN => n348);
   pc_target_reg_23_25_inst : DFFR_X1 port map( D => n5774, CK => Clk, RN => 
                           n3885, Q => net113572, QN => n347);
   pc_target_reg_23_23_inst : DFFR_X1 port map( D => n5773, CK => Clk, RN => 
                           n3886, Q => net113571, QN => n346);
   pc_target_reg_23_21_inst : DFFR_X1 port map( D => n5772, CK => Clk, RN => 
                           n3886, Q => net113570, QN => n345);
   pc_target_reg_23_19_inst : DFFR_X1 port map( D => n5771, CK => Clk, RN => 
                           n3886, Q => net113569, QN => n344);
   pc_target_reg_23_17_inst : DFFR_X1 port map( D => n5770, CK => Clk, RN => 
                           n3886, Q => net113568, QN => n343);
   pc_target_reg_23_15_inst : DFFR_X1 port map( D => n5769, CK => Clk, RN => 
                           n3886, Q => net113567, QN => n342);
   pc_target_reg_23_13_inst : DFFR_X1 port map( D => n5768, CK => Clk, RN => 
                           n3886, Q => net113566, QN => n341);
   pc_target_reg_23_11_inst : DFFR_X1 port map( D => n5767, CK => Clk, RN => 
                           n3886, Q => net113565, QN => n340);
   pc_target_reg_23_9_inst : DFFR_X1 port map( D => n5766, CK => Clk, RN => 
                           n3886, Q => net113564, QN => n339);
   pc_target_reg_23_7_inst : DFFR_X1 port map( D => n5765, CK => Clk, RN => 
                           n3886, Q => net113563, QN => n338);
   pc_target_reg_23_5_inst : DFFR_X1 port map( D => n5764, CK => Clk, RN => 
                           n3886, Q => n_1094, QN => n337);
   pc_target_reg_23_3_inst : DFFR_X1 port map( D => n5763, CK => Clk, RN => 
                           n3886, Q => net113561, QN => n336);
   pc_target_reg_23_1_inst : DFFR_X1 port map( D => n5762, CK => Clk, RN => 
                           n3886, Q => n_1095, QN => n335);
   pc_target_reg_23_0_inst : DFFR_X1 port map( D => n5761, CK => Clk, RN => 
                           n3887, Q => n_1096, QN => n334);
   pc_target_reg_23_2_inst : DFFR_X1 port map( D => n5760, CK => Clk, RN => 
                           n3887, Q => net113558, QN => n333);
   pc_target_reg_23_4_inst : DFFR_X1 port map( D => n5759, CK => Clk, RN => 
                           n3887, Q => n_1097, QN => n332);
   pc_target_reg_23_6_inst : DFFR_X1 port map( D => n5758, CK => Clk, RN => 
                           n3887, Q => n_1098, QN => n331);
   pc_target_reg_23_8_inst : DFFR_X1 port map( D => n5757, CK => Clk, RN => 
                           n3887, Q => net113555, QN => n330);
   pc_target_reg_23_10_inst : DFFR_X1 port map( D => n5756, CK => Clk, RN => 
                           n3887, Q => net113554, QN => n329);
   pc_target_reg_23_12_inst : DFFR_X1 port map( D => n5755, CK => Clk, RN => 
                           n3887, Q => net113553, QN => n328);
   pc_target_reg_23_14_inst : DFFR_X1 port map( D => n5754, CK => Clk, RN => 
                           n3887, Q => net113552, QN => n327);
   pc_target_reg_23_16_inst : DFFR_X1 port map( D => n5753, CK => Clk, RN => 
                           n3887, Q => net113551, QN => n326);
   pc_target_reg_23_18_inst : DFFR_X1 port map( D => n5752, CK => Clk, RN => 
                           n3887, Q => net113550, QN => n325);
   pc_target_reg_23_20_inst : DFFR_X1 port map( D => n5751, CK => Clk, RN => 
                           n3887, Q => net113549, QN => n324);
   pc_target_reg_23_22_inst : DFFR_X1 port map( D => n5750, CK => Clk, RN => 
                           n3887, Q => net113548, QN => n323);
   pc_target_reg_23_24_inst : DFFR_X1 port map( D => n5749, CK => Clk, RN => 
                           n3872, Q => net113547, QN => n322);
   pc_target_reg_23_26_inst : DFFR_X1 port map( D => n5748, CK => Clk, RN => 
                           n3872, Q => net113546, QN => n321);
   pc_target_reg_23_28_inst : DFFR_X1 port map( D => n5747, CK => Clk, RN => 
                           n3872, Q => net113545, QN => n320);
   pc_target_reg_24_31_inst : DFFR_X1 port map( D => n5745, CK => Clk, RN => 
                           n3865, Q => net113544, QN => n315);
   pc_target_reg_24_29_inst : DFFR_X1 port map( D => n5744, CK => Clk, RN => 
                           n3887, Q => net113543, QN => n314);
   pc_target_reg_24_27_inst : DFFR_X1 port map( D => n5743, CK => Clk, RN => 
                           n3887, Q => net113542, QN => n313);
   pc_target_reg_24_25_inst : DFFR_X1 port map( D => n5742, CK => Clk, RN => 
                           n3887, Q => net113541, QN => n312);
   pc_target_reg_24_23_inst : DFFR_X1 port map( D => n5741, CK => Clk, RN => 
                           n3888, Q => net113540, QN => n311);
   pc_target_reg_24_21_inst : DFFR_X1 port map( D => n5740, CK => Clk, RN => 
                           n3888, Q => net113539, QN => n310);
   pc_target_reg_24_19_inst : DFFR_X1 port map( D => n5739, CK => Clk, RN => 
                           n3888, Q => net113538, QN => n309);
   pc_target_reg_24_17_inst : DFFR_X1 port map( D => n5738, CK => Clk, RN => 
                           n3875, Q => net113537, QN => n308);
   pc_target_reg_24_15_inst : DFFR_X1 port map( D => n5737, CK => Clk, RN => 
                           n3871, Q => net113536, QN => n307);
   pc_target_reg_24_13_inst : DFFR_X1 port map( D => n5736, CK => Clk, RN => 
                           n3872, Q => net113535, QN => n306);
   pc_target_reg_24_11_inst : DFFR_X1 port map( D => n5735, CK => Clk, RN => 
                           n3872, Q => net113534, QN => n305);
   pc_target_reg_24_9_inst : DFFR_X1 port map( D => n5734, CK => Clk, RN => 
                           n3872, Q => net113533, QN => n304);
   pc_target_reg_24_7_inst : DFFR_X1 port map( D => n5733, CK => Clk, RN => 
                           n3872, Q => net113532, QN => n303);
   pc_target_reg_24_3_inst : DFFR_X1 port map( D => n5731, CK => Clk, RN => 
                           n3872, Q => net113531, QN => n301);
   pc_target_reg_24_1_inst : DFFR_X1 port map( D => n5730, CK => Clk, RN => 
                           n3872, Q => n_1099, QN => n300);
   pc_target_reg_24_0_inst : DFFR_X1 port map( D => n5729, CK => Clk, RN => 
                           n3872, Q => n_1100, QN => n299);
   pc_target_reg_24_2_inst : DFFR_X1 port map( D => n5728, CK => Clk, RN => 
                           n3872, Q => net113528, QN => n298);
   pc_target_reg_24_6_inst : DFFR_X1 port map( D => n5726, CK => Clk, RN => 
                           n3872, Q => n_1101, QN => n296);
   pc_target_reg_24_8_inst : DFFR_X1 port map( D => n5725, CK => Clk, RN => 
                           n3872, Q => net113526, QN => n295);
   pc_target_reg_24_10_inst : DFFR_X1 port map( D => n5724, CK => Clk, RN => 
                           n3872, Q => net113525, QN => n294);
   pc_target_reg_24_12_inst : DFFR_X1 port map( D => n5723, CK => Clk, RN => 
                           n3873, Q => net113524, QN => n293);
   pc_target_reg_24_14_inst : DFFR_X1 port map( D => n5722, CK => Clk, RN => 
                           n3873, Q => net113523, QN => n292);
   pc_target_reg_24_16_inst : DFFR_X1 port map( D => n5721, CK => Clk, RN => 
                           n3873, Q => net113522, QN => n291);
   pc_target_reg_24_18_inst : DFFR_X1 port map( D => n5720, CK => Clk, RN => 
                           n3873, Q => net113521, QN => n290);
   pc_target_reg_24_20_inst : DFFR_X1 port map( D => n5719, CK => Clk, RN => 
                           n3873, Q => net113520, QN => n289);
   pc_target_reg_24_22_inst : DFFR_X1 port map( D => n5718, CK => Clk, RN => 
                           n3873, Q => net113519, QN => n288);
   pc_target_reg_24_24_inst : DFFR_X1 port map( D => n5717, CK => Clk, RN => 
                           n3873, Q => net113518, QN => n287);
   pc_target_reg_24_26_inst : DFFR_X1 port map( D => n5716, CK => Clk, RN => 
                           n3873, Q => net113517, QN => n286);
   pc_target_reg_24_28_inst : DFFR_X1 port map( D => n5715, CK => Clk, RN => 
                           n3873, Q => net113516, QN => n285);
   pc_target_reg_25_31_inst : DFFR_X1 port map( D => n5713, CK => Clk, RN => 
                           n3865, Q => net113515, QN => n281);
   pc_target_reg_25_29_inst : DFFR_X1 port map( D => n5712, CK => Clk, RN => 
                           n3872, Q => net113514, QN => n280);
   pc_target_reg_25_27_inst : DFFR_X1 port map( D => n5711, CK => Clk, RN => 
                           n3873, Q => net113513, QN => n279);
   pc_target_reg_25_25_inst : DFFR_X1 port map( D => n5710, CK => Clk, RN => 
                           n3873, Q => net113512, QN => n278);
   pc_target_reg_25_23_inst : DFFR_X1 port map( D => n5709, CK => Clk, RN => 
                           n3873, Q => net113511, QN => n277);
   pc_target_reg_25_21_inst : DFFR_X1 port map( D => n5708, CK => Clk, RN => 
                           n3873, Q => net113510, QN => n276);
   pc_target_reg_25_19_inst : DFFR_X1 port map( D => n5707, CK => Clk, RN => 
                           n3873, Q => net113509, QN => n275);
   pc_target_reg_25_17_inst : DFFR_X1 port map( D => n5706, CK => Clk, RN => 
                           n3873, Q => net113508, QN => n274);
   pc_target_reg_25_15_inst : DFFR_X1 port map( D => n5705, CK => Clk, RN => 
                           n3874, Q => net113507, QN => n273);
   pc_target_reg_25_13_inst : DFFR_X1 port map( D => n5704, CK => Clk, RN => 
                           n3874, Q => net113506, QN => n272);
   pc_target_reg_25_11_inst : DFFR_X1 port map( D => n5703, CK => Clk, RN => 
                           n3874, Q => net113505, QN => n271);
   pc_target_reg_25_9_inst : DFFR_X1 port map( D => n5702, CK => Clk, RN => 
                           n3874, Q => net113504, QN => n270);
   pc_target_reg_25_7_inst : DFFR_X1 port map( D => n5701, CK => Clk, RN => 
                           n3874, Q => net113503, QN => n269);
   pc_target_reg_25_5_inst : DFFR_X1 port map( D => n5700, CK => Clk, RN => 
                           n3874, Q => net113502, QN => n268);
   pc_target_reg_25_3_inst : DFFR_X1 port map( D => n5699, CK => Clk, RN => 
                           n3874, Q => net113501, QN => n267);
   pc_target_reg_25_1_inst : DFFR_X1 port map( D => n5698, CK => Clk, RN => 
                           n3874, Q => net113500, QN => n266);
   pc_target_reg_25_0_inst : DFFR_X1 port map( D => n5697, CK => Clk, RN => 
                           n3875, Q => net113499, QN => n265);
   pc_target_reg_25_2_inst : DFFR_X1 port map( D => n5696, CK => Clk, RN => 
                           n3874, Q => net113498, QN => n264);
   pc_target_reg_25_4_inst : DFFR_X1 port map( D => n5695, CK => Clk, RN => 
                           n3874, Q => net113497, QN => n263);
   pc_target_reg_25_6_inst : DFFR_X1 port map( D => n5694, CK => Clk, RN => 
                           n3874, Q => net113496, QN => n262);
   pc_target_reg_25_8_inst : DFFR_X1 port map( D => n5693, CK => Clk, RN => 
                           n3874, Q => net113495, QN => n261);
   pc_target_reg_25_10_inst : DFFR_X1 port map( D => n5692, CK => Clk, RN => 
                           n3874, Q => net113494, QN => n260);
   pc_target_reg_25_12_inst : DFFR_X1 port map( D => n5691, CK => Clk, RN => 
                           n3874, Q => net113493, QN => n259);
   pc_target_reg_25_14_inst : DFFR_X1 port map( D => n5690, CK => Clk, RN => 
                           n3874, Q => net113492, QN => n258);
   pc_target_reg_25_16_inst : DFFR_X1 port map( D => n5689, CK => Clk, RN => 
                           n3875, Q => net113491, QN => n257);
   pc_target_reg_25_18_inst : DFFR_X1 port map( D => n5688, CK => Clk, RN => 
                           n3875, Q => net113490, QN => n256);
   pc_target_reg_25_20_inst : DFFR_X1 port map( D => n5687, CK => Clk, RN => 
                           n3875, Q => net113489, QN => n255);
   pc_target_reg_25_22_inst : DFFR_X1 port map( D => n5686, CK => Clk, RN => 
                           n3875, Q => net113488, QN => n254);
   pc_target_reg_25_24_inst : DFFR_X1 port map( D => n5685, CK => Clk, RN => 
                           n3875, Q => net113487, QN => n253);
   pc_target_reg_25_26_inst : DFFR_X1 port map( D => n5684, CK => Clk, RN => 
                           n3875, Q => net113486, QN => n252);
   pc_target_reg_25_28_inst : DFFR_X1 port map( D => n5683, CK => Clk, RN => 
                           n3875, Q => net113485, QN => n251);
   pc_target_reg_26_31_inst : DFFR_X1 port map( D => n5681, CK => Clk, RN => 
                           n3871, Q => pc_target_26_31_port, QN => net113484);
   pc_target_reg_26_29_inst : DFFR_X1 port map( D => n5680, CK => Clk, RN => 
                           n3875, Q => pc_target_26_29_port, QN => net113483);
   pc_target_reg_26_27_inst : DFFR_X1 port map( D => n5679, CK => Clk, RN => 
                           n3875, Q => pc_target_26_27_port, QN => net113482);
   pc_target_reg_26_25_inst : DFFR_X1 port map( D => n5678, CK => Clk, RN => 
                           n3875, Q => pc_target_26_25_port, QN => net113481);
   pc_target_reg_26_23_inst : DFFR_X1 port map( D => n5677, CK => Clk, RN => 
                           n3875, Q => pc_target_26_23_port, QN => net113480);
   pc_target_reg_26_21_inst : DFFR_X1 port map( D => n5676, CK => Clk, RN => 
                           n3875, Q => pc_target_26_21_port, QN => net113479);
   pc_target_reg_26_19_inst : DFFR_X1 port map( D => n5675, CK => Clk, RN => 
                           n3875, Q => pc_target_26_19_port, QN => net113478);
   pc_target_reg_26_17_inst : DFFR_X1 port map( D => n5674, CK => Clk, RN => 
                           n3876, Q => pc_target_26_17_port, QN => net113477);
   pc_target_reg_26_15_inst : DFFR_X1 port map( D => n5673, CK => Clk, RN => 
                           n3876, Q => pc_target_26_15_port, QN => net113476);
   pc_target_reg_26_13_inst : DFFR_X1 port map( D => n5672, CK => Clk, RN => 
                           n3876, Q => pc_target_26_13_port, QN => net113475);
   pc_target_reg_26_11_inst : DFFR_X1 port map( D => n5671, CK => Clk, RN => 
                           n3876, Q => pc_target_26_11_port, QN => net113474);
   pc_target_reg_26_9_inst : DFFR_X1 port map( D => n5670, CK => Clk, RN => 
                           n3876, Q => pc_target_26_9_port, QN => net113473);
   pc_target_reg_26_7_inst : DFFR_X1 port map( D => n5669, CK => Clk, RN => 
                           n3876, Q => pc_target_26_7_port, QN => net113472);
   pc_target_reg_26_5_inst : DFFR_X1 port map( D => n5668, CK => Clk, RN => 
                           n3876, Q => pc_target_26_5_port, QN => net113471);
   pc_target_reg_26_3_inst : DFFR_X1 port map( D => n5667, CK => Clk, RN => 
                           n3876, Q => pc_target_26_3_port, QN => net113470);
   pc_target_reg_26_1_inst : DFFR_X1 port map( D => n5666, CK => Clk, RN => 
                           n3876, Q => pc_target_26_1_port, QN => net113469);
   pc_target_reg_26_0_inst : DFFR_X1 port map( D => n5665, CK => Clk, RN => 
                           n3876, Q => pc_target_26_0_port, QN => net113468);
   pc_target_reg_26_2_inst : DFFR_X1 port map( D => n5664, CK => Clk, RN => 
                           n3876, Q => pc_target_26_2_port, QN => net113467);
   pc_target_reg_26_4_inst : DFFR_X1 port map( D => n5663, CK => Clk, RN => 
                           n3876, Q => pc_target_26_4_port, QN => net113466);
   pc_target_reg_26_6_inst : DFFR_X1 port map( D => n5662, CK => Clk, RN => 
                           n3876, Q => pc_target_26_6_port, QN => net113465);
   pc_target_reg_26_8_inst : DFFR_X1 port map( D => n5661, CK => Clk, RN => 
                           n3876, Q => pc_target_26_8_port, QN => net113464);
   pc_target_reg_26_10_inst : DFFR_X1 port map( D => n5660, CK => Clk, RN => 
                           n3876, Q => pc_target_26_10_port, QN => net113463);
   pc_target_reg_26_12_inst : DFFR_X1 port map( D => n5659, CK => Clk, RN => 
                           n3877, Q => pc_target_26_12_port, QN => net113462);
   pc_target_reg_26_14_inst : DFFR_X1 port map( D => n5658, CK => Clk, RN => 
                           n3877, Q => pc_target_26_14_port, QN => net113461);
   pc_target_reg_26_16_inst : DFFR_X1 port map( D => n5657, CK => Clk, RN => 
                           n3877, Q => pc_target_26_16_port, QN => net113460);
   pc_target_reg_26_18_inst : DFFR_X1 port map( D => n5656, CK => Clk, RN => 
                           n3877, Q => pc_target_26_18_port, QN => net113459);
   pc_target_reg_26_20_inst : DFFR_X1 port map( D => n5655, CK => Clk, RN => 
                           n3877, Q => pc_target_26_20_port, QN => net113458);
   pc_target_reg_26_22_inst : DFFR_X1 port map( D => n5654, CK => Clk, RN => 
                           n3877, Q => pc_target_26_22_port, QN => net113457);
   pc_target_reg_26_24_inst : DFFR_X1 port map( D => n5653, CK => Clk, RN => 
                           n3877, Q => pc_target_26_24_port, QN => net113456);
   pc_target_reg_26_26_inst : DFFR_X1 port map( D => n5652, CK => Clk, RN => 
                           n3877, Q => pc_target_26_26_port, QN => net113455);
   pc_target_reg_26_28_inst : DFFR_X1 port map( D => n5651, CK => Clk, RN => 
                           n3877, Q => pc_target_26_28_port, QN => net113454);
   pc_target_reg_26_30_inst : DFFR_X1 port map( D => n5650, CK => Clk, RN => 
                           n3866, Q => pc_target_26_30_port, QN => net113453);
   pc_target_reg_27_31_inst : DFFR_X1 port map( D => n5649, CK => Clk, RN => 
                           n3888, Q => pc_target_27_31_port, QN => net113452);
   pc_target_reg_27_29_inst : DFFR_X1 port map( D => n5648, CK => Clk, RN => 
                           n3865, Q => pc_target_27_29_port, QN => net113451);
   pc_target_reg_27_27_inst : DFFR_X1 port map( D => n5647, CK => Clk, RN => 
                           n3865, Q => pc_target_27_27_port, QN => net113450);
   pc_target_reg_27_25_inst : DFFR_X1 port map( D => n5646, CK => Clk, RN => 
                           n3866, Q => pc_target_27_25_port, QN => net113449);
   pc_target_reg_27_23_inst : DFFR_X1 port map( D => n5645, CK => Clk, RN => 
                           n3866, Q => pc_target_27_23_port, QN => net113448);
   pc_target_reg_27_21_inst : DFFR_X1 port map( D => n5644, CK => Clk, RN => 
                           n3866, Q => pc_target_27_21_port, QN => net113447);
   pc_target_reg_27_19_inst : DFFR_X1 port map( D => n5643, CK => Clk, RN => 
                           n3866, Q => pc_target_27_19_port, QN => net113446);
   pc_target_reg_27_17_inst : DFFR_X1 port map( D => n5642, CK => Clk, RN => 
                           n3866, Q => pc_target_27_17_port, QN => net113445);
   pc_target_reg_27_15_inst : DFFR_X1 port map( D => n5641, CK => Clk, RN => 
                           n3866, Q => pc_target_27_15_port, QN => net113444);
   pc_target_reg_27_13_inst : DFFR_X1 port map( D => n5640, CK => Clk, RN => 
                           n3866, Q => pc_target_27_13_port, QN => net113443);
   pc_target_reg_27_11_inst : DFFR_X1 port map( D => n5639, CK => Clk, RN => 
                           n3866, Q => pc_target_27_11_port, QN => net113442);
   pc_target_reg_27_9_inst : DFFR_X1 port map( D => n5638, CK => Clk, RN => 
                           n3866, Q => pc_target_27_9_port, QN => net113441);
   pc_target_reg_27_7_inst : DFFR_X1 port map( D => n5637, CK => Clk, RN => 
                           n3866, Q => pc_target_27_7_port, QN => net113440);
   pc_target_reg_27_5_inst : DFFR_X1 port map( D => n5636, CK => Clk, RN => 
                           n3866, Q => pc_target_27_5_port, QN => net113439);
   pc_target_reg_27_3_inst : DFFR_X1 port map( D => n5635, CK => Clk, RN => 
                           n3866, Q => pc_target_27_3_port, QN => net113438);
   pc_target_reg_27_1_inst : DFFR_X1 port map( D => n5634, CK => Clk, RN => 
                           n3866, Q => pc_target_27_1_port, QN => net113437);
   pc_target_reg_27_0_inst : DFFR_X1 port map( D => n5633, CK => Clk, RN => 
                           n3867, Q => pc_target_27_0_port, QN => net113436);
   pc_target_reg_27_2_inst : DFFR_X1 port map( D => n5632, CK => Clk, RN => 
                           n3866, Q => pc_target_27_2_port, QN => net113435);
   pc_target_reg_27_4_inst : DFFR_X1 port map( D => n5631, CK => Clk, RN => 
                           n3867, Q => pc_target_27_4_port, QN => net113434);
   pc_target_reg_27_6_inst : DFFR_X1 port map( D => n5630, CK => Clk, RN => 
                           n3867, Q => pc_target_27_6_port, QN => net113433);
   pc_target_reg_27_8_inst : DFFR_X1 port map( D => n5629, CK => Clk, RN => 
                           n3867, Q => pc_target_27_8_port, QN => net113432);
   pc_target_reg_27_10_inst : DFFR_X1 port map( D => n5628, CK => Clk, RN => 
                           n3867, Q => pc_target_27_10_port, QN => net113431);
   pc_target_reg_27_12_inst : DFFR_X1 port map( D => n5627, CK => Clk, RN => 
                           n3867, Q => pc_target_27_12_port, QN => net113430);
   pc_target_reg_27_14_inst : DFFR_X1 port map( D => n5626, CK => Clk, RN => 
                           n3867, Q => pc_target_27_14_port, QN => net113429);
   pc_target_reg_27_16_inst : DFFR_X1 port map( D => n5625, CK => Clk, RN => 
                           n3867, Q => pc_target_27_16_port, QN => net113428);
   pc_target_reg_27_18_inst : DFFR_X1 port map( D => n5624, CK => Clk, RN => 
                           n3867, Q => pc_target_27_18_port, QN => net113427);
   pc_target_reg_27_20_inst : DFFR_X1 port map( D => n5623, CK => Clk, RN => 
                           n3867, Q => pc_target_27_20_port, QN => net113426);
   pc_target_reg_27_22_inst : DFFR_X1 port map( D => n5622, CK => Clk, RN => 
                           n3867, Q => pc_target_27_22_port, QN => net113425);
   pc_target_reg_27_24_inst : DFFR_X1 port map( D => n5621, CK => Clk, RN => 
                           n3867, Q => pc_target_27_24_port, QN => net113424);
   pc_target_reg_27_26_inst : DFFR_X1 port map( D => n5620, CK => Clk, RN => 
                           n3867, Q => pc_target_27_26_port, QN => net113423);
   pc_target_reg_27_28_inst : DFFR_X1 port map( D => n5619, CK => Clk, RN => 
                           n3867, Q => pc_target_27_28_port, QN => net113422);
   pc_target_reg_27_30_inst : DFFR_X1 port map( D => n5618, CK => Clk, RN => 
                           n3868, Q => pc_target_27_30_port, QN => net113421);
   pc_target_reg_28_31_inst : DFFR_X1 port map( D => n5617, CK => Clk, RN => 
                           n3865, Q => net113420, QN => n175);
   pc_target_reg_28_29_inst : DFFR_X1 port map( D => n5616, CK => Clk, RN => 
                           n3868, Q => net113419, QN => n174);
   pc_target_reg_28_27_inst : DFFR_X1 port map( D => n5615, CK => Clk, RN => 
                           n3868, Q => net113418, QN => n173);
   pc_target_reg_28_25_inst : DFFR_X1 port map( D => n5614, CK => Clk, RN => 
                           n3868, Q => net113417, QN => n172);
   pc_target_reg_28_23_inst : DFFR_X1 port map( D => n5613, CK => Clk, RN => 
                           n3868, Q => net113416, QN => n171);
   pc_target_reg_28_21_inst : DFFR_X1 port map( D => n5612, CK => Clk, RN => 
                           n3868, Q => net113415, QN => n170);
   pc_target_reg_28_19_inst : DFFR_X1 port map( D => n5611, CK => Clk, RN => 
                           n3868, Q => net113414, QN => n169);
   pc_target_reg_28_17_inst : DFFR_X1 port map( D => n5610, CK => Clk, RN => 
                           n3868, Q => net113413, QN => n168);
   pc_target_reg_28_15_inst : DFFR_X1 port map( D => n5609, CK => Clk, RN => 
                           n3868, Q => net113412, QN => n167);
   pc_target_reg_28_13_inst : DFFR_X1 port map( D => n5608, CK => Clk, RN => 
                           n3868, Q => net113411, QN => n166);
   pc_target_reg_28_11_inst : DFFR_X1 port map( D => n5607, CK => Clk, RN => 
                           n3868, Q => net113410, QN => n165);
   pc_target_reg_28_9_inst : DFFR_X1 port map( D => n5606, CK => Clk, RN => 
                           n3868, Q => net113409, QN => n164);
   pc_target_reg_28_7_inst : DFFR_X1 port map( D => n5605, CK => Clk, RN => 
                           n3868, Q => net113408, QN => n163);
   pc_target_reg_28_5_inst : DFFR_X1 port map( D => n5604, CK => Clk, RN => 
                           n3868, Q => n_1102, QN => n162);
   pc_target_reg_28_3_inst : DFFR_X1 port map( D => n5603, CK => Clk, RN => 
                           n3868, Q => net113406, QN => n161);
   pc_target_reg_28_1_inst : DFFR_X1 port map( D => n5602, CK => Clk, RN => 
                           n3869, Q => n_1103, QN => n160);
   pc_target_reg_28_0_inst : DFFR_X1 port map( D => n5601, CK => Clk, RN => 
                           n3869, Q => n_1104, QN => n159);
   pc_target_reg_28_2_inst : DFFR_X1 port map( D => n5600, CK => Clk, RN => 
                           n3869, Q => net113403, QN => n158);
   pc_target_reg_28_4_inst : DFFR_X1 port map( D => n5599, CK => Clk, RN => 
                           n3869, Q => n_1105, QN => n157);
   pc_target_reg_28_6_inst : DFFR_X1 port map( D => n5598, CK => Clk, RN => 
                           n3869, Q => n_1106, QN => n156);
   pc_target_reg_28_8_inst : DFFR_X1 port map( D => n5597, CK => Clk, RN => 
                           n3869, Q => net113400, QN => n155);
   pc_target_reg_28_10_inst : DFFR_X1 port map( D => n5596, CK => Clk, RN => 
                           n3869, Q => net113399, QN => n154);
   pc_target_reg_28_12_inst : DFFR_X1 port map( D => n5595, CK => Clk, RN => 
                           n3869, Q => net113398, QN => n153);
   pc_target_reg_28_14_inst : DFFR_X1 port map( D => n5594, CK => Clk, RN => 
                           n3869, Q => net113397, QN => n152);
   pc_target_reg_28_16_inst : DFFR_X1 port map( D => n5593, CK => Clk, RN => 
                           n3869, Q => net113396, QN => n151);
   pc_target_reg_28_18_inst : DFFR_X1 port map( D => n5592, CK => Clk, RN => 
                           n3869, Q => net113395, QN => n150);
   pc_target_reg_28_20_inst : DFFR_X1 port map( D => n5591, CK => Clk, RN => 
                           n3869, Q => net113394, QN => n149);
   pc_target_reg_28_22_inst : DFFR_X1 port map( D => n5590, CK => Clk, RN => 
                           n3869, Q => net113393, QN => n148);
   pc_target_reg_28_24_inst : DFFR_X1 port map( D => n5589, CK => Clk, RN => 
                           n3869, Q => net113392, QN => n147);
   pc_target_reg_28_26_inst : DFFR_X1 port map( D => n5588, CK => Clk, RN => 
                           n3869, Q => net113391, QN => n146);
   pc_target_reg_28_28_inst : DFFR_X1 port map( D => n5587, CK => Clk, RN => 
                           n3870, Q => net113390, QN => n145);
   pc_target_reg_29_31_inst : DFFR_X1 port map( D => n5585, CK => Clk, RN => 
                           n3865, Q => net113389, QN => n140);
   pc_target_reg_29_29_inst : DFFR_X1 port map( D => n5584, CK => Clk, RN => 
                           n3870, Q => net113388, QN => n138);
   pc_target_reg_29_27_inst : DFFR_X1 port map( D => n5583, CK => Clk, RN => 
                           n3870, Q => net113387, QN => n136);
   pc_target_reg_29_25_inst : DFFR_X1 port map( D => n5582, CK => Clk, RN => 
                           n3870, Q => net113386, QN => n134);
   pc_target_reg_29_23_inst : DFFR_X1 port map( D => n5581, CK => Clk, RN => 
                           n3870, Q => net113385, QN => n132);
   pc_target_reg_29_21_inst : DFFR_X1 port map( D => n5580, CK => Clk, RN => 
                           n3870, Q => net113384, QN => n130);
   pc_target_reg_29_19_inst : DFFR_X1 port map( D => n5579, CK => Clk, RN => 
                           n3870, Q => net113383, QN => n128);
   pc_target_reg_29_17_inst : DFFR_X1 port map( D => n5578, CK => Clk, RN => 
                           n3870, Q => net113382, QN => n126_port);
   pc_target_reg_29_15_inst : DFFR_X1 port map( D => n5577, CK => Clk, RN => 
                           n3870, Q => net113381, QN => n124_port);
   pc_target_reg_29_13_inst : DFFR_X1 port map( D => n5576, CK => Clk, RN => 
                           n3870, Q => net113380, QN => n122_port);
   pc_target_reg_29_11_inst : DFFR_X1 port map( D => n5575, CK => Clk, RN => 
                           n3870, Q => net113379, QN => n120_port);
   pc_target_reg_29_9_inst : DFFR_X1 port map( D => n5574, CK => Clk, RN => 
                           n3870, Q => net113378, QN => n118_port);
   pc_target_reg_29_7_inst : DFFR_X1 port map( D => n5573, CK => Clk, RN => 
                           n3870, Q => net113377, QN => n116_port);
   pc_target_reg_29_5_inst : DFFR_X1 port map( D => n5572, CK => Clk, RN => 
                           n3870, Q => n_1107, QN => n114_port);
   pc_target_reg_29_3_inst : DFFR_X1 port map( D => n5571, CK => Clk, RN => 
                           n3870, Q => net113375, QN => n112_port);
   pc_target_reg_29_1_inst : DFFR_X1 port map( D => n5570, CK => Clk, RN => 
                           n3871, Q => n_1108, QN => n110_port);
   pc_target_reg_29_0_inst : DFFR_X1 port map( D => n5569, CK => Clk, RN => 
                           n3871, Q => n_1109, QN => n108_port);
   pc_target_reg_29_2_inst : DFFR_X1 port map( D => n5568, CK => Clk, RN => 
                           n3871, Q => net113372, QN => n106_port);
   pc_target_reg_29_4_inst : DFFR_X1 port map( D => n5567, CK => Clk, RN => 
                           n3871, Q => n_1110, QN => n104_port);
   pc_target_reg_29_6_inst : DFFR_X1 port map( D => n5566, CK => Clk, RN => 
                           n3871, Q => n_1111, QN => n102_port);
   pc_target_reg_29_8_inst : DFFR_X1 port map( D => n5565, CK => Clk, RN => 
                           n3871, Q => net113369, QN => n100_port);
   pc_target_reg_29_10_inst : DFFR_X1 port map( D => n5564, CK => Clk, RN => 
                           n3871, Q => net113368, QN => n98_port);
   pc_target_reg_29_12_inst : DFFR_X1 port map( D => n5563, CK => Clk, RN => 
                           n3871, Q => net113367, QN => n96_port);
   pc_target_reg_29_14_inst : DFFR_X1 port map( D => n5562, CK => Clk, RN => 
                           n3871, Q => net113366, QN => n94);
   pc_target_reg_29_16_inst : DFFR_X1 port map( D => n5561, CK => Clk, RN => 
                           n3871, Q => net113365, QN => n92);
   pc_target_reg_29_18_inst : DFFR_X1 port map( D => n5560, CK => Clk, RN => 
                           n3871, Q => net113364, QN => n90);
   pc_target_reg_29_20_inst : DFFR_X1 port map( D => n5559, CK => Clk, RN => 
                           n3859, Q => net113363, QN => n88);
   pc_target_reg_29_22_inst : DFFR_X1 port map( D => n5558, CK => Clk, RN => 
                           n3855, Q => net113362, QN => n86);
   pc_target_reg_29_24_inst : DFFR_X1 port map( D => n5557, CK => Clk, RN => 
                           n3855, Q => net113361, QN => n84);
   pc_target_reg_29_26_inst : DFFR_X1 port map( D => n5556, CK => Clk, RN => 
                           n3855, Q => net113360, QN => n82);
   pc_target_reg_29_28_inst : DFFR_X1 port map( D => n5555, CK => Clk, RN => 
                           n3855, Q => net113359, QN => n80);
   pc_target_reg_30_31_inst : DFFR_X1 port map( D => n5553, CK => Clk, RN => 
                           n3867, Q => pc_target_30_31_port, QN => net113358);
   pc_target_reg_30_29_inst : DFFR_X1 port map( D => n5552, CK => Clk, RN => 
                           n3871, Q => pc_target_30_29_port, QN => net113357);
   pc_target_reg_30_27_inst : DFFR_X1 port map( D => n5551, CK => Clk, RN => 
                           n3871, Q => pc_target_30_27_port, QN => net113356);
   pc_target_reg_30_25_inst : DFFR_X1 port map( D => n5550, CK => Clk, RN => 
                           n3855, Q => pc_target_30_25_port, QN => net113355);
   pc_target_reg_30_23_inst : DFFR_X1 port map( D => n5549, CK => Clk, RN => 
                           n3856, Q => pc_target_30_23_port, QN => net113354);
   pc_target_reg_30_21_inst : DFFR_X1 port map( D => n5548, CK => Clk, RN => 
                           n3856, Q => pc_target_30_21_port, QN => net113353);
   pc_target_reg_30_19_inst : DFFR_X1 port map( D => n5547, CK => Clk, RN => 
                           n3856, Q => pc_target_30_19_port, QN => net113352);
   pc_target_reg_30_17_inst : DFFR_X1 port map( D => n5546, CK => Clk, RN => 
                           n3856, Q => pc_target_30_17_port, QN => net113351);
   pc_target_reg_30_15_inst : DFFR_X1 port map( D => n5545, CK => Clk, RN => 
                           n3856, Q => pc_target_30_15_port, QN => net113350);
   pc_target_reg_30_13_inst : DFFR_X1 port map( D => n5544, CK => Clk, RN => 
                           n3856, Q => pc_target_30_13_port, QN => net113349);
   pc_target_reg_30_11_inst : DFFR_X1 port map( D => n5543, CK => Clk, RN => 
                           n3856, Q => pc_target_30_11_port, QN => net113348);
   pc_target_reg_30_9_inst : DFFR_X1 port map( D => n5542, CK => Clk, RN => 
                           n3856, Q => pc_target_30_9_port, QN => net113347);
   pc_target_reg_30_7_inst : DFFR_X1 port map( D => n5541, CK => Clk, RN => 
                           n3856, Q => pc_target_30_7_port, QN => net113346);
   pc_target_reg_30_5_inst : DFFR_X1 port map( D => n5540, CK => Clk, RN => 
                           n3856, Q => pc_target_30_5_port, QN => net113345);
   pc_target_reg_30_3_inst : DFFR_X1 port map( D => n5539, CK => Clk, RN => 
                           n3856, Q => pc_target_30_3_port, QN => net113344);
   pc_target_reg_30_1_inst : DFFR_X1 port map( D => n5538, CK => Clk, RN => 
                           n3856, Q => pc_target_30_1_port, QN => net113343);
   pc_target_reg_30_0_inst : DFFR_X1 port map( D => n5537, CK => Clk, RN => 
                           n3857, Q => pc_target_30_0_port, QN => net113342);
   pc_target_reg_30_2_inst : DFFR_X1 port map( D => n5536, CK => Clk, RN => 
                           n3856, Q => pc_target_30_2_port, QN => net113341);
   pc_target_reg_30_4_inst : DFFR_X1 port map( D => n5535, CK => Clk, RN => 
                           n3856, Q => pc_target_30_4_port, QN => net113340);
   pc_target_reg_30_6_inst : DFFR_X1 port map( D => n5534, CK => Clk, RN => 
                           n3856, Q => pc_target_30_6_port, QN => net113339);
   pc_target_reg_30_8_inst : DFFR_X1 port map( D => n5533, CK => Clk, RN => 
                           n3857, Q => pc_target_30_8_port, QN => net113338);
   pc_target_reg_30_10_inst : DFFR_X1 port map( D => n5532, CK => Clk, RN => 
                           n3857, Q => pc_target_30_10_port, QN => net113337);
   pc_target_reg_30_12_inst : DFFR_X1 port map( D => n5531, CK => Clk, RN => 
                           n3857, Q => pc_target_30_12_port, QN => net113336);
   pc_target_reg_30_14_inst : DFFR_X1 port map( D => n5530, CK => Clk, RN => 
                           n3857, Q => pc_target_30_14_port, QN => net113335);
   pc_target_reg_30_16_inst : DFFR_X1 port map( D => n5529, CK => Clk, RN => 
                           n3857, Q => pc_target_30_16_port, QN => net113334);
   pc_target_reg_30_18_inst : DFFR_X1 port map( D => n5528, CK => Clk, RN => 
                           n3857, Q => pc_target_30_18_port, QN => net113333);
   pc_target_reg_30_20_inst : DFFR_X1 port map( D => n5527, CK => Clk, RN => 
                           n3857, Q => pc_target_30_20_port, QN => net113332);
   pc_target_reg_30_22_inst : DFFR_X1 port map( D => n5526, CK => Clk, RN => 
                           n3857, Q => pc_target_30_22_port, QN => net113331);
   pc_target_reg_30_24_inst : DFFR_X1 port map( D => n5525, CK => Clk, RN => 
                           n3857, Q => pc_target_30_24_port, QN => net113330);
   pc_target_reg_30_26_inst : DFFR_X1 port map( D => n5524, CK => Clk, RN => 
                           n3857, Q => pc_target_30_26_port, QN => net113329);
   pc_target_reg_30_28_inst : DFFR_X1 port map( D => n5523, CK => Clk, RN => 
                           n3857, Q => pc_target_30_28_port, QN => net113328);
   pc_target_reg_30_30_inst : DFFR_X1 port map( D => n5522, CK => Clk, RN => 
                           n3857, Q => pc_target_30_30_port, QN => net113327);
   pc_target_reg_31_31_inst : DFFR_X1 port map( D => n5521, CK => Clk, RN => 
                           n3863, Q => pc_target_31_31_port, QN => net113326);
   OUT_PC_target_reg_31_inst : DLH_X1 port map( G => Enable, D => N96, Q => 
                           OUT_PC_target(31));
   pc_target_reg_31_29_inst : DFFR_X1 port map( D => n5520, CK => Clk, RN => 
                           n3857, Q => pc_target_31_29_port, QN => net113325);
   OUT_PC_target_reg_29_inst : DLH_X1 port map( G => Enable, D => N98, Q => 
                           OUT_PC_target(29));
   pc_target_reg_31_27_inst : DFFR_X1 port map( D => n5519, CK => Clk, RN => 
                           n3857, Q => pc_target_31_27_port, QN => net113324);
   OUT_PC_target_reg_27_inst : DLH_X1 port map( G => Enable, D => N100, Q => 
                           OUT_PC_target(27));
   pc_target_reg_31_25_inst : DFFR_X1 port map( D => n5518, CK => Clk, RN => 
                           n3858, Q => pc_target_31_25_port, QN => net113323);
   OUT_PC_target_reg_25_inst : DLH_X1 port map( G => Enable, D => N102, Q => 
                           OUT_PC_target(25));
   pc_target_reg_31_23_inst : DFFR_X1 port map( D => n5517, CK => Clk, RN => 
                           n3858, Q => pc_target_31_23_port, QN => net113322);
   OUT_PC_target_reg_23_inst : DLH_X1 port map( G => Enable, D => N104, Q => 
                           OUT_PC_target(23));
   pc_target_reg_31_21_inst : DFFR_X1 port map( D => n5516, CK => Clk, RN => 
                           n3858, Q => pc_target_31_21_port, QN => net113321);
   OUT_PC_target_reg_21_inst : DLH_X1 port map( G => Enable, D => N106, Q => 
                           OUT_PC_target(21));
   pc_target_reg_31_19_inst : DFFR_X1 port map( D => n5515, CK => Clk, RN => 
                           n3858, Q => pc_target_31_19_port, QN => net113320);
   OUT_PC_target_reg_19_inst : DLH_X1 port map( G => Enable, D => N108, Q => 
                           OUT_PC_target(19));
   pc_target_reg_31_17_inst : DFFR_X1 port map( D => n5514, CK => Clk, RN => 
                           n3858, Q => pc_target_31_17_port, QN => net113319);
   OUT_PC_target_reg_17_inst : DLH_X1 port map( G => Enable, D => N110, Q => 
                           OUT_PC_target(17));
   pc_target_reg_31_15_inst : DFFR_X1 port map( D => n5513, CK => Clk, RN => 
                           n3858, Q => pc_target_31_15_port, QN => net113318);
   OUT_PC_target_reg_15_inst : DLH_X1 port map( G => Enable, D => N112, Q => 
                           OUT_PC_target(15));
   pc_target_reg_31_13_inst : DFFR_X1 port map( D => n5512, CK => Clk, RN => 
                           n3858, Q => pc_target_31_13_port, QN => net113317);
   OUT_PC_target_reg_13_inst : DLH_X1 port map( G => Enable, D => N114, Q => 
                           OUT_PC_target(13));
   pc_target_reg_31_11_inst : DFFR_X1 port map( D => n5511, CK => Clk, RN => 
                           n3858, Q => pc_target_31_11_port, QN => net113316);
   OUT_PC_target_reg_11_inst : DLH_X1 port map( G => Enable, D => N116, Q => 
                           OUT_PC_target(11));
   pc_target_reg_31_9_inst : DFFR_X1 port map( D => n5510, CK => Clk, RN => 
                           n3858, Q => pc_target_31_9_port, QN => net113315);
   OUT_PC_target_reg_9_inst : DLH_X1 port map( G => Enable, D => N118, Q => 
                           OUT_PC_target(9));
   pc_target_reg_31_7_inst : DFFR_X1 port map( D => n5509, CK => Clk, RN => 
                           n3858, Q => pc_target_31_7_port, QN => net113314);
   OUT_PC_target_reg_7_inst : DLH_X1 port map( G => Enable, D => N120, Q => 
                           OUT_PC_target(7));
   pc_target_reg_31_5_inst : DFFR_X1 port map( D => n5508, CK => Clk, RN => 
                           n3858, Q => pc_target_31_5_port, QN => net113313);
   OUT_PC_target_reg_5_inst : DLH_X1 port map( G => Enable, D => N122, Q => 
                           OUT_PC_target(5));
   pc_target_reg_31_3_inst : DFFR_X1 port map( D => n5507, CK => Clk, RN => 
                           n3860, Q => pc_target_31_3_port, QN => net113312);
   OUT_PC_target_reg_3_inst : DLH_X1 port map( G => Enable, D => N124, Q => 
                           OUT_PC_target(3));
   pc_target_reg_31_1_inst : DFFR_X1 port map( D => n5506, CK => Clk, RN => 
                           n3860, Q => pc_target_31_1_port, QN => net113311);
   OUT_PC_target_reg_1_inst : DLH_X1 port map( G => Enable, D => N126, Q => 
                           OUT_PC_target(1));
   pc_target_reg_31_0_inst : DFFR_X1 port map( D => n5505, CK => Clk, RN => 
                           n3861, Q => pc_target_31_0_port, QN => net113310);
   OUT_PC_target_reg_0_inst : DLH_X1 port map( G => Enable, D => N127, Q => 
                           OUT_PC_target(0));
   pc_target_reg_31_2_inst : DFFR_X1 port map( D => n5504, CK => Clk, RN => 
                           n3860, Q => pc_target_31_2_port, QN => net113309);
   OUT_PC_target_reg_2_inst : DLH_X1 port map( G => Enable, D => N125, Q => 
                           OUT_PC_target(2));
   pc_target_reg_31_4_inst : DFFR_X1 port map( D => n5503, CK => Clk, RN => 
                           n3861, Q => pc_target_31_4_port, QN => net113308);
   OUT_PC_target_reg_4_inst : DLH_X1 port map( G => Enable, D => N123, Q => 
                           OUT_PC_target(4));
   pc_target_reg_31_6_inst : DFFR_X1 port map( D => n5502, CK => Clk, RN => 
                           n3861, Q => pc_target_31_6_port, QN => net113307);
   OUT_PC_target_reg_6_inst : DLH_X1 port map( G => Enable, D => N121, Q => 
                           OUT_PC_target(6));
   pc_target_reg_31_8_inst : DFFR_X1 port map( D => n5501, CK => Clk, RN => 
                           n3861, Q => pc_target_31_8_port, QN => net113306);
   OUT_PC_target_reg_8_inst : DLH_X1 port map( G => Enable, D => N119, Q => 
                           OUT_PC_target(8));
   pc_target_reg_31_10_inst : DFFR_X1 port map( D => n5500, CK => Clk, RN => 
                           n3861, Q => pc_target_31_10_port, QN => net113305);
   OUT_PC_target_reg_10_inst : DLH_X1 port map( G => Enable, D => N117, Q => 
                           OUT_PC_target(10));
   pc_target_reg_31_12_inst : DFFR_X1 port map( D => n5499, CK => Clk, RN => 
                           n3861, Q => pc_target_31_12_port, QN => net113304);
   OUT_PC_target_reg_12_inst : DLH_X1 port map( G => Enable, D => N115, Q => 
                           OUT_PC_target(12));
   pc_target_reg_31_14_inst : DFFR_X1 port map( D => n5498, CK => Clk, RN => 
                           n3861, Q => pc_target_31_14_port, QN => net113303);
   OUT_PC_target_reg_14_inst : DLH_X1 port map( G => Enable, D => N113, Q => 
                           OUT_PC_target(14));
   pc_target_reg_31_16_inst : DFFR_X1 port map( D => n5497, CK => Clk, RN => 
                           n3861, Q => pc_target_31_16_port, QN => net113302);
   OUT_PC_target_reg_16_inst : DLH_X1 port map( G => Enable, D => N111, Q => 
                           OUT_PC_target(16));
   pc_target_reg_31_18_inst : DFFR_X1 port map( D => n5496, CK => Clk, RN => 
                           n3861, Q => pc_target_31_18_port, QN => net113301);
   OUT_PC_target_reg_18_inst : DLH_X1 port map( G => Enable, D => N109, Q => 
                           OUT_PC_target(18));
   pc_target_reg_31_20_inst : DFFR_X1 port map( D => n5495, CK => Clk, RN => 
                           n3863, Q => pc_target_31_20_port, QN => net113300);
   OUT_PC_target_reg_20_inst : DLH_X1 port map( G => Enable, D => N107, Q => 
                           OUT_PC_target(20));
   pc_target_reg_31_22_inst : DFFR_X1 port map( D => n5494, CK => Clk, RN => 
                           n3863, Q => pc_target_31_22_port, QN => net113299);
   OUT_PC_target_reg_22_inst : DLH_X1 port map( G => Enable, D => N105, Q => 
                           OUT_PC_target(22));
   pc_target_reg_31_24_inst : DFFR_X1 port map( D => n5493, CK => Clk, RN => 
                           n3863, Q => pc_target_31_24_port, QN => net113298);
   OUT_PC_target_reg_24_inst : DLH_X1 port map( G => Enable, D => N103, Q => 
                           OUT_PC_target(24));
   pc_target_reg_31_26_inst : DFFR_X1 port map( D => n5492, CK => Clk, RN => 
                           n3863, Q => pc_target_31_26_port, QN => net113297);
   OUT_PC_target_reg_26_inst : DLH_X1 port map( G => Enable, D => N101, Q => 
                           OUT_PC_target(26));
   pc_target_reg_31_28_inst : DFFR_X1 port map( D => n5491, CK => Clk, RN => 
                           n3864, Q => pc_target_31_28_port, QN => net113296);
   OUT_PC_target_reg_28_inst : DLH_X1 port map( G => Enable, D => N99, Q => 
                           OUT_PC_target(28));
   pc_target_reg_31_30_inst : DFFR_X1 port map( D => n5490, CK => Clk, RN => 
                           n3864, Q => pc_target_31_30_port, QN => net113295);
   OUT_PC_target_reg_30_inst : DLH_X1 port map( G => Enable, D => N97, Q => 
                           OUT_PC_target(30));
   U3 : INV_X1 port map( A => n4, ZN => n5490);
   U5 : AOI22_X1 port map( A1 => n5, A2 => Set_target(30), B1 => n6, B2 => 
                           pc_target_31_30_port, ZN => n4);
   U6 : INV_X1 port map( A => n7, ZN => n5491);
   U7 : AOI22_X1 port map( A1 => n5, A2 => Set_target(28), B1 => n6, B2 => 
                           pc_target_31_28_port, ZN => n7);
   U8 : INV_X1 port map( A => n8, ZN => n5492);
   U9 : AOI22_X1 port map( A1 => n5, A2 => Set_target(26), B1 => n6, B2 => 
                           pc_target_31_26_port, ZN => n8);
   U10 : INV_X1 port map( A => n9, ZN => n5493);
   U11 : AOI22_X1 port map( A1 => n5, A2 => Set_target(24), B1 => n6, B2 => 
                           pc_target_31_24_port, ZN => n9);
   U12 : INV_X1 port map( A => n10, ZN => n5494);
   U13 : AOI22_X1 port map( A1 => n5, A2 => Set_target(22), B1 => n6, B2 => 
                           pc_target_31_22_port, ZN => n10);
   U14 : INV_X1 port map( A => n11, ZN => n5495);
   U15 : AOI22_X1 port map( A1 => n5, A2 => Set_target(20), B1 => n6, B2 => 
                           pc_target_31_20_port, ZN => n11);
   U16 : INV_X1 port map( A => n12, ZN => n5496);
   U17 : AOI22_X1 port map( A1 => n5, A2 => Set_target(18), B1 => n6, B2 => 
                           pc_target_31_18_port, ZN => n12);
   U18 : INV_X1 port map( A => n13, ZN => n5497);
   U19 : AOI22_X1 port map( A1 => n5, A2 => Set_target(16), B1 => n6, B2 => 
                           pc_target_31_16_port, ZN => n13);
   U20 : INV_X1 port map( A => n14, ZN => n5498);
   U21 : AOI22_X1 port map( A1 => n5, A2 => Set_target(14), B1 => n6, B2 => 
                           pc_target_31_14_port, ZN => n14);
   U22 : INV_X1 port map( A => n15, ZN => n5499);
   U23 : AOI22_X1 port map( A1 => n5, A2 => Set_target(12), B1 => n6, B2 => 
                           pc_target_31_12_port, ZN => n15);
   U24 : INV_X1 port map( A => n16, ZN => n5500);
   U25 : AOI22_X1 port map( A1 => n5, A2 => Set_target(10), B1 => n6, B2 => 
                           pc_target_31_10_port, ZN => n16);
   U26 : INV_X1 port map( A => n17, ZN => n5501);
   U27 : AOI22_X1 port map( A1 => n5, A2 => Set_target(8), B1 => n6, B2 => 
                           pc_target_31_8_port, ZN => n17);
   U28 : INV_X1 port map( A => n18, ZN => n5502);
   U29 : AOI22_X1 port map( A1 => n5, A2 => Set_target(6), B1 => n6, B2 => 
                           pc_target_31_6_port, ZN => n18);
   U30 : INV_X1 port map( A => n19, ZN => n5503);
   U31 : AOI22_X1 port map( A1 => n5, A2 => Set_target(4), B1 => n6, B2 => 
                           pc_target_31_4_port, ZN => n19);
   U32 : INV_X1 port map( A => n20, ZN => n5504);
   U33 : AOI22_X1 port map( A1 => n5, A2 => Set_target(2), B1 => n6, B2 => 
                           pc_target_31_2_port, ZN => n20);
   U34 : INV_X1 port map( A => n21, ZN => n5505);
   U35 : AOI22_X1 port map( A1 => n5, A2 => Set_target(0), B1 => n6, B2 => 
                           pc_target_31_0_port, ZN => n21);
   U36 : INV_X1 port map( A => n22, ZN => n5506);
   U37 : AOI22_X1 port map( A1 => n5, A2 => Set_target(1), B1 => n6, B2 => 
                           pc_target_31_1_port, ZN => n22);
   U38 : INV_X1 port map( A => n23, ZN => n5507);
   U39 : AOI22_X1 port map( A1 => n5, A2 => Set_target(3), B1 => n6, B2 => 
                           pc_target_31_3_port, ZN => n23);
   U40 : INV_X1 port map( A => n24, ZN => n5508);
   U41 : AOI22_X1 port map( A1 => n5, A2 => Set_target(5), B1 => n6, B2 => 
                           pc_target_31_5_port, ZN => n24);
   U42 : INV_X1 port map( A => n25, ZN => n5509);
   U43 : AOI22_X1 port map( A1 => n5, A2 => Set_target(7), B1 => n6, B2 => 
                           pc_target_31_7_port, ZN => n25);
   U44 : INV_X1 port map( A => n26, ZN => n5510);
   U45 : AOI22_X1 port map( A1 => n5, A2 => Set_target(9), B1 => n6, B2 => 
                           pc_target_31_9_port, ZN => n26);
   U46 : INV_X1 port map( A => n27, ZN => n5511);
   U47 : AOI22_X1 port map( A1 => n5, A2 => Set_target(11), B1 => n6, B2 => 
                           pc_target_31_11_port, ZN => n27);
   U48 : INV_X1 port map( A => n28, ZN => n5512);
   U49 : AOI22_X1 port map( A1 => n5, A2 => Set_target(13), B1 => n6, B2 => 
                           pc_target_31_13_port, ZN => n28);
   U50 : INV_X1 port map( A => n29, ZN => n5513);
   U51 : AOI22_X1 port map( A1 => n5, A2 => Set_target(15), B1 => n6, B2 => 
                           pc_target_31_15_port, ZN => n29);
   U52 : INV_X1 port map( A => n30, ZN => n5514);
   U53 : AOI22_X1 port map( A1 => n5, A2 => Set_target(17), B1 => n6, B2 => 
                           pc_target_31_17_port, ZN => n30);
   U54 : INV_X1 port map( A => n31, ZN => n5515);
   U55 : AOI22_X1 port map( A1 => n5, A2 => Set_target(19), B1 => n6, B2 => 
                           pc_target_31_19_port, ZN => n31);
   U56 : INV_X1 port map( A => n32, ZN => n5516);
   U57 : AOI22_X1 port map( A1 => n5, A2 => Set_target(21), B1 => n6, B2 => 
                           pc_target_31_21_port, ZN => n32);
   U58 : INV_X1 port map( A => n33, ZN => n5517);
   U59 : AOI22_X1 port map( A1 => n5, A2 => Set_target(23), B1 => n6, B2 => 
                           pc_target_31_23_port, ZN => n33);
   U60 : INV_X1 port map( A => n34, ZN => n5518);
   U61 : AOI22_X1 port map( A1 => n5, A2 => Set_target(25), B1 => n6, B2 => 
                           pc_target_31_25_port, ZN => n34);
   U62 : INV_X1 port map( A => n35, ZN => n5519);
   U63 : AOI22_X1 port map( A1 => n5, A2 => Set_target(27), B1 => n6, B2 => 
                           pc_target_31_27_port, ZN => n35);
   U64 : INV_X1 port map( A => n36, ZN => n5520);
   U65 : AOI22_X1 port map( A1 => n5, A2 => Set_target(29), B1 => n6, B2 => 
                           pc_target_31_29_port, ZN => n36);
   U66 : INV_X1 port map( A => n37, ZN => n5521);
   U67 : AOI22_X1 port map( A1 => n5, A2 => Set_target(31), B1 => n6, B2 => 
                           pc_target_31_31_port, ZN => n37);
   U70 : INV_X1 port map( A => n40, ZN => n5522);
   U71 : AOI22_X1 port map( A1 => Set_target(30), A2 => n3798, B1 => n42, B2 =>
                           pc_target_30_30_port, ZN => n40);
   U72 : INV_X1 port map( A => n43, ZN => n5523);
   U73 : AOI22_X1 port map( A1 => Set_target(28), A2 => n3798, B1 => n42, B2 =>
                           pc_target_30_28_port, ZN => n43);
   U74 : INV_X1 port map( A => n44, ZN => n5524);
   U75 : AOI22_X1 port map( A1 => Set_target(26), A2 => n3798, B1 => n42, B2 =>
                           pc_target_30_26_port, ZN => n44);
   U76 : INV_X1 port map( A => n45, ZN => n5525);
   U77 : AOI22_X1 port map( A1 => Set_target(24), A2 => n3798, B1 => n42, B2 =>
                           pc_target_30_24_port, ZN => n45);
   U78 : INV_X1 port map( A => n46, ZN => n5526);
   U79 : AOI22_X1 port map( A1 => Set_target(22), A2 => n3798, B1 => n42, B2 =>
                           pc_target_30_22_port, ZN => n46);
   U80 : INV_X1 port map( A => n47, ZN => n5527);
   U81 : AOI22_X1 port map( A1 => Set_target(20), A2 => n3798, B1 => n42, B2 =>
                           pc_target_30_20_port, ZN => n47);
   U82 : INV_X1 port map( A => n48, ZN => n5528);
   U83 : AOI22_X1 port map( A1 => Set_target(18), A2 => n3798, B1 => n42, B2 =>
                           pc_target_30_18_port, ZN => n48);
   U84 : INV_X1 port map( A => n49, ZN => n5529);
   U85 : AOI22_X1 port map( A1 => Set_target(16), A2 => n3798, B1 => n42, B2 =>
                           pc_target_30_16_port, ZN => n49);
   U86 : INV_X1 port map( A => n50, ZN => n5530);
   U87 : AOI22_X1 port map( A1 => Set_target(14), A2 => n3798, B1 => n42, B2 =>
                           pc_target_30_14_port, ZN => n50);
   U88 : INV_X1 port map( A => n51, ZN => n5531);
   U89 : AOI22_X1 port map( A1 => Set_target(12), A2 => n3798, B1 => n42, B2 =>
                           pc_target_30_12_port, ZN => n51);
   U90 : INV_X1 port map( A => n52, ZN => n5532);
   U91 : AOI22_X1 port map( A1 => Set_target(10), A2 => n3798, B1 => n42, B2 =>
                           pc_target_30_10_port, ZN => n52);
   U92 : INV_X1 port map( A => n53, ZN => n5533);
   U93 : AOI22_X1 port map( A1 => Set_target(8), A2 => n3798, B1 => n42, B2 => 
                           pc_target_30_8_port, ZN => n53);
   U94 : INV_X1 port map( A => n54, ZN => n5534);
   U95 : AOI22_X1 port map( A1 => Set_target(6), A2 => n3798, B1 => n42, B2 => 
                           pc_target_30_6_port, ZN => n54);
   U96 : INV_X1 port map( A => n55, ZN => n5535);
   U97 : AOI22_X1 port map( A1 => Set_target(4), A2 => n3798, B1 => n42, B2 => 
                           pc_target_30_4_port, ZN => n55);
   U98 : INV_X1 port map( A => n56, ZN => n5536);
   U99 : AOI22_X1 port map( A1 => Set_target(2), A2 => n3798, B1 => n42, B2 => 
                           pc_target_30_2_port, ZN => n56);
   U100 : INV_X1 port map( A => n57, ZN => n5537);
   U101 : AOI22_X1 port map( A1 => Set_target(0), A2 => n3798, B1 => n42, B2 =>
                           pc_target_30_0_port, ZN => n57);
   U102 : INV_X1 port map( A => n58, ZN => n5538);
   U103 : AOI22_X1 port map( A1 => Set_target(1), A2 => n3798, B1 => n42, B2 =>
                           pc_target_30_1_port, ZN => n58);
   U104 : INV_X1 port map( A => n59, ZN => n5539);
   U105 : AOI22_X1 port map( A1 => Set_target(3), A2 => n3798, B1 => n42, B2 =>
                           pc_target_30_3_port, ZN => n59);
   U106 : INV_X1 port map( A => n60, ZN => n5540);
   U107 : AOI22_X1 port map( A1 => Set_target(5), A2 => n3798, B1 => n42, B2 =>
                           pc_target_30_5_port, ZN => n60);
   U108 : INV_X1 port map( A => n61, ZN => n5541);
   U109 : AOI22_X1 port map( A1 => Set_target(7), A2 => n3798, B1 => n42, B2 =>
                           pc_target_30_7_port, ZN => n61);
   U110 : INV_X1 port map( A => n62, ZN => n5542);
   U111 : AOI22_X1 port map( A1 => Set_target(9), A2 => n3798, B1 => n42, B2 =>
                           pc_target_30_9_port, ZN => n62);
   U112 : INV_X1 port map( A => n63, ZN => n5543);
   U113 : AOI22_X1 port map( A1 => Set_target(11), A2 => n3798, B1 => n42, B2 
                           => pc_target_30_11_port, ZN => n63);
   U114 : INV_X1 port map( A => n64, ZN => n5544);
   U115 : AOI22_X1 port map( A1 => Set_target(13), A2 => n3798, B1 => n42, B2 
                           => pc_target_30_13_port, ZN => n64);
   U116 : INV_X1 port map( A => n65, ZN => n5545);
   U117 : AOI22_X1 port map( A1 => Set_target(15), A2 => n3798, B1 => n42, B2 
                           => pc_target_30_15_port, ZN => n65);
   U118 : INV_X1 port map( A => n66, ZN => n5546);
   U119 : AOI22_X1 port map( A1 => Set_target(17), A2 => n3798, B1 => n42, B2 
                           => pc_target_30_17_port, ZN => n66);
   U120 : INV_X1 port map( A => n67, ZN => n5547);
   U121 : AOI22_X1 port map( A1 => Set_target(19), A2 => n3798, B1 => n42, B2 
                           => pc_target_30_19_port, ZN => n67);
   U122 : INV_X1 port map( A => n68, ZN => n5548);
   U123 : AOI22_X1 port map( A1 => Set_target(21), A2 => n3798, B1 => n42, B2 
                           => pc_target_30_21_port, ZN => n68);
   U124 : INV_X1 port map( A => n69, ZN => n5549);
   U125 : AOI22_X1 port map( A1 => Set_target(23), A2 => n3798, B1 => n42, B2 
                           => pc_target_30_23_port, ZN => n69);
   U126 : INV_X1 port map( A => n70, ZN => n5550);
   U127 : AOI22_X1 port map( A1 => Set_target(25), A2 => n3798, B1 => n42, B2 
                           => pc_target_30_25_port, ZN => n70);
   U128 : INV_X1 port map( A => n71, ZN => n5551);
   U129 : AOI22_X1 port map( A1 => Set_target(27), A2 => n3798, B1 => n42, B2 
                           => pc_target_30_27_port, ZN => n71);
   U130 : INV_X1 port map( A => n72, ZN => n5552);
   U131 : AOI22_X1 port map( A1 => Set_target(29), A2 => n3798, B1 => n42, B2 
                           => pc_target_30_29_port, ZN => n72);
   U132 : INV_X1 port map( A => n73, ZN => n5553);
   U133 : AOI22_X1 port map( A1 => Set_target(31), A2 => n3798, B1 => n42, B2 
                           => pc_target_30_31_port, ZN => n73);
   U136 : OAI22_X1 port map( A1 => n75, A2 => n76, B1 => n77, B2 => n78, ZN => 
                           n5554);
   U137 : OAI22_X1 port map( A1 => n79, A2 => n76, B1 => n77, B2 => n80, ZN => 
                           n5555);
   U138 : OAI22_X1 port map( A1 => n81, A2 => n76, B1 => n77, B2 => n82, ZN => 
                           n5556);
   U139 : OAI22_X1 port map( A1 => n83, A2 => n76, B1 => n77, B2 => n84, ZN => 
                           n5557);
   U140 : OAI22_X1 port map( A1 => n85, A2 => n76, B1 => n77, B2 => n86, ZN => 
                           n5558);
   U141 : OAI22_X1 port map( A1 => n87, A2 => n76, B1 => n77, B2 => n88, ZN => 
                           n5559);
   U142 : OAI22_X1 port map( A1 => n89, A2 => n76, B1 => n77, B2 => n90, ZN => 
                           n5560);
   U143 : OAI22_X1 port map( A1 => n91, A2 => n76, B1 => n77, B2 => n92, ZN => 
                           n5561);
   U144 : OAI22_X1 port map( A1 => n93, A2 => n76, B1 => n77, B2 => n94, ZN => 
                           n5562);
   U145 : OAI22_X1 port map( A1 => n95, A2 => n76, B1 => n77, B2 => n96_port, 
                           ZN => n5563);
   U146 : OAI22_X1 port map( A1 => n97_port, A2 => n76, B1 => n77, B2 => 
                           n98_port, ZN => n5564);
   U147 : OAI22_X1 port map( A1 => n99_port, A2 => n76, B1 => n77, B2 => 
                           n100_port, ZN => n5565);
   U148 : OAI22_X1 port map( A1 => n101_port, A2 => n76, B1 => n77, B2 => 
                           n102_port, ZN => n5566);
   U149 : OAI22_X1 port map( A1 => n103_port, A2 => n76, B1 => n77, B2 => 
                           n104_port, ZN => n5567);
   U150 : OAI22_X1 port map( A1 => n105_port, A2 => n76, B1 => n77, B2 => 
                           n106_port, ZN => n5568);
   U151 : OAI22_X1 port map( A1 => n107_port, A2 => n76, B1 => n77, B2 => 
                           n108_port, ZN => n5569);
   U152 : OAI22_X1 port map( A1 => n109_port, A2 => n76, B1 => n77, B2 => 
                           n110_port, ZN => n5570);
   U153 : OAI22_X1 port map( A1 => n111_port, A2 => n76, B1 => n77, B2 => 
                           n112_port, ZN => n5571);
   U154 : OAI22_X1 port map( A1 => n113_port, A2 => n76, B1 => n77, B2 => 
                           n114_port, ZN => n5572);
   U155 : OAI22_X1 port map( A1 => n115_port, A2 => n76, B1 => n77, B2 => 
                           n116_port, ZN => n5573);
   U156 : OAI22_X1 port map( A1 => n117_port, A2 => n76, B1 => n77, B2 => 
                           n118_port, ZN => n5574);
   U157 : OAI22_X1 port map( A1 => n119_port, A2 => n76, B1 => n77, B2 => 
                           n120_port, ZN => n5575);
   U158 : OAI22_X1 port map( A1 => n121_port, A2 => n76, B1 => n77, B2 => 
                           n122_port, ZN => n5576);
   U159 : OAI22_X1 port map( A1 => n123_port, A2 => n76, B1 => n77, B2 => 
                           n124_port, ZN => n5577);
   U160 : OAI22_X1 port map( A1 => n125_port, A2 => n76, B1 => n77, B2 => 
                           n126_port, ZN => n5578);
   U161 : OAI22_X1 port map( A1 => n127_port, A2 => n76, B1 => n77, B2 => n128,
                           ZN => n5579);
   U162 : OAI22_X1 port map( A1 => n129, A2 => n76, B1 => n77, B2 => n130, ZN 
                           => n5580);
   U163 : OAI22_X1 port map( A1 => n131, A2 => n76, B1 => n77, B2 => n132, ZN 
                           => n5581);
   U164 : OAI22_X1 port map( A1 => n133, A2 => n76, B1 => n77, B2 => n134, ZN 
                           => n5582);
   U165 : OAI22_X1 port map( A1 => n135, A2 => n76, B1 => n77, B2 => n136, ZN 
                           => n5583);
   U166 : OAI22_X1 port map( A1 => n137, A2 => n76, B1 => n77, B2 => n138, ZN 
                           => n5584);
   U167 : OAI22_X1 port map( A1 => n139, A2 => n76, B1 => n77, B2 => n140, ZN 
                           => n5585);
   U170 : OAI22_X1 port map( A1 => n75, A2 => n142, B1 => n143, B2 => n144, ZN 
                           => n5586);
   U171 : OAI22_X1 port map( A1 => n79, A2 => n142, B1 => n143, B2 => n145, ZN 
                           => n5587);
   U172 : OAI22_X1 port map( A1 => n81, A2 => n142, B1 => n143, B2 => n146, ZN 
                           => n5588);
   U173 : OAI22_X1 port map( A1 => n83, A2 => n142, B1 => n143, B2 => n147, ZN 
                           => n5589);
   U174 : OAI22_X1 port map( A1 => n85, A2 => n142, B1 => n143, B2 => n148, ZN 
                           => n5590);
   U175 : OAI22_X1 port map( A1 => n87, A2 => n142, B1 => n143, B2 => n149, ZN 
                           => n5591);
   U176 : OAI22_X1 port map( A1 => n89, A2 => n142, B1 => n143, B2 => n150, ZN 
                           => n5592);
   U177 : OAI22_X1 port map( A1 => n91, A2 => n142, B1 => n143, B2 => n151, ZN 
                           => n5593);
   U178 : OAI22_X1 port map( A1 => n93, A2 => n142, B1 => n143, B2 => n152, ZN 
                           => n5594);
   U179 : OAI22_X1 port map( A1 => n95, A2 => n142, B1 => n143, B2 => n153, ZN 
                           => n5595);
   U180 : OAI22_X1 port map( A1 => n97_port, A2 => n142, B1 => n143, B2 => n154
                           , ZN => n5596);
   U181 : OAI22_X1 port map( A1 => n99_port, A2 => n142, B1 => n143, B2 => n155
                           , ZN => n5597);
   U182 : OAI22_X1 port map( A1 => n101_port, A2 => n142, B1 => n143, B2 => 
                           n156, ZN => n5598);
   U183 : OAI22_X1 port map( A1 => n103_port, A2 => n142, B1 => n143, B2 => 
                           n157, ZN => n5599);
   U184 : OAI22_X1 port map( A1 => n105_port, A2 => n142, B1 => n143, B2 => 
                           n158, ZN => n5600);
   U185 : OAI22_X1 port map( A1 => n107_port, A2 => n142, B1 => n143, B2 => 
                           n159, ZN => n5601);
   U186 : OAI22_X1 port map( A1 => n109_port, A2 => n142, B1 => n143, B2 => 
                           n160, ZN => n5602);
   U187 : OAI22_X1 port map( A1 => n111_port, A2 => n142, B1 => n143, B2 => 
                           n161, ZN => n5603);
   U188 : OAI22_X1 port map( A1 => n113_port, A2 => n142, B1 => n143, B2 => 
                           n162, ZN => n5604);
   U189 : OAI22_X1 port map( A1 => n115_port, A2 => n142, B1 => n143, B2 => 
                           n163, ZN => n5605);
   U190 : OAI22_X1 port map( A1 => n117_port, A2 => n142, B1 => n143, B2 => 
                           n164, ZN => n5606);
   U191 : OAI22_X1 port map( A1 => n119_port, A2 => n142, B1 => n143, B2 => 
                           n165, ZN => n5607);
   U192 : OAI22_X1 port map( A1 => n121_port, A2 => n142, B1 => n143, B2 => 
                           n166, ZN => n5608);
   U193 : OAI22_X1 port map( A1 => n123_port, A2 => n142, B1 => n143, B2 => 
                           n167, ZN => n5609);
   U194 : OAI22_X1 port map( A1 => n125_port, A2 => n142, B1 => n143, B2 => 
                           n168, ZN => n5610);
   U195 : OAI22_X1 port map( A1 => n127_port, A2 => n142, B1 => n143, B2 => 
                           n169, ZN => n5611);
   U196 : OAI22_X1 port map( A1 => n129, A2 => n142, B1 => n143, B2 => n170, ZN
                           => n5612);
   U197 : OAI22_X1 port map( A1 => n131, A2 => n142, B1 => n143, B2 => n171, ZN
                           => n5613);
   U198 : OAI22_X1 port map( A1 => n133, A2 => n142, B1 => n143, B2 => n172, ZN
                           => n5614);
   U199 : OAI22_X1 port map( A1 => n135, A2 => n142, B1 => n143, B2 => n173, ZN
                           => n5615);
   U200 : OAI22_X1 port map( A1 => n137, A2 => n142, B1 => n143, B2 => n174, ZN
                           => n5616);
   U201 : OAI22_X1 port map( A1 => n139, A2 => n142, B1 => n143, B2 => n175, ZN
                           => n5617);
   U205 : INV_X1 port map( A => n179, ZN => n5618);
   U206 : AOI22_X1 port map( A1 => Set_target(30), A2 => n3797, B1 => n181, B2 
                           => pc_target_27_30_port, ZN => n179);
   U207 : INV_X1 port map( A => n182, ZN => n5619);
   U208 : AOI22_X1 port map( A1 => Set_target(28), A2 => n3797, B1 => n181, B2 
                           => pc_target_27_28_port, ZN => n182);
   U209 : INV_X1 port map( A => n183, ZN => n5620);
   U210 : AOI22_X1 port map( A1 => Set_target(26), A2 => n3797, B1 => n181, B2 
                           => pc_target_27_26_port, ZN => n183);
   U211 : INV_X1 port map( A => n184, ZN => n5621);
   U212 : AOI22_X1 port map( A1 => Set_target(24), A2 => n3797, B1 => n181, B2 
                           => pc_target_27_24_port, ZN => n184);
   U213 : INV_X1 port map( A => n185, ZN => n5622);
   U214 : AOI22_X1 port map( A1 => Set_target(22), A2 => n3797, B1 => n181, B2 
                           => pc_target_27_22_port, ZN => n185);
   U215 : INV_X1 port map( A => n186, ZN => n5623);
   U216 : AOI22_X1 port map( A1 => Set_target(20), A2 => n3797, B1 => n181, B2 
                           => pc_target_27_20_port, ZN => n186);
   U217 : INV_X1 port map( A => n187, ZN => n5624);
   U218 : AOI22_X1 port map( A1 => Set_target(18), A2 => n3797, B1 => n181, B2 
                           => pc_target_27_18_port, ZN => n187);
   U219 : INV_X1 port map( A => n188_port, ZN => n5625);
   U220 : AOI22_X1 port map( A1 => Set_target(16), A2 => n3797, B1 => n181, B2 
                           => pc_target_27_16_port, ZN => n188_port);
   U221 : INV_X1 port map( A => n189_port, ZN => n5626);
   U222 : AOI22_X1 port map( A1 => Set_target(14), A2 => n3797, B1 => n181, B2 
                           => pc_target_27_14_port, ZN => n189_port);
   U223 : INV_X1 port map( A => n190_port, ZN => n5627);
   U224 : AOI22_X1 port map( A1 => Set_target(12), A2 => n3797, B1 => n181, B2 
                           => pc_target_27_12_port, ZN => n190_port);
   U225 : INV_X1 port map( A => n191_port, ZN => n5628);
   U226 : AOI22_X1 port map( A1 => Set_target(10), A2 => n3797, B1 => n181, B2 
                           => pc_target_27_10_port, ZN => n191_port);
   U227 : INV_X1 port map( A => n192_port, ZN => n5629);
   U228 : AOI22_X1 port map( A1 => Set_target(8), A2 => n3797, B1 => n181, B2 
                           => pc_target_27_8_port, ZN => n192_port);
   U229 : INV_X1 port map( A => n193_port, ZN => n5630);
   U230 : AOI22_X1 port map( A1 => Set_target(6), A2 => n3797, B1 => n181, B2 
                           => pc_target_27_6_port, ZN => n193_port);
   U231 : INV_X1 port map( A => n194_port, ZN => n5631);
   U232 : AOI22_X1 port map( A1 => Set_target(4), A2 => n3797, B1 => n181, B2 
                           => pc_target_27_4_port, ZN => n194_port);
   U233 : INV_X1 port map( A => n195_port, ZN => n5632);
   U234 : AOI22_X1 port map( A1 => Set_target(2), A2 => n3797, B1 => n181, B2 
                           => pc_target_27_2_port, ZN => n195_port);
   U235 : INV_X1 port map( A => n196_port, ZN => n5633);
   U236 : AOI22_X1 port map( A1 => Set_target(0), A2 => n3797, B1 => n181, B2 
                           => pc_target_27_0_port, ZN => n196_port);
   U237 : INV_X1 port map( A => n197_port, ZN => n5634);
   U238 : AOI22_X1 port map( A1 => Set_target(1), A2 => n3797, B1 => n181, B2 
                           => pc_target_27_1_port, ZN => n197_port);
   U239 : INV_X1 port map( A => n198_port, ZN => n5635);
   U240 : AOI22_X1 port map( A1 => Set_target(3), A2 => n3797, B1 => n181, B2 
                           => pc_target_27_3_port, ZN => n198_port);
   U241 : INV_X1 port map( A => n199_port, ZN => n5636);
   U242 : AOI22_X1 port map( A1 => Set_target(5), A2 => n3797, B1 => n181, B2 
                           => pc_target_27_5_port, ZN => n199_port);
   U243 : INV_X1 port map( A => n200_port, ZN => n5637);
   U244 : AOI22_X1 port map( A1 => Set_target(7), A2 => n3797, B1 => n181, B2 
                           => pc_target_27_7_port, ZN => n200_port);
   U245 : INV_X1 port map( A => n201_port, ZN => n5638);
   U246 : AOI22_X1 port map( A1 => Set_target(9), A2 => n3797, B1 => n181, B2 
                           => pc_target_27_9_port, ZN => n201_port);
   U247 : INV_X1 port map( A => n202_port, ZN => n5639);
   U248 : AOI22_X1 port map( A1 => Set_target(11), A2 => n3797, B1 => n181, B2 
                           => pc_target_27_11_port, ZN => n202_port);
   U249 : INV_X1 port map( A => n203_port, ZN => n5640);
   U250 : AOI22_X1 port map( A1 => Set_target(13), A2 => n3797, B1 => n181, B2 
                           => pc_target_27_13_port, ZN => n203_port);
   U251 : INV_X1 port map( A => n204_port, ZN => n5641);
   U252 : AOI22_X1 port map( A1 => Set_target(15), A2 => n3797, B1 => n181, B2 
                           => pc_target_27_15_port, ZN => n204_port);
   U253 : INV_X1 port map( A => n205_port, ZN => n5642);
   U254 : AOI22_X1 port map( A1 => Set_target(17), A2 => n3797, B1 => n181, B2 
                           => pc_target_27_17_port, ZN => n205_port);
   U255 : INV_X1 port map( A => n206_port, ZN => n5643);
   U256 : AOI22_X1 port map( A1 => Set_target(19), A2 => n3797, B1 => n181, B2 
                           => pc_target_27_19_port, ZN => n206_port);
   U257 : INV_X1 port map( A => n207_port, ZN => n5644);
   U258 : AOI22_X1 port map( A1 => Set_target(21), A2 => n3797, B1 => n181, B2 
                           => pc_target_27_21_port, ZN => n207_port);
   U259 : INV_X1 port map( A => n208_port, ZN => n5645);
   U260 : AOI22_X1 port map( A1 => Set_target(23), A2 => n3797, B1 => n181, B2 
                           => pc_target_27_23_port, ZN => n208_port);
   U261 : INV_X1 port map( A => n209_port, ZN => n5646);
   U262 : AOI22_X1 port map( A1 => Set_target(25), A2 => n3797, B1 => n181, B2 
                           => pc_target_27_25_port, ZN => n209_port);
   U263 : INV_X1 port map( A => n210_port, ZN => n5647);
   U264 : AOI22_X1 port map( A1 => Set_target(27), A2 => n3797, B1 => n181, B2 
                           => pc_target_27_27_port, ZN => n210_port);
   U265 : INV_X1 port map( A => n211_port, ZN => n5648);
   U266 : AOI22_X1 port map( A1 => Set_target(29), A2 => n3797, B1 => n181, B2 
                           => pc_target_27_29_port, ZN => n211_port);
   U267 : INV_X1 port map( A => n212_port, ZN => n5649);
   U268 : AOI22_X1 port map( A1 => Set_target(31), A2 => n3797, B1 => n181, B2 
                           => pc_target_27_31_port, ZN => n212_port);
   U271 : INV_X1 port map( A => n214_port, ZN => n5650);
   U272 : AOI22_X1 port map( A1 => Set_target(30), A2 => n215_port, B1 => 
                           n216_port, B2 => pc_target_26_30_port, ZN => 
                           n214_port);
   U273 : INV_X1 port map( A => n217_port, ZN => n5651);
   U274 : AOI22_X1 port map( A1 => Set_target(28), A2 => n215_port, B1 => 
                           n216_port, B2 => pc_target_26_28_port, ZN => 
                           n217_port);
   U275 : INV_X1 port map( A => n218_port, ZN => n5652);
   U276 : AOI22_X1 port map( A1 => Set_target(26), A2 => n215_port, B1 => 
                           n216_port, B2 => pc_target_26_26_port, ZN => 
                           n218_port);
   U277 : INV_X1 port map( A => n219_port, ZN => n5653);
   U278 : AOI22_X1 port map( A1 => Set_target(24), A2 => n215_port, B1 => 
                           n216_port, B2 => pc_target_26_24_port, ZN => 
                           n219_port);
   U279 : INV_X1 port map( A => n220_port, ZN => n5654);
   U280 : AOI22_X1 port map( A1 => Set_target(22), A2 => n215_port, B1 => 
                           n216_port, B2 => pc_target_26_22_port, ZN => 
                           n220_port);
   U281 : INV_X1 port map( A => n221, ZN => n5655);
   U282 : AOI22_X1 port map( A1 => Set_target(20), A2 => n215_port, B1 => 
                           n216_port, B2 => pc_target_26_20_port, ZN => n221);
   U283 : INV_X1 port map( A => n222, ZN => n5656);
   U284 : AOI22_X1 port map( A1 => Set_target(18), A2 => n215_port, B1 => 
                           n216_port, B2 => pc_target_26_18_port, ZN => n222);
   U285 : INV_X1 port map( A => n223, ZN => n5657);
   U286 : AOI22_X1 port map( A1 => Set_target(16), A2 => n215_port, B1 => 
                           n216_port, B2 => pc_target_26_16_port, ZN => n223);
   U287 : INV_X1 port map( A => n224, ZN => n5658);
   U288 : AOI22_X1 port map( A1 => Set_target(14), A2 => n215_port, B1 => 
                           n216_port, B2 => pc_target_26_14_port, ZN => n224);
   U289 : INV_X1 port map( A => n225, ZN => n5659);
   U290 : AOI22_X1 port map( A1 => Set_target(12), A2 => n215_port, B1 => 
                           n216_port, B2 => pc_target_26_12_port, ZN => n225);
   U291 : INV_X1 port map( A => n226, ZN => n5660);
   U292 : AOI22_X1 port map( A1 => Set_target(10), A2 => n215_port, B1 => 
                           n216_port, B2 => pc_target_26_10_port, ZN => n226);
   U293 : INV_X1 port map( A => n227, ZN => n5661);
   U294 : AOI22_X1 port map( A1 => Set_target(8), A2 => n215_port, B1 => 
                           n216_port, B2 => pc_target_26_8_port, ZN => n227);
   U295 : INV_X1 port map( A => n228, ZN => n5662);
   U296 : AOI22_X1 port map( A1 => Set_target(6), A2 => n215_port, B1 => 
                           n216_port, B2 => pc_target_26_6_port, ZN => n228);
   U297 : INV_X1 port map( A => n229, ZN => n5663);
   U298 : AOI22_X1 port map( A1 => Set_target(4), A2 => n215_port, B1 => 
                           n216_port, B2 => pc_target_26_4_port, ZN => n229);
   U299 : INV_X1 port map( A => n230, ZN => n5664);
   U300 : AOI22_X1 port map( A1 => Set_target(2), A2 => n215_port, B1 => 
                           n216_port, B2 => pc_target_26_2_port, ZN => n230);
   U301 : INV_X1 port map( A => n231, ZN => n5665);
   U302 : AOI22_X1 port map( A1 => Set_target(0), A2 => n215_port, B1 => 
                           n216_port, B2 => pc_target_26_0_port, ZN => n231);
   U303 : INV_X1 port map( A => n232, ZN => n5666);
   U304 : AOI22_X1 port map( A1 => Set_target(1), A2 => n215_port, B1 => 
                           n216_port, B2 => pc_target_26_1_port, ZN => n232);
   U305 : INV_X1 port map( A => n233, ZN => n5667);
   U306 : AOI22_X1 port map( A1 => Set_target(3), A2 => n215_port, B1 => 
                           n216_port, B2 => pc_target_26_3_port, ZN => n233);
   U307 : INV_X1 port map( A => n234, ZN => n5668);
   U308 : AOI22_X1 port map( A1 => Set_target(5), A2 => n215_port, B1 => 
                           n216_port, B2 => pc_target_26_5_port, ZN => n234);
   U309 : INV_X1 port map( A => n235, ZN => n5669);
   U310 : AOI22_X1 port map( A1 => Set_target(7), A2 => n215_port, B1 => 
                           n216_port, B2 => pc_target_26_7_port, ZN => n235);
   U311 : INV_X1 port map( A => n236, ZN => n5670);
   U312 : AOI22_X1 port map( A1 => Set_target(9), A2 => n215_port, B1 => 
                           n216_port, B2 => pc_target_26_9_port, ZN => n236);
   U313 : INV_X1 port map( A => n237, ZN => n5671);
   U314 : AOI22_X1 port map( A1 => Set_target(11), A2 => n215_port, B1 => 
                           n216_port, B2 => pc_target_26_11_port, ZN => n237);
   U315 : INV_X1 port map( A => n238, ZN => n5672);
   U316 : AOI22_X1 port map( A1 => Set_target(13), A2 => n215_port, B1 => 
                           n216_port, B2 => pc_target_26_13_port, ZN => n238);
   U317 : INV_X1 port map( A => n239, ZN => n5673);
   U318 : AOI22_X1 port map( A1 => Set_target(15), A2 => n215_port, B1 => 
                           n216_port, B2 => pc_target_26_15_port, ZN => n239);
   U319 : INV_X1 port map( A => n240, ZN => n5674);
   U320 : AOI22_X1 port map( A1 => Set_target(17), A2 => n215_port, B1 => 
                           n216_port, B2 => pc_target_26_17_port, ZN => n240);
   U321 : INV_X1 port map( A => n241, ZN => n5675);
   U322 : AOI22_X1 port map( A1 => Set_target(19), A2 => n215_port, B1 => 
                           n216_port, B2 => pc_target_26_19_port, ZN => n241);
   U323 : INV_X1 port map( A => n242, ZN => n5676);
   U324 : AOI22_X1 port map( A1 => Set_target(21), A2 => n215_port, B1 => 
                           n216_port, B2 => pc_target_26_21_port, ZN => n242);
   U325 : INV_X1 port map( A => n243, ZN => n5677);
   U326 : AOI22_X1 port map( A1 => Set_target(23), A2 => n215_port, B1 => 
                           n216_port, B2 => pc_target_26_23_port, ZN => n243);
   U327 : INV_X1 port map( A => n244, ZN => n5678);
   U328 : AOI22_X1 port map( A1 => Set_target(25), A2 => n215_port, B1 => 
                           n216_port, B2 => pc_target_26_25_port, ZN => n244);
   U329 : INV_X1 port map( A => n245, ZN => n5679);
   U330 : AOI22_X1 port map( A1 => Set_target(27), A2 => n215_port, B1 => 
                           n216_port, B2 => pc_target_26_27_port, ZN => n245);
   U331 : INV_X1 port map( A => n246, ZN => n5680);
   U332 : AOI22_X1 port map( A1 => Set_target(29), A2 => n215_port, B1 => 
                           n216_port, B2 => pc_target_26_29_port, ZN => n246);
   U333 : INV_X1 port map( A => n247, ZN => n5681);
   U334 : AOI22_X1 port map( A1 => Set_target(31), A2 => n215_port, B1 => 
                           n216_port, B2 => pc_target_26_31_port, ZN => n247);
   U337 : OAI22_X1 port map( A1 => n75, A2 => n248, B1 => n249, B2 => n250, ZN 
                           => n5682);
   U338 : OAI22_X1 port map( A1 => n79, A2 => n248, B1 => n249, B2 => n251, ZN 
                           => n5683);
   U339 : OAI22_X1 port map( A1 => n81, A2 => n248, B1 => n249, B2 => n252, ZN 
                           => n5684);
   U340 : OAI22_X1 port map( A1 => n83, A2 => n248, B1 => n249, B2 => n253, ZN 
                           => n5685);
   U341 : OAI22_X1 port map( A1 => n85, A2 => n248, B1 => n249, B2 => n254, ZN 
                           => n5686);
   U342 : OAI22_X1 port map( A1 => n87, A2 => n248, B1 => n249, B2 => n255, ZN 
                           => n5687);
   U343 : OAI22_X1 port map( A1 => n89, A2 => n248, B1 => n249, B2 => n256, ZN 
                           => n5688);
   U344 : OAI22_X1 port map( A1 => n91, A2 => n248, B1 => n249, B2 => n257, ZN 
                           => n5689);
   U345 : OAI22_X1 port map( A1 => n93, A2 => n248, B1 => n249, B2 => n258, ZN 
                           => n5690);
   U346 : OAI22_X1 port map( A1 => n95, A2 => n248, B1 => n249, B2 => n259, ZN 
                           => n5691);
   U347 : OAI22_X1 port map( A1 => n97_port, A2 => n248, B1 => n249, B2 => n260
                           , ZN => n5692);
   U348 : OAI22_X1 port map( A1 => n99_port, A2 => n248, B1 => n249, B2 => n261
                           , ZN => n5693);
   U349 : OAI22_X1 port map( A1 => n101_port, A2 => n248, B1 => n249, B2 => 
                           n262, ZN => n5694);
   U350 : OAI22_X1 port map( A1 => n103_port, A2 => n248, B1 => n249, B2 => 
                           n263, ZN => n5695);
   U351 : OAI22_X1 port map( A1 => n105_port, A2 => n248, B1 => n249, B2 => 
                           n264, ZN => n5696);
   U352 : OAI22_X1 port map( A1 => n107_port, A2 => n248, B1 => n249, B2 => 
                           n265, ZN => n5697);
   U353 : OAI22_X1 port map( A1 => n109_port, A2 => n248, B1 => n249, B2 => 
                           n266, ZN => n5698);
   U354 : OAI22_X1 port map( A1 => n111_port, A2 => n248, B1 => n249, B2 => 
                           n267, ZN => n5699);
   U355 : OAI22_X1 port map( A1 => n113_port, A2 => n248, B1 => n249, B2 => 
                           n268, ZN => n5700);
   U356 : OAI22_X1 port map( A1 => n115_port, A2 => n248, B1 => n249, B2 => 
                           n269, ZN => n5701);
   U357 : OAI22_X1 port map( A1 => n117_port, A2 => n248, B1 => n249, B2 => 
                           n270, ZN => n5702);
   U358 : OAI22_X1 port map( A1 => n119_port, A2 => n248, B1 => n249, B2 => 
                           n271, ZN => n5703);
   U359 : OAI22_X1 port map( A1 => n121_port, A2 => n248, B1 => n249, B2 => 
                           n272, ZN => n5704);
   U360 : OAI22_X1 port map( A1 => n123_port, A2 => n248, B1 => n249, B2 => 
                           n273, ZN => n5705);
   U361 : OAI22_X1 port map( A1 => n125_port, A2 => n248, B1 => n249, B2 => 
                           n274, ZN => n5706);
   U362 : OAI22_X1 port map( A1 => n127_port, A2 => n248, B1 => n249, B2 => 
                           n275, ZN => n5707);
   U363 : OAI22_X1 port map( A1 => n129, A2 => n248, B1 => n249, B2 => n276, ZN
                           => n5708);
   U364 : OAI22_X1 port map( A1 => n131, A2 => n248, B1 => n249, B2 => n277, ZN
                           => n5709);
   U365 : OAI22_X1 port map( A1 => n133, A2 => n248, B1 => n249, B2 => n278, ZN
                           => n5710);
   U366 : OAI22_X1 port map( A1 => n135, A2 => n248, B1 => n249, B2 => n279, ZN
                           => n5711);
   U367 : OAI22_X1 port map( A1 => n137, A2 => n248, B1 => n249, B2 => n280, ZN
                           => n5712);
   U368 : OAI22_X1 port map( A1 => n139, A2 => n248, B1 => n249, B2 => n281, ZN
                           => n5713);
   U371 : OAI22_X1 port map( A1 => n75, A2 => n282, B1 => n3444, B2 => n284, ZN
                           => n5714);
   U372 : OAI22_X1 port map( A1 => n79, A2 => n282, B1 => n3444, B2 => n285, ZN
                           => n5715);
   U373 : OAI22_X1 port map( A1 => n81, A2 => n282, B1 => n3444, B2 => n286, ZN
                           => n5716);
   U374 : OAI22_X1 port map( A1 => n83, A2 => n282, B1 => n3444, B2 => n287, ZN
                           => n5717);
   U375 : OAI22_X1 port map( A1 => n85, A2 => n282, B1 => n3444, B2 => n288, ZN
                           => n5718);
   U376 : OAI22_X1 port map( A1 => n87, A2 => n282, B1 => n3444, B2 => n289, ZN
                           => n5719);
   U377 : OAI22_X1 port map( A1 => n89, A2 => n282, B1 => n3444, B2 => n290, ZN
                           => n5720);
   U378 : OAI22_X1 port map( A1 => n91, A2 => n282, B1 => n3444, B2 => n291, ZN
                           => n5721);
   U379 : OAI22_X1 port map( A1 => n93, A2 => n282, B1 => n3444, B2 => n292, ZN
                           => n5722);
   U380 : OAI22_X1 port map( A1 => n95, A2 => n282, B1 => n3444, B2 => n293, ZN
                           => n5723);
   U381 : OAI22_X1 port map( A1 => n97_port, A2 => n282, B1 => n3444, B2 => 
                           n294, ZN => n5724);
   U382 : OAI22_X1 port map( A1 => n99_port, A2 => n282, B1 => n3444, B2 => 
                           n295, ZN => n5725);
   U383 : OAI22_X1 port map( A1 => n101_port, A2 => n282, B1 => n3444, B2 => 
                           n296, ZN => n5726);
   U384 : OAI22_X1 port map( A1 => n103_port, A2 => n282, B1 => n3444, B2 => 
                           n297, ZN => n5727);
   U385 : OAI22_X1 port map( A1 => n105_port, A2 => n282, B1 => n3444, B2 => 
                           n298, ZN => n5728);
   U386 : OAI22_X1 port map( A1 => n107_port, A2 => n282, B1 => n3444, B2 => 
                           n299, ZN => n5729);
   U387 : OAI22_X1 port map( A1 => n109_port, A2 => n282, B1 => n3444, B2 => 
                           n300, ZN => n5730);
   U388 : OAI22_X1 port map( A1 => n111_port, A2 => n282, B1 => n3444, B2 => 
                           n301, ZN => n5731);
   U389 : OAI22_X1 port map( A1 => n113_port, A2 => n282, B1 => n3444, B2 => 
                           n302, ZN => n5732);
   U390 : OAI22_X1 port map( A1 => n115_port, A2 => n282, B1 => n3444, B2 => 
                           n303, ZN => n5733);
   U391 : OAI22_X1 port map( A1 => n117_port, A2 => n282, B1 => n3444, B2 => 
                           n304, ZN => n5734);
   U392 : OAI22_X1 port map( A1 => n119_port, A2 => n282, B1 => n3444, B2 => 
                           n305, ZN => n5735);
   U393 : OAI22_X1 port map( A1 => n121_port, A2 => n282, B1 => n3444, B2 => 
                           n306, ZN => n5736);
   U394 : OAI22_X1 port map( A1 => n123_port, A2 => n282, B1 => n3444, B2 => 
                           n307, ZN => n5737);
   U395 : OAI22_X1 port map( A1 => n125_port, A2 => n282, B1 => n3444, B2 => 
                           n308, ZN => n5738);
   U396 : OAI22_X1 port map( A1 => n127_port, A2 => n282, B1 => n3444, B2 => 
                           n309, ZN => n5739);
   U397 : OAI22_X1 port map( A1 => n129, A2 => n282, B1 => n3444, B2 => n310, 
                           ZN => n5740);
   U398 : OAI22_X1 port map( A1 => n131, A2 => n282, B1 => n3444, B2 => n311, 
                           ZN => n5741);
   U399 : OAI22_X1 port map( A1 => n133, A2 => n282, B1 => n3444, B2 => n312, 
                           ZN => n5742);
   U400 : OAI22_X1 port map( A1 => n135, A2 => n282, B1 => n3444, B2 => n313, 
                           ZN => n5743);
   U401 : OAI22_X1 port map( A1 => n137, A2 => n282, B1 => n3444, B2 => n314, 
                           ZN => n5744);
   U402 : OAI22_X1 port map( A1 => n139, A2 => n282, B1 => n3444, B2 => n315, 
                           ZN => n5745);
   U406 : OAI22_X1 port map( A1 => n75, A2 => n317, B1 => n318, B2 => n319, ZN 
                           => n5746);
   U407 : OAI22_X1 port map( A1 => n79, A2 => n317, B1 => n318, B2 => n320, ZN 
                           => n5747);
   U408 : OAI22_X1 port map( A1 => n81, A2 => n317, B1 => n318, B2 => n321, ZN 
                           => n5748);
   U409 : OAI22_X1 port map( A1 => n83, A2 => n317, B1 => n318, B2 => n322, ZN 
                           => n5749);
   U410 : OAI22_X1 port map( A1 => n85, A2 => n317, B1 => n318, B2 => n323, ZN 
                           => n5750);
   U411 : OAI22_X1 port map( A1 => n87, A2 => n317, B1 => n318, B2 => n324, ZN 
                           => n5751);
   U412 : OAI22_X1 port map( A1 => n89, A2 => n317, B1 => n318, B2 => n325, ZN 
                           => n5752);
   U413 : OAI22_X1 port map( A1 => n91, A2 => n317, B1 => n318, B2 => n326, ZN 
                           => n5753);
   U414 : OAI22_X1 port map( A1 => n93, A2 => n317, B1 => n318, B2 => n327, ZN 
                           => n5754);
   U415 : OAI22_X1 port map( A1 => n95, A2 => n317, B1 => n318, B2 => n328, ZN 
                           => n5755);
   U416 : OAI22_X1 port map( A1 => n97_port, A2 => n317, B1 => n318, B2 => n329
                           , ZN => n5756);
   U417 : OAI22_X1 port map( A1 => n99_port, A2 => n317, B1 => n318, B2 => n330
                           , ZN => n5757);
   U418 : OAI22_X1 port map( A1 => n101_port, A2 => n317, B1 => n318, B2 => 
                           n331, ZN => n5758);
   U419 : OAI22_X1 port map( A1 => n103_port, A2 => n317, B1 => n318, B2 => 
                           n332, ZN => n5759);
   U420 : OAI22_X1 port map( A1 => n105_port, A2 => n317, B1 => n318, B2 => 
                           n333, ZN => n5760);
   U421 : OAI22_X1 port map( A1 => n107_port, A2 => n317, B1 => n318, B2 => 
                           n334, ZN => n5761);
   U422 : OAI22_X1 port map( A1 => n109_port, A2 => n317, B1 => n318, B2 => 
                           n335, ZN => n5762);
   U423 : OAI22_X1 port map( A1 => n111_port, A2 => n317, B1 => n318, B2 => 
                           n336, ZN => n5763);
   U424 : OAI22_X1 port map( A1 => n113_port, A2 => n317, B1 => n318, B2 => 
                           n337, ZN => n5764);
   U425 : OAI22_X1 port map( A1 => n115_port, A2 => n317, B1 => n318, B2 => 
                           n338, ZN => n5765);
   U426 : OAI22_X1 port map( A1 => n117_port, A2 => n317, B1 => n318, B2 => 
                           n339, ZN => n5766);
   U427 : OAI22_X1 port map( A1 => n119_port, A2 => n317, B1 => n318, B2 => 
                           n340, ZN => n5767);
   U428 : OAI22_X1 port map( A1 => n121_port, A2 => n317, B1 => n318, B2 => 
                           n341, ZN => n5768);
   U429 : OAI22_X1 port map( A1 => n123_port, A2 => n317, B1 => n318, B2 => 
                           n342, ZN => n5769);
   U430 : OAI22_X1 port map( A1 => n125_port, A2 => n317, B1 => n318, B2 => 
                           n343, ZN => n5770);
   U431 : OAI22_X1 port map( A1 => n127_port, A2 => n317, B1 => n318, B2 => 
                           n344, ZN => n5771);
   U432 : OAI22_X1 port map( A1 => n129, A2 => n317, B1 => n318, B2 => n345, ZN
                           => n5772);
   U433 : OAI22_X1 port map( A1 => n131, A2 => n317, B1 => n318, B2 => n346, ZN
                           => n5773);
   U434 : OAI22_X1 port map( A1 => n133, A2 => n317, B1 => n318, B2 => n347, ZN
                           => n5774);
   U435 : OAI22_X1 port map( A1 => n135, A2 => n317, B1 => n318, B2 => n348, ZN
                           => n5775);
   U436 : OAI22_X1 port map( A1 => n137, A2 => n317, B1 => n318, B2 => n349, ZN
                           => n5776);
   U437 : OAI22_X1 port map( A1 => n139, A2 => n317, B1 => n318, B2 => n350, ZN
                           => n5777);
   U440 : OAI22_X1 port map( A1 => n75, A2 => n352, B1 => n353, B2 => n354, ZN 
                           => n5778);
   U441 : OAI22_X1 port map( A1 => n79, A2 => n352, B1 => n353, B2 => n355, ZN 
                           => n5779);
   U442 : OAI22_X1 port map( A1 => n81, A2 => n352, B1 => n353, B2 => n356, ZN 
                           => n5780);
   U443 : OAI22_X1 port map( A1 => n83, A2 => n352, B1 => n353, B2 => n357, ZN 
                           => n5781);
   U444 : OAI22_X1 port map( A1 => n85, A2 => n352, B1 => n353, B2 => n358, ZN 
                           => n5782);
   U445 : OAI22_X1 port map( A1 => n87, A2 => n352, B1 => n353, B2 => n359, ZN 
                           => n5783);
   U446 : OAI22_X1 port map( A1 => n89, A2 => n352, B1 => n353, B2 => n360, ZN 
                           => n5784);
   U447 : OAI22_X1 port map( A1 => n91, A2 => n352, B1 => n353, B2 => n361, ZN 
                           => n5785);
   U448 : OAI22_X1 port map( A1 => n93, A2 => n352, B1 => n353, B2 => n362, ZN 
                           => n5786);
   U449 : OAI22_X1 port map( A1 => n95, A2 => n352, B1 => n353, B2 => n363, ZN 
                           => n5787);
   U450 : OAI22_X1 port map( A1 => n97_port, A2 => n352, B1 => n353, B2 => n364
                           , ZN => n5788);
   U451 : OAI22_X1 port map( A1 => n99_port, A2 => n352, B1 => n353, B2 => n365
                           , ZN => n5789);
   U452 : OAI22_X1 port map( A1 => n101_port, A2 => n352, B1 => n353, B2 => 
                           n366, ZN => n5790);
   U453 : OAI22_X1 port map( A1 => n103_port, A2 => n352, B1 => n353, B2 => 
                           n367, ZN => n5791);
   U454 : OAI22_X1 port map( A1 => n105_port, A2 => n352, B1 => n353, B2 => 
                           n368, ZN => n5792);
   U455 : OAI22_X1 port map( A1 => n107_port, A2 => n352, B1 => n353, B2 => 
                           n369, ZN => n5793);
   U456 : OAI22_X1 port map( A1 => n109_port, A2 => n352, B1 => n353, B2 => 
                           n370, ZN => n5794);
   U457 : OAI22_X1 port map( A1 => n111_port, A2 => n352, B1 => n353, B2 => 
                           n371, ZN => n5795);
   U458 : OAI22_X1 port map( A1 => n113_port, A2 => n352, B1 => n353, B2 => 
                           n372, ZN => n5796);
   U459 : OAI22_X1 port map( A1 => n115_port, A2 => n352, B1 => n353, B2 => 
                           n373, ZN => n5797);
   U460 : OAI22_X1 port map( A1 => n117_port, A2 => n352, B1 => n353, B2 => 
                           n374, ZN => n5798);
   U461 : OAI22_X1 port map( A1 => n119_port, A2 => n352, B1 => n353, B2 => 
                           n375, ZN => n5799);
   U462 : OAI22_X1 port map( A1 => n121_port, A2 => n352, B1 => n353, B2 => 
                           n376, ZN => n5800);
   U463 : OAI22_X1 port map( A1 => n123_port, A2 => n352, B1 => n353, B2 => 
                           n377, ZN => n5801);
   U464 : OAI22_X1 port map( A1 => n125_port, A2 => n352, B1 => n353, B2 => 
                           n378, ZN => n5802);
   U465 : OAI22_X1 port map( A1 => n127_port, A2 => n352, B1 => n353, B2 => 
                           n379, ZN => n5803);
   U466 : OAI22_X1 port map( A1 => n129, A2 => n352, B1 => n353, B2 => n380, ZN
                           => n5804);
   U467 : OAI22_X1 port map( A1 => n131, A2 => n352, B1 => n353, B2 => n381, ZN
                           => n5805);
   U468 : OAI22_X1 port map( A1 => n133, A2 => n352, B1 => n353, B2 => n382, ZN
                           => n5806);
   U469 : OAI22_X1 port map( A1 => n135, A2 => n352, B1 => n353, B2 => n383, ZN
                           => n5807);
   U470 : OAI22_X1 port map( A1 => n137, A2 => n352, B1 => n353, B2 => n384, ZN
                           => n5808);
   U471 : OAI22_X1 port map( A1 => n139, A2 => n352, B1 => n353, B2 => n385, ZN
                           => n5809);
   U474 : INV_X1 port map( A => n386, ZN => n5810);
   U475 : AOI22_X1 port map( A1 => Set_target(30), A2 => n3799, B1 => n388, B2 
                           => pc_target_21_30_port, ZN => n386);
   U476 : INV_X1 port map( A => n389, ZN => n5811);
   U477 : AOI22_X1 port map( A1 => Set_target(28), A2 => n3799, B1 => n388, B2 
                           => pc_target_21_28_port, ZN => n389);
   U478 : INV_X1 port map( A => n390, ZN => n5812);
   U479 : AOI22_X1 port map( A1 => Set_target(26), A2 => n3799, B1 => n388, B2 
                           => pc_target_21_26_port, ZN => n390);
   U480 : INV_X1 port map( A => n391, ZN => n5813);
   U481 : AOI22_X1 port map( A1 => Set_target(24), A2 => n3799, B1 => n388, B2 
                           => pc_target_21_24_port, ZN => n391);
   U482 : INV_X1 port map( A => n392, ZN => n5814);
   U483 : AOI22_X1 port map( A1 => Set_target(22), A2 => n3799, B1 => n388, B2 
                           => pc_target_21_22_port, ZN => n392);
   U484 : INV_X1 port map( A => n393, ZN => n5815);
   U485 : AOI22_X1 port map( A1 => Set_target(20), A2 => n3799, B1 => n388, B2 
                           => pc_target_21_20_port, ZN => n393);
   U486 : INV_X1 port map( A => n394, ZN => n5816);
   U487 : AOI22_X1 port map( A1 => Set_target(18), A2 => n3799, B1 => n388, B2 
                           => pc_target_21_18_port, ZN => n394);
   U488 : INV_X1 port map( A => n395, ZN => n5817);
   U489 : AOI22_X1 port map( A1 => Set_target(16), A2 => n3799, B1 => n388, B2 
                           => pc_target_21_16_port, ZN => n395);
   U490 : INV_X1 port map( A => n396, ZN => n5818);
   U491 : AOI22_X1 port map( A1 => Set_target(14), A2 => n3799, B1 => n388, B2 
                           => pc_target_21_14_port, ZN => n396);
   U492 : INV_X1 port map( A => n397, ZN => n5819);
   U493 : AOI22_X1 port map( A1 => Set_target(12), A2 => n3799, B1 => n388, B2 
                           => pc_target_21_12_port, ZN => n397);
   U494 : INV_X1 port map( A => n398, ZN => n5820);
   U495 : AOI22_X1 port map( A1 => Set_target(10), A2 => n3799, B1 => n388, B2 
                           => pc_target_21_10_port, ZN => n398);
   U496 : INV_X1 port map( A => n399, ZN => n5821);
   U497 : AOI22_X1 port map( A1 => Set_target(8), A2 => n3799, B1 => n388, B2 
                           => pc_target_21_8_port, ZN => n399);
   U498 : INV_X1 port map( A => n400, ZN => n5822);
   U499 : AOI22_X1 port map( A1 => Set_target(6), A2 => n3799, B1 => n388, B2 
                           => pc_target_21_6_port, ZN => n400);
   U500 : INV_X1 port map( A => n401, ZN => n5823);
   U501 : AOI22_X1 port map( A1 => Set_target(4), A2 => n3799, B1 => n388, B2 
                           => pc_target_21_4_port, ZN => n401);
   U502 : INV_X1 port map( A => n402, ZN => n5824);
   U503 : AOI22_X1 port map( A1 => Set_target(2), A2 => n3799, B1 => n388, B2 
                           => pc_target_21_2_port, ZN => n402);
   U504 : INV_X1 port map( A => n403, ZN => n5825);
   U505 : AOI22_X1 port map( A1 => Set_target(0), A2 => n3799, B1 => n388, B2 
                           => pc_target_21_0_port, ZN => n403);
   U506 : INV_X1 port map( A => n404, ZN => n5826);
   U507 : AOI22_X1 port map( A1 => Set_target(1), A2 => n3799, B1 => n388, B2 
                           => pc_target_21_1_port, ZN => n404);
   U508 : INV_X1 port map( A => n405, ZN => n5827);
   U509 : AOI22_X1 port map( A1 => Set_target(3), A2 => n3799, B1 => n388, B2 
                           => pc_target_21_3_port, ZN => n405);
   U510 : INV_X1 port map( A => n406, ZN => n5828);
   U511 : AOI22_X1 port map( A1 => Set_target(5), A2 => n3799, B1 => n388, B2 
                           => pc_target_21_5_port, ZN => n406);
   U512 : INV_X1 port map( A => n407, ZN => n5829);
   U513 : AOI22_X1 port map( A1 => Set_target(7), A2 => n3799, B1 => n388, B2 
                           => pc_target_21_7_port, ZN => n407);
   U514 : INV_X1 port map( A => n408, ZN => n5830);
   U515 : AOI22_X1 port map( A1 => Set_target(9), A2 => n3799, B1 => n388, B2 
                           => pc_target_21_9_port, ZN => n408);
   U516 : INV_X1 port map( A => n409, ZN => n5831);
   U517 : AOI22_X1 port map( A1 => Set_target(11), A2 => n3799, B1 => n388, B2 
                           => pc_target_21_11_port, ZN => n409);
   U518 : INV_X1 port map( A => n410, ZN => n5832);
   U519 : AOI22_X1 port map( A1 => Set_target(13), A2 => n3799, B1 => n388, B2 
                           => pc_target_21_13_port, ZN => n410);
   U520 : INV_X1 port map( A => n411, ZN => n5833);
   U521 : AOI22_X1 port map( A1 => Set_target(15), A2 => n3799, B1 => n388, B2 
                           => pc_target_21_15_port, ZN => n411);
   U522 : INV_X1 port map( A => n412, ZN => n5834);
   U523 : AOI22_X1 port map( A1 => Set_target(17), A2 => n3799, B1 => n388, B2 
                           => pc_target_21_17_port, ZN => n412);
   U524 : INV_X1 port map( A => n413, ZN => n5835);
   U525 : AOI22_X1 port map( A1 => Set_target(19), A2 => n3799, B1 => n388, B2 
                           => pc_target_21_19_port, ZN => n413);
   U526 : INV_X1 port map( A => n414, ZN => n5836);
   U527 : AOI22_X1 port map( A1 => Set_target(21), A2 => n3799, B1 => n388, B2 
                           => pc_target_21_21_port, ZN => n414);
   U528 : INV_X1 port map( A => n415, ZN => n5837);
   U529 : AOI22_X1 port map( A1 => Set_target(23), A2 => n3799, B1 => n388, B2 
                           => pc_target_21_23_port, ZN => n415);
   U530 : INV_X1 port map( A => n416, ZN => n5838);
   U531 : AOI22_X1 port map( A1 => Set_target(25), A2 => n3799, B1 => n388, B2 
                           => pc_target_21_25_port, ZN => n416);
   U532 : INV_X1 port map( A => n417, ZN => n5839);
   U533 : AOI22_X1 port map( A1 => Set_target(27), A2 => n3799, B1 => n388, B2 
                           => pc_target_21_27_port, ZN => n417);
   U534 : INV_X1 port map( A => n418, ZN => n5840);
   U535 : AOI22_X1 port map( A1 => Set_target(29), A2 => n3799, B1 => n388, B2 
                           => pc_target_21_29_port, ZN => n418);
   U536 : INV_X1 port map( A => n419, ZN => n5841);
   U537 : AOI22_X1 port map( A1 => Set_target(31), A2 => n3799, B1 => n388, B2 
                           => pc_target_21_31_port, ZN => n419);
   U540 : INV_X1 port map( A => n420, ZN => n5842);
   U541 : AOI22_X1 port map( A1 => Set_target(30), A2 => n421, B1 => n422, B2 
                           => pc_target_20_30_port, ZN => n420);
   U542 : INV_X1 port map( A => n423, ZN => n5843);
   U543 : AOI22_X1 port map( A1 => Set_target(28), A2 => n421, B1 => n422, B2 
                           => pc_target_20_28_port, ZN => n423);
   U544 : INV_X1 port map( A => n424, ZN => n5844);
   U545 : AOI22_X1 port map( A1 => Set_target(26), A2 => n421, B1 => n422, B2 
                           => pc_target_20_26_port, ZN => n424);
   U546 : INV_X1 port map( A => n425, ZN => n5845);
   U547 : AOI22_X1 port map( A1 => Set_target(24), A2 => n421, B1 => n422, B2 
                           => pc_target_20_24_port, ZN => n425);
   U548 : INV_X1 port map( A => n426, ZN => n5846);
   U549 : AOI22_X1 port map( A1 => Set_target(22), A2 => n421, B1 => n422, B2 
                           => pc_target_20_22_port, ZN => n426);
   U550 : INV_X1 port map( A => n427, ZN => n5847);
   U551 : AOI22_X1 port map( A1 => Set_target(20), A2 => n421, B1 => n422, B2 
                           => pc_target_20_20_port, ZN => n427);
   U552 : INV_X1 port map( A => n428, ZN => n5848);
   U553 : AOI22_X1 port map( A1 => Set_target(18), A2 => n421, B1 => n422, B2 
                           => pc_target_20_18_port, ZN => n428);
   U554 : INV_X1 port map( A => n429, ZN => n5849);
   U555 : AOI22_X1 port map( A1 => Set_target(16), A2 => n421, B1 => n422, B2 
                           => pc_target_20_16_port, ZN => n429);
   U556 : INV_X1 port map( A => n430, ZN => n5850);
   U557 : AOI22_X1 port map( A1 => Set_target(14), A2 => n421, B1 => n422, B2 
                           => pc_target_20_14_port, ZN => n430);
   U558 : INV_X1 port map( A => n431, ZN => n5851);
   U559 : AOI22_X1 port map( A1 => Set_target(12), A2 => n421, B1 => n422, B2 
                           => pc_target_20_12_port, ZN => n431);
   U560 : INV_X1 port map( A => n432, ZN => n5852);
   U561 : AOI22_X1 port map( A1 => Set_target(10), A2 => n421, B1 => n422, B2 
                           => pc_target_20_10_port, ZN => n432);
   U562 : INV_X1 port map( A => n433, ZN => n5853);
   U563 : AOI22_X1 port map( A1 => Set_target(8), A2 => n421, B1 => n422, B2 =>
                           pc_target_20_8_port, ZN => n433);
   U564 : INV_X1 port map( A => n434, ZN => n5854);
   U565 : AOI22_X1 port map( A1 => Set_target(6), A2 => n421, B1 => n422, B2 =>
                           pc_target_20_6_port, ZN => n434);
   U566 : INV_X1 port map( A => n435, ZN => n5855);
   U567 : AOI22_X1 port map( A1 => Set_target(4), A2 => n421, B1 => n422, B2 =>
                           pc_target_20_4_port, ZN => n435);
   U568 : INV_X1 port map( A => n436, ZN => n5856);
   U569 : AOI22_X1 port map( A1 => Set_target(2), A2 => n421, B1 => n422, B2 =>
                           pc_target_20_2_port, ZN => n436);
   U570 : INV_X1 port map( A => n437, ZN => n5857);
   U571 : AOI22_X1 port map( A1 => Set_target(0), A2 => n421, B1 => n422, B2 =>
                           pc_target_20_0_port, ZN => n437);
   U572 : INV_X1 port map( A => n438, ZN => n5858);
   U573 : AOI22_X1 port map( A1 => Set_target(1), A2 => n421, B1 => n422, B2 =>
                           pc_target_20_1_port, ZN => n438);
   U574 : INV_X1 port map( A => n439, ZN => n5859);
   U575 : AOI22_X1 port map( A1 => Set_target(3), A2 => n421, B1 => n422, B2 =>
                           pc_target_20_3_port, ZN => n439);
   U576 : INV_X1 port map( A => n440, ZN => n5860);
   U577 : AOI22_X1 port map( A1 => Set_target(5), A2 => n421, B1 => n422, B2 =>
                           pc_target_20_5_port, ZN => n440);
   U578 : INV_X1 port map( A => n441, ZN => n5861);
   U579 : AOI22_X1 port map( A1 => Set_target(7), A2 => n421, B1 => n422, B2 =>
                           pc_target_20_7_port, ZN => n441);
   U580 : INV_X1 port map( A => n442, ZN => n5862);
   U581 : AOI22_X1 port map( A1 => Set_target(9), A2 => n421, B1 => n422, B2 =>
                           pc_target_20_9_port, ZN => n442);
   U582 : INV_X1 port map( A => n443, ZN => n5863);
   U583 : AOI22_X1 port map( A1 => Set_target(11), A2 => n421, B1 => n422, B2 
                           => pc_target_20_11_port, ZN => n443);
   U584 : INV_X1 port map( A => n444, ZN => n5864);
   U585 : AOI22_X1 port map( A1 => Set_target(13), A2 => n421, B1 => n422, B2 
                           => pc_target_20_13_port, ZN => n444);
   U586 : INV_X1 port map( A => n445, ZN => n5865);
   U587 : AOI22_X1 port map( A1 => Set_target(15), A2 => n421, B1 => n422, B2 
                           => pc_target_20_15_port, ZN => n445);
   U588 : INV_X1 port map( A => n446, ZN => n5866);
   U589 : AOI22_X1 port map( A1 => Set_target(17), A2 => n421, B1 => n422, B2 
                           => pc_target_20_17_port, ZN => n446);
   U590 : INV_X1 port map( A => n447, ZN => n5867);
   U591 : AOI22_X1 port map( A1 => Set_target(19), A2 => n421, B1 => n422, B2 
                           => pc_target_20_19_port, ZN => n447);
   U592 : INV_X1 port map( A => n448, ZN => n5868);
   U593 : AOI22_X1 port map( A1 => Set_target(21), A2 => n421, B1 => n422, B2 
                           => pc_target_20_21_port, ZN => n448);
   U594 : INV_X1 port map( A => n449, ZN => n5869);
   U595 : AOI22_X1 port map( A1 => Set_target(23), A2 => n421, B1 => n422, B2 
                           => pc_target_20_23_port, ZN => n449);
   U596 : INV_X1 port map( A => n450, ZN => n5870);
   U597 : AOI22_X1 port map( A1 => Set_target(25), A2 => n421, B1 => n422, B2 
                           => pc_target_20_25_port, ZN => n450);
   U598 : INV_X1 port map( A => n451, ZN => n5871);
   U599 : AOI22_X1 port map( A1 => Set_target(27), A2 => n421, B1 => n422, B2 
                           => pc_target_20_27_port, ZN => n451);
   U600 : INV_X1 port map( A => n452, ZN => n5872);
   U601 : AOI22_X1 port map( A1 => Set_target(29), A2 => n421, B1 => n422, B2 
                           => pc_target_20_29_port, ZN => n452);
   U602 : INV_X1 port map( A => n453, ZN => n5873);
   U603 : AOI22_X1 port map( A1 => Set_target(31), A2 => n421, B1 => n422, B2 
                           => pc_target_20_31_port, ZN => n453);
   U607 : INV_X1 port map( A => n455, ZN => n5874);
   U608 : AOI22_X1 port map( A1 => Set_target(30), A2 => n456, B1 => n457, B2 
                           => pc_target_19_30_port, ZN => n455);
   U609 : INV_X1 port map( A => n458, ZN => n5875);
   U610 : AOI22_X1 port map( A1 => Set_target(28), A2 => n456, B1 => n457, B2 
                           => pc_target_19_28_port, ZN => n458);
   U611 : INV_X1 port map( A => n459, ZN => n5876);
   U612 : AOI22_X1 port map( A1 => Set_target(26), A2 => n456, B1 => n457, B2 
                           => pc_target_19_26_port, ZN => n459);
   U613 : INV_X1 port map( A => n460, ZN => n5877);
   U614 : AOI22_X1 port map( A1 => Set_target(24), A2 => n456, B1 => n457, B2 
                           => pc_target_19_24_port, ZN => n460);
   U615 : INV_X1 port map( A => n461, ZN => n5878);
   U616 : AOI22_X1 port map( A1 => Set_target(22), A2 => n456, B1 => n457, B2 
                           => pc_target_19_22_port, ZN => n461);
   U617 : INV_X1 port map( A => n462, ZN => n5879);
   U618 : AOI22_X1 port map( A1 => Set_target(20), A2 => n456, B1 => n457, B2 
                           => pc_target_19_20_port, ZN => n462);
   U619 : INV_X1 port map( A => n463, ZN => n5880);
   U620 : AOI22_X1 port map( A1 => Set_target(18), A2 => n456, B1 => n457, B2 
                           => pc_target_19_18_port, ZN => n463);
   U621 : INV_X1 port map( A => n464, ZN => n5881);
   U622 : AOI22_X1 port map( A1 => Set_target(16), A2 => n456, B1 => n457, B2 
                           => pc_target_19_16_port, ZN => n464);
   U623 : INV_X1 port map( A => n465, ZN => n5882);
   U624 : AOI22_X1 port map( A1 => Set_target(14), A2 => n456, B1 => n457, B2 
                           => pc_target_19_14_port, ZN => n465);
   U625 : INV_X1 port map( A => n466, ZN => n5883);
   U626 : AOI22_X1 port map( A1 => Set_target(12), A2 => n456, B1 => n457, B2 
                           => pc_target_19_12_port, ZN => n466);
   U627 : INV_X1 port map( A => n467, ZN => n5884);
   U628 : AOI22_X1 port map( A1 => Set_target(10), A2 => n456, B1 => n457, B2 
                           => pc_target_19_10_port, ZN => n467);
   U629 : INV_X1 port map( A => n468, ZN => n5885);
   U630 : AOI22_X1 port map( A1 => Set_target(8), A2 => n456, B1 => n457, B2 =>
                           pc_target_19_8_port, ZN => n468);
   U631 : INV_X1 port map( A => n469, ZN => n5886);
   U632 : AOI22_X1 port map( A1 => Set_target(6), A2 => n456, B1 => n457, B2 =>
                           pc_target_19_6_port, ZN => n469);
   U633 : INV_X1 port map( A => n470, ZN => n5887);
   U634 : AOI22_X1 port map( A1 => Set_target(4), A2 => n456, B1 => n457, B2 =>
                           pc_target_19_4_port, ZN => n470);
   U635 : INV_X1 port map( A => n471, ZN => n5888);
   U636 : AOI22_X1 port map( A1 => Set_target(2), A2 => n456, B1 => n457, B2 =>
                           pc_target_19_2_port, ZN => n471);
   U637 : INV_X1 port map( A => n472, ZN => n5889);
   U638 : AOI22_X1 port map( A1 => Set_target(0), A2 => n456, B1 => n457, B2 =>
                           pc_target_19_0_port, ZN => n472);
   U639 : INV_X1 port map( A => n473, ZN => n5890);
   U640 : AOI22_X1 port map( A1 => Set_target(1), A2 => n456, B1 => n457, B2 =>
                           pc_target_19_1_port, ZN => n473);
   U641 : INV_X1 port map( A => n474, ZN => n5891);
   U642 : AOI22_X1 port map( A1 => Set_target(3), A2 => n456, B1 => n457, B2 =>
                           pc_target_19_3_port, ZN => n474);
   U643 : INV_X1 port map( A => n475, ZN => n5892);
   U644 : AOI22_X1 port map( A1 => Set_target(5), A2 => n456, B1 => n457, B2 =>
                           pc_target_19_5_port, ZN => n475);
   U645 : INV_X1 port map( A => n476, ZN => n5893);
   U646 : AOI22_X1 port map( A1 => Set_target(7), A2 => n456, B1 => n457, B2 =>
                           pc_target_19_7_port, ZN => n476);
   U647 : INV_X1 port map( A => n477, ZN => n5894);
   U648 : AOI22_X1 port map( A1 => Set_target(9), A2 => n456, B1 => n457, B2 =>
                           pc_target_19_9_port, ZN => n477);
   U649 : INV_X1 port map( A => n478, ZN => n5895);
   U650 : AOI22_X1 port map( A1 => Set_target(11), A2 => n456, B1 => n457, B2 
                           => pc_target_19_11_port, ZN => n478);
   U651 : INV_X1 port map( A => n479, ZN => n5896);
   U652 : AOI22_X1 port map( A1 => Set_target(13), A2 => n456, B1 => n457, B2 
                           => pc_target_19_13_port, ZN => n479);
   U653 : INV_X1 port map( A => n480, ZN => n5897);
   U654 : AOI22_X1 port map( A1 => Set_target(15), A2 => n456, B1 => n457, B2 
                           => pc_target_19_15_port, ZN => n480);
   U655 : INV_X1 port map( A => n481, ZN => n5898);
   U656 : AOI22_X1 port map( A1 => Set_target(17), A2 => n456, B1 => n457, B2 
                           => pc_target_19_17_port, ZN => n481);
   U657 : INV_X1 port map( A => n482, ZN => n5899);
   U658 : AOI22_X1 port map( A1 => Set_target(19), A2 => n456, B1 => n457, B2 
                           => pc_target_19_19_port, ZN => n482);
   U659 : INV_X1 port map( A => n483, ZN => n5900);
   U660 : AOI22_X1 port map( A1 => Set_target(21), A2 => n456, B1 => n457, B2 
                           => pc_target_19_21_port, ZN => n483);
   U661 : INV_X1 port map( A => n484, ZN => n5901);
   U662 : AOI22_X1 port map( A1 => Set_target(23), A2 => n456, B1 => n457, B2 
                           => pc_target_19_23_port, ZN => n484);
   U663 : INV_X1 port map( A => n485, ZN => n5902);
   U664 : AOI22_X1 port map( A1 => Set_target(25), A2 => n456, B1 => n457, B2 
                           => pc_target_19_25_port, ZN => n485);
   U665 : INV_X1 port map( A => n486, ZN => n5903);
   U666 : AOI22_X1 port map( A1 => Set_target(27), A2 => n456, B1 => n457, B2 
                           => pc_target_19_27_port, ZN => n486);
   U667 : INV_X1 port map( A => n487, ZN => n5904);
   U668 : AOI22_X1 port map( A1 => Set_target(29), A2 => n456, B1 => n457, B2 
                           => pc_target_19_29_port, ZN => n487);
   U669 : INV_X1 port map( A => n488, ZN => n5905);
   U670 : AOI22_X1 port map( A1 => Set_target(31), A2 => n456, B1 => n457, B2 
                           => pc_target_19_31_port, ZN => n488);
   U673 : INV_X1 port map( A => n490, ZN => n5906);
   U674 : AOI22_X1 port map( A1 => Set_target(30), A2 => n491, B1 => n492, B2 
                           => pc_target_18_30_port, ZN => n490);
   U675 : INV_X1 port map( A => n493, ZN => n5907);
   U676 : AOI22_X1 port map( A1 => Set_target(28), A2 => n491, B1 => n492, B2 
                           => pc_target_18_28_port, ZN => n493);
   U677 : INV_X1 port map( A => n494, ZN => n5908);
   U678 : AOI22_X1 port map( A1 => Set_target(26), A2 => n491, B1 => n492, B2 
                           => pc_target_18_26_port, ZN => n494);
   U679 : INV_X1 port map( A => n495, ZN => n5909);
   U680 : AOI22_X1 port map( A1 => Set_target(24), A2 => n491, B1 => n492, B2 
                           => pc_target_18_24_port, ZN => n495);
   U681 : INV_X1 port map( A => n496, ZN => n5910);
   U682 : AOI22_X1 port map( A1 => Set_target(22), A2 => n491, B1 => n492, B2 
                           => pc_target_18_22_port, ZN => n496);
   U683 : INV_X1 port map( A => n497, ZN => n5911);
   U684 : AOI22_X1 port map( A1 => Set_target(20), A2 => n491, B1 => n492, B2 
                           => pc_target_18_20_port, ZN => n497);
   U685 : INV_X1 port map( A => n498, ZN => n5912);
   U686 : AOI22_X1 port map( A1 => Set_target(18), A2 => n491, B1 => n492, B2 
                           => pc_target_18_18_port, ZN => n498);
   U687 : INV_X1 port map( A => n499, ZN => n5913);
   U688 : AOI22_X1 port map( A1 => Set_target(16), A2 => n491, B1 => n492, B2 
                           => pc_target_18_16_port, ZN => n499);
   U689 : INV_X1 port map( A => n500, ZN => n5914);
   U690 : AOI22_X1 port map( A1 => Set_target(14), A2 => n491, B1 => n492, B2 
                           => pc_target_18_14_port, ZN => n500);
   U691 : INV_X1 port map( A => n501, ZN => n5915);
   U692 : AOI22_X1 port map( A1 => Set_target(12), A2 => n491, B1 => n492, B2 
                           => pc_target_18_12_port, ZN => n501);
   U693 : INV_X1 port map( A => n502, ZN => n5916);
   U694 : AOI22_X1 port map( A1 => Set_target(10), A2 => n491, B1 => n492, B2 
                           => pc_target_18_10_port, ZN => n502);
   U695 : INV_X1 port map( A => n503, ZN => n5917);
   U696 : AOI22_X1 port map( A1 => Set_target(8), A2 => n491, B1 => n492, B2 =>
                           pc_target_18_8_port, ZN => n503);
   U697 : INV_X1 port map( A => n504, ZN => n5918);
   U698 : AOI22_X1 port map( A1 => Set_target(6), A2 => n491, B1 => n492, B2 =>
                           pc_target_18_6_port, ZN => n504);
   U699 : INV_X1 port map( A => n505, ZN => n5919);
   U700 : AOI22_X1 port map( A1 => Set_target(4), A2 => n491, B1 => n492, B2 =>
                           pc_target_18_4_port, ZN => n505);
   U701 : INV_X1 port map( A => n506, ZN => n5920);
   U702 : AOI22_X1 port map( A1 => Set_target(2), A2 => n491, B1 => n492, B2 =>
                           pc_target_18_2_port, ZN => n506);
   U703 : INV_X1 port map( A => n507, ZN => n5921);
   U704 : AOI22_X1 port map( A1 => Set_target(0), A2 => n491, B1 => n492, B2 =>
                           pc_target_18_0_port, ZN => n507);
   U705 : INV_X1 port map( A => n508, ZN => n5922);
   U706 : AOI22_X1 port map( A1 => Set_target(1), A2 => n491, B1 => n492, B2 =>
                           pc_target_18_1_port, ZN => n508);
   U707 : INV_X1 port map( A => n509, ZN => n5923);
   U708 : AOI22_X1 port map( A1 => Set_target(3), A2 => n491, B1 => n492, B2 =>
                           pc_target_18_3_port, ZN => n509);
   U709 : INV_X1 port map( A => n510, ZN => n5924);
   U710 : AOI22_X1 port map( A1 => Set_target(5), A2 => n491, B1 => n492, B2 =>
                           pc_target_18_5_port, ZN => n510);
   U711 : INV_X1 port map( A => n511, ZN => n5925);
   U712 : AOI22_X1 port map( A1 => Set_target(7), A2 => n491, B1 => n492, B2 =>
                           pc_target_18_7_port, ZN => n511);
   U713 : INV_X1 port map( A => n512, ZN => n5926);
   U714 : AOI22_X1 port map( A1 => Set_target(9), A2 => n491, B1 => n492, B2 =>
                           pc_target_18_9_port, ZN => n512);
   U715 : INV_X1 port map( A => n513, ZN => n5927);
   U716 : AOI22_X1 port map( A1 => Set_target(11), A2 => n491, B1 => n492, B2 
                           => pc_target_18_11_port, ZN => n513);
   U717 : INV_X1 port map( A => n514, ZN => n5928);
   U718 : AOI22_X1 port map( A1 => Set_target(13), A2 => n491, B1 => n492, B2 
                           => pc_target_18_13_port, ZN => n514);
   U719 : INV_X1 port map( A => n515, ZN => n5929);
   U720 : AOI22_X1 port map( A1 => Set_target(15), A2 => n491, B1 => n492, B2 
                           => pc_target_18_15_port, ZN => n515);
   U721 : INV_X1 port map( A => n516, ZN => n5930);
   U722 : AOI22_X1 port map( A1 => Set_target(17), A2 => n491, B1 => n492, B2 
                           => pc_target_18_17_port, ZN => n516);
   U723 : INV_X1 port map( A => n517, ZN => n5931);
   U724 : AOI22_X1 port map( A1 => Set_target(19), A2 => n491, B1 => n492, B2 
                           => pc_target_18_19_port, ZN => n517);
   U725 : INV_X1 port map( A => n518, ZN => n5932);
   U726 : AOI22_X1 port map( A1 => Set_target(21), A2 => n491, B1 => n492, B2 
                           => pc_target_18_21_port, ZN => n518);
   U727 : INV_X1 port map( A => n519, ZN => n5933);
   U728 : AOI22_X1 port map( A1 => Set_target(23), A2 => n491, B1 => n492, B2 
                           => pc_target_18_23_port, ZN => n519);
   U729 : INV_X1 port map( A => n520, ZN => n5934);
   U730 : AOI22_X1 port map( A1 => Set_target(25), A2 => n491, B1 => n492, B2 
                           => pc_target_18_25_port, ZN => n520);
   U731 : INV_X1 port map( A => n521, ZN => n5935);
   U732 : AOI22_X1 port map( A1 => Set_target(27), A2 => n491, B1 => n492, B2 
                           => pc_target_18_27_port, ZN => n521);
   U733 : INV_X1 port map( A => n522, ZN => n5936);
   U734 : AOI22_X1 port map( A1 => Set_target(29), A2 => n491, B1 => n492, B2 
                           => pc_target_18_29_port, ZN => n522);
   U735 : INV_X1 port map( A => n523, ZN => n5937);
   U736 : AOI22_X1 port map( A1 => Set_target(31), A2 => n491, B1 => n492, B2 
                           => pc_target_18_31_port, ZN => n523);
   U739 : OAI22_X1 port map( A1 => n75, A2 => n524, B1 => n3445, B2 => n526, ZN
                           => n5938);
   U740 : OAI22_X1 port map( A1 => n79, A2 => n524, B1 => n3445, B2 => n527, ZN
                           => n5939);
   U741 : OAI22_X1 port map( A1 => n81, A2 => n524, B1 => n3445, B2 => n528, ZN
                           => n5940);
   U742 : OAI22_X1 port map( A1 => n83, A2 => n524, B1 => n3445, B2 => n529, ZN
                           => n5941);
   U743 : OAI22_X1 port map( A1 => n85, A2 => n524, B1 => n3445, B2 => n530, ZN
                           => n5942);
   U744 : OAI22_X1 port map( A1 => n87, A2 => n524, B1 => n3445, B2 => n531, ZN
                           => n5943);
   U745 : OAI22_X1 port map( A1 => n89, A2 => n524, B1 => n3445, B2 => n532, ZN
                           => n5944);
   U746 : OAI22_X1 port map( A1 => n91, A2 => n524, B1 => n3445, B2 => n533, ZN
                           => n5945);
   U747 : OAI22_X1 port map( A1 => n93, A2 => n524, B1 => n3445, B2 => n534, ZN
                           => n5946);
   U748 : OAI22_X1 port map( A1 => n95, A2 => n524, B1 => n3445, B2 => n535, ZN
                           => n5947);
   U749 : OAI22_X1 port map( A1 => n97_port, A2 => n524, B1 => n3445, B2 => 
                           n536, ZN => n5948);
   U750 : OAI22_X1 port map( A1 => n99_port, A2 => n524, B1 => n3445, B2 => 
                           n537, ZN => n5949);
   U751 : OAI22_X1 port map( A1 => n101_port, A2 => n524, B1 => n3445, B2 => 
                           n538, ZN => n5950);
   U752 : OAI22_X1 port map( A1 => n103_port, A2 => n524, B1 => n3445, B2 => 
                           n539, ZN => n5951);
   U753 : OAI22_X1 port map( A1 => n105_port, A2 => n524, B1 => n3445, B2 => 
                           n540, ZN => n5952);
   U754 : OAI22_X1 port map( A1 => n107_port, A2 => n524, B1 => n3445, B2 => 
                           n541, ZN => n5953);
   U755 : OAI22_X1 port map( A1 => n109_port, A2 => n524, B1 => n3445, B2 => 
                           n542, ZN => n5954);
   U756 : OAI22_X1 port map( A1 => n111_port, A2 => n524, B1 => n3445, B2 => 
                           n543, ZN => n5955);
   U757 : OAI22_X1 port map( A1 => n113_port, A2 => n524, B1 => n3445, B2 => 
                           n544, ZN => n5956);
   U758 : OAI22_X1 port map( A1 => n115_port, A2 => n524, B1 => n3445, B2 => 
                           n545, ZN => n5957);
   U759 : OAI22_X1 port map( A1 => n117_port, A2 => n524, B1 => n3445, B2 => 
                           n546, ZN => n5958);
   U760 : OAI22_X1 port map( A1 => n119_port, A2 => n524, B1 => n3445, B2 => 
                           n547, ZN => n5959);
   U761 : OAI22_X1 port map( A1 => n121_port, A2 => n524, B1 => n3445, B2 => 
                           n548, ZN => n5960);
   U762 : OAI22_X1 port map( A1 => n123_port, A2 => n524, B1 => n3445, B2 => 
                           n549, ZN => n5961);
   U763 : OAI22_X1 port map( A1 => n125_port, A2 => n524, B1 => n3445, B2 => 
                           n550, ZN => n5962);
   U764 : OAI22_X1 port map( A1 => n127_port, A2 => n524, B1 => n3445, B2 => 
                           n551, ZN => n5963);
   U765 : OAI22_X1 port map( A1 => n129, A2 => n524, B1 => n3445, B2 => n552, 
                           ZN => n5964);
   U766 : OAI22_X1 port map( A1 => n131, A2 => n524, B1 => n3445, B2 => n553, 
                           ZN => n5965);
   U767 : OAI22_X1 port map( A1 => n133, A2 => n524, B1 => n3445, B2 => n554, 
                           ZN => n5966);
   U768 : OAI22_X1 port map( A1 => n135, A2 => n524, B1 => n3445, B2 => n555, 
                           ZN => n5967);
   U769 : OAI22_X1 port map( A1 => n137, A2 => n524, B1 => n3445, B2 => n556, 
                           ZN => n5968);
   U770 : OAI22_X1 port map( A1 => n139, A2 => n524, B1 => n3445, B2 => n557, 
                           ZN => n5969);
   U773 : OAI22_X1 port map( A1 => n75, A2 => n1463, B1 => n559, B2 => n560, ZN
                           => n5970);
   U774 : OAI22_X1 port map( A1 => n79, A2 => n1481, B1 => n559, B2 => n561, ZN
                           => n5971);
   U775 : OAI22_X1 port map( A1 => n81, A2 => n1481, B1 => n559, B2 => n562, ZN
                           => n5972);
   U776 : OAI22_X1 port map( A1 => n83, A2 => n1481, B1 => n559, B2 => n563, ZN
                           => n5973);
   U778 : OAI22_X1 port map( A1 => n87, A2 => n1463, B1 => n559, B2 => n565, ZN
                           => n5975);
   U779 : OAI22_X1 port map( A1 => n89, A2 => n1481, B1 => n559, B2 => n566, ZN
                           => n5976);
   U780 : OAI22_X1 port map( A1 => n91, A2 => n1463, B1 => n559, B2 => n567, ZN
                           => n5977);
   U781 : OAI22_X1 port map( A1 => n93, A2 => n1481, B1 => n559, B2 => n568, ZN
                           => n5978);
   U782 : OAI22_X1 port map( A1 => n95, A2 => n1463, B1 => n559, B2 => n569, ZN
                           => n5979);
   U783 : OAI22_X1 port map( A1 => n97_port, A2 => n1481, B1 => n559, B2 => 
                           n570, ZN => n5980);
   U784 : OAI22_X1 port map( A1 => n99_port, A2 => n1481, B1 => n559, B2 => 
                           n571, ZN => n5981);
   U785 : OAI22_X1 port map( A1 => n101_port, A2 => n1481, B1 => n559, B2 => 
                           n572, ZN => n5982);
   U786 : OAI22_X1 port map( A1 => n103_port, A2 => n1481, B1 => n559, B2 => 
                           n573, ZN => n5983);
   U787 : OAI22_X1 port map( A1 => n105_port, A2 => n1481, B1 => n559, B2 => 
                           n574, ZN => n5984);
   U788 : OAI22_X1 port map( A1 => n107_port, A2 => n1481, B1 => n559, B2 => 
                           n575, ZN => n5985);
   U789 : OAI22_X1 port map( A1 => n109_port, A2 => n1481, B1 => n559, B2 => 
                           n576, ZN => n5986);
   U790 : OAI22_X1 port map( A1 => n111_port, A2 => n1481, B1 => n559, B2 => 
                           n577, ZN => n5987);
   U791 : OAI22_X1 port map( A1 => n113_port, A2 => n1481, B1 => n559, B2 => 
                           n578, ZN => n5988);
   U792 : OAI22_X1 port map( A1 => n115_port, A2 => n1481, B1 => n559, B2 => 
                           n579, ZN => n5989);
   U793 : OAI22_X1 port map( A1 => n117_port, A2 => n1481, B1 => n559, B2 => 
                           n580, ZN => n5990);
   U794 : OAI22_X1 port map( A1 => n119_port, A2 => n1481, B1 => n559, B2 => 
                           n581, ZN => n5991);
   U795 : OAI22_X1 port map( A1 => n121_port, A2 => n1481, B1 => n559, B2 => 
                           n582, ZN => n5992);
   U796 : OAI22_X1 port map( A1 => n123_port, A2 => n1481, B1 => n559, B2 => 
                           n583, ZN => n5993);
   U797 : OAI22_X1 port map( A1 => n125_port, A2 => n1481, B1 => n559, B2 => 
                           n584, ZN => n5994);
   U798 : OAI22_X1 port map( A1 => n127_port, A2 => n1481, B1 => n559, B2 => 
                           n585, ZN => n5995);
   U799 : OAI22_X1 port map( A1 => n129, A2 => n1481, B1 => n559, B2 => n586, 
                           ZN => n5996);
   U800 : OAI22_X1 port map( A1 => n131, A2 => n1481, B1 => n559, B2 => n587, 
                           ZN => n5997);
   U801 : OAI22_X1 port map( A1 => n133, A2 => n1481, B1 => n559, B2 => n588, 
                           ZN => n5998);
   U802 : OAI22_X1 port map( A1 => n135, A2 => n1463, B1 => n559, B2 => n589, 
                           ZN => n5999);
   U803 : OAI22_X1 port map( A1 => n137, A2 => n1481, B1 => n559, B2 => n590, 
                           ZN => n6000);
   U804 : OAI22_X1 port map( A1 => n139, A2 => n1481, B1 => n559, B2 => n591, 
                           ZN => n6001);
   U809 : INV_X1 port map( A => n594, ZN => n6002);
   U810 : AOI22_X1 port map( A1 => Set_target(30), A2 => n595, B1 => n596, B2 
                           => pc_target_15_30_port, ZN => n594);
   U811 : INV_X1 port map( A => n597, ZN => n6003);
   U812 : AOI22_X1 port map( A1 => Set_target(28), A2 => n595, B1 => n596, B2 
                           => pc_target_15_28_port, ZN => n597);
   U813 : INV_X1 port map( A => n598, ZN => n6004);
   U814 : AOI22_X1 port map( A1 => Set_target(26), A2 => n595, B1 => n596, B2 
                           => pc_target_15_26_port, ZN => n598);
   U815 : INV_X1 port map( A => n599, ZN => n6005);
   U816 : AOI22_X1 port map( A1 => Set_target(24), A2 => n595, B1 => n596, B2 
                           => pc_target_15_24_port, ZN => n599);
   U817 : INV_X1 port map( A => n600, ZN => n6006);
   U818 : AOI22_X1 port map( A1 => Set_target(22), A2 => n595, B1 => n596, B2 
                           => pc_target_15_22_port, ZN => n600);
   U819 : INV_X1 port map( A => n601, ZN => n6007);
   U820 : AOI22_X1 port map( A1 => Set_target(20), A2 => n595, B1 => n596, B2 
                           => pc_target_15_20_port, ZN => n601);
   U821 : INV_X1 port map( A => n602, ZN => n6008);
   U822 : AOI22_X1 port map( A1 => Set_target(18), A2 => n595, B1 => n596, B2 
                           => pc_target_15_18_port, ZN => n602);
   U823 : INV_X1 port map( A => n603, ZN => n6009);
   U824 : AOI22_X1 port map( A1 => Set_target(16), A2 => n595, B1 => n596, B2 
                           => pc_target_15_16_port, ZN => n603);
   U825 : INV_X1 port map( A => n604, ZN => n6010);
   U826 : AOI22_X1 port map( A1 => Set_target(14), A2 => n595, B1 => n596, B2 
                           => pc_target_15_14_port, ZN => n604);
   U827 : INV_X1 port map( A => n605, ZN => n6011);
   U828 : AOI22_X1 port map( A1 => Set_target(12), A2 => n595, B1 => n596, B2 
                           => pc_target_15_12_port, ZN => n605);
   U829 : INV_X1 port map( A => n606, ZN => n6012);
   U830 : AOI22_X1 port map( A1 => Set_target(10), A2 => n595, B1 => n596, B2 
                           => pc_target_15_10_port, ZN => n606);
   U831 : INV_X1 port map( A => n607, ZN => n6013);
   U832 : AOI22_X1 port map( A1 => Set_target(8), A2 => n595, B1 => n596, B2 =>
                           pc_target_15_8_port, ZN => n607);
   U833 : INV_X1 port map( A => n608, ZN => n6014);
   U834 : AOI22_X1 port map( A1 => Set_target(6), A2 => n595, B1 => n596, B2 =>
                           pc_target_15_6_port, ZN => n608);
   U835 : INV_X1 port map( A => n609, ZN => n6015);
   U836 : AOI22_X1 port map( A1 => Set_target(4), A2 => n595, B1 => n596, B2 =>
                           pc_target_15_4_port, ZN => n609);
   U837 : INV_X1 port map( A => n610, ZN => n6016);
   U838 : AOI22_X1 port map( A1 => Set_target(2), A2 => n595, B1 => n596, B2 =>
                           pc_target_15_2_port, ZN => n610);
   U839 : INV_X1 port map( A => n611, ZN => n6017);
   U840 : AOI22_X1 port map( A1 => Set_target(0), A2 => n595, B1 => n596, B2 =>
                           pc_target_15_0_port, ZN => n611);
   U841 : INV_X1 port map( A => n612, ZN => n6018);
   U842 : AOI22_X1 port map( A1 => Set_target(1), A2 => n595, B1 => n596, B2 =>
                           pc_target_15_1_port, ZN => n612);
   U843 : INV_X1 port map( A => n613, ZN => n6019);
   U844 : AOI22_X1 port map( A1 => Set_target(3), A2 => n595, B1 => n596, B2 =>
                           pc_target_15_3_port, ZN => n613);
   U845 : INV_X1 port map( A => n614, ZN => n6020);
   U846 : AOI22_X1 port map( A1 => Set_target(5), A2 => n595, B1 => n596, B2 =>
                           pc_target_15_5_port, ZN => n614);
   U847 : INV_X1 port map( A => n615, ZN => n6021);
   U848 : AOI22_X1 port map( A1 => Set_target(7), A2 => n595, B1 => n596, B2 =>
                           pc_target_15_7_port, ZN => n615);
   U849 : INV_X1 port map( A => n616, ZN => n6022);
   U850 : AOI22_X1 port map( A1 => Set_target(9), A2 => n595, B1 => n596, B2 =>
                           pc_target_15_9_port, ZN => n616);
   U851 : INV_X1 port map( A => n617, ZN => n6023);
   U852 : AOI22_X1 port map( A1 => Set_target(11), A2 => n595, B1 => n596, B2 
                           => pc_target_15_11_port, ZN => n617);
   U853 : INV_X1 port map( A => n618, ZN => n6024);
   U854 : AOI22_X1 port map( A1 => Set_target(13), A2 => n595, B1 => n596, B2 
                           => pc_target_15_13_port, ZN => n618);
   U855 : INV_X1 port map( A => n619, ZN => n6025);
   U856 : AOI22_X1 port map( A1 => Set_target(15), A2 => n595, B1 => n596, B2 
                           => pc_target_15_15_port, ZN => n619);
   U857 : INV_X1 port map( A => n620, ZN => n6026);
   U858 : AOI22_X1 port map( A1 => Set_target(17), A2 => n595, B1 => n596, B2 
                           => pc_target_15_17_port, ZN => n620);
   U859 : INV_X1 port map( A => n621, ZN => n6027);
   U860 : AOI22_X1 port map( A1 => Set_target(19), A2 => n595, B1 => n596, B2 
                           => pc_target_15_19_port, ZN => n621);
   U861 : INV_X1 port map( A => n622, ZN => n6028);
   U862 : AOI22_X1 port map( A1 => Set_target(21), A2 => n595, B1 => n596, B2 
                           => pc_target_15_21_port, ZN => n622);
   U863 : INV_X1 port map( A => n623, ZN => n6029);
   U864 : AOI22_X1 port map( A1 => Set_target(23), A2 => n595, B1 => n596, B2 
                           => pc_target_15_23_port, ZN => n623);
   U865 : INV_X1 port map( A => n624, ZN => n6030);
   U866 : AOI22_X1 port map( A1 => Set_target(25), A2 => n595, B1 => n596, B2 
                           => pc_target_15_25_port, ZN => n624);
   U867 : INV_X1 port map( A => n625, ZN => n6031);
   U868 : AOI22_X1 port map( A1 => Set_target(27), A2 => n595, B1 => n596, B2 
                           => pc_target_15_27_port, ZN => n625);
   U869 : INV_X1 port map( A => n626, ZN => n6032);
   U870 : AOI22_X1 port map( A1 => Set_target(29), A2 => n595, B1 => n596, B2 
                           => pc_target_15_29_port, ZN => n626);
   U871 : INV_X1 port map( A => n627, ZN => n6033);
   U872 : AOI22_X1 port map( A1 => Set_target(31), A2 => n595, B1 => n596, B2 
                           => pc_target_15_31_port, ZN => n627);
   U875 : INV_X1 port map( A => n629, ZN => n6034);
   U876 : AOI22_X1 port map( A1 => Set_target(30), A2 => n630, B1 => n631, B2 
                           => pc_target_14_30_port, ZN => n629);
   U877 : INV_X1 port map( A => n632, ZN => n6035);
   U878 : AOI22_X1 port map( A1 => Set_target(28), A2 => n630, B1 => n631, B2 
                           => pc_target_14_28_port, ZN => n632);
   U879 : INV_X1 port map( A => n633, ZN => n6036);
   U880 : AOI22_X1 port map( A1 => Set_target(26), A2 => n630, B1 => n631, B2 
                           => pc_target_14_26_port, ZN => n633);
   U881 : INV_X1 port map( A => n634, ZN => n6037);
   U882 : AOI22_X1 port map( A1 => Set_target(24), A2 => n630, B1 => n631, B2 
                           => pc_target_14_24_port, ZN => n634);
   U883 : INV_X1 port map( A => n635, ZN => n6038);
   U884 : AOI22_X1 port map( A1 => Set_target(22), A2 => n630, B1 => n631, B2 
                           => pc_target_14_22_port, ZN => n635);
   U885 : INV_X1 port map( A => n636, ZN => n6039);
   U886 : AOI22_X1 port map( A1 => Set_target(20), A2 => n630, B1 => n631, B2 
                           => pc_target_14_20_port, ZN => n636);
   U887 : INV_X1 port map( A => n637, ZN => n6040);
   U888 : AOI22_X1 port map( A1 => Set_target(18), A2 => n630, B1 => n631, B2 
                           => pc_target_14_18_port, ZN => n637);
   U889 : INV_X1 port map( A => n638, ZN => n6041);
   U890 : AOI22_X1 port map( A1 => Set_target(16), A2 => n630, B1 => n631, B2 
                           => pc_target_14_16_port, ZN => n638);
   U891 : INV_X1 port map( A => n639, ZN => n6042);
   U892 : AOI22_X1 port map( A1 => Set_target(14), A2 => n630, B1 => n631, B2 
                           => pc_target_14_14_port, ZN => n639);
   U893 : INV_X1 port map( A => n640, ZN => n6043);
   U894 : AOI22_X1 port map( A1 => Set_target(12), A2 => n630, B1 => n631, B2 
                           => pc_target_14_12_port, ZN => n640);
   U895 : INV_X1 port map( A => n641, ZN => n6044);
   U896 : AOI22_X1 port map( A1 => Set_target(10), A2 => n630, B1 => n631, B2 
                           => pc_target_14_10_port, ZN => n641);
   U897 : INV_X1 port map( A => n642, ZN => n6045);
   U898 : AOI22_X1 port map( A1 => Set_target(8), A2 => n630, B1 => n631, B2 =>
                           pc_target_14_8_port, ZN => n642);
   U899 : INV_X1 port map( A => n643, ZN => n6046);
   U900 : AOI22_X1 port map( A1 => Set_target(6), A2 => n630, B1 => n631, B2 =>
                           pc_target_14_6_port, ZN => n643);
   U901 : INV_X1 port map( A => n644, ZN => n6047);
   U902 : AOI22_X1 port map( A1 => Set_target(4), A2 => n630, B1 => n631, B2 =>
                           pc_target_14_4_port, ZN => n644);
   U903 : INV_X1 port map( A => n645, ZN => n6048);
   U904 : AOI22_X1 port map( A1 => Set_target(2), A2 => n630, B1 => n631, B2 =>
                           pc_target_14_2_port, ZN => n645);
   U905 : INV_X1 port map( A => n646, ZN => n6049);
   U906 : AOI22_X1 port map( A1 => Set_target(0), A2 => n630, B1 => n631, B2 =>
                           pc_target_14_0_port, ZN => n646);
   U907 : INV_X1 port map( A => n647, ZN => n6050);
   U908 : AOI22_X1 port map( A1 => Set_target(1), A2 => n630, B1 => n631, B2 =>
                           pc_target_14_1_port, ZN => n647);
   U909 : INV_X1 port map( A => n648, ZN => n6051);
   U910 : AOI22_X1 port map( A1 => Set_target(3), A2 => n630, B1 => n631, B2 =>
                           pc_target_14_3_port, ZN => n648);
   U911 : INV_X1 port map( A => n649, ZN => n6052);
   U912 : AOI22_X1 port map( A1 => Set_target(5), A2 => n630, B1 => n631, B2 =>
                           pc_target_14_5_port, ZN => n649);
   U913 : INV_X1 port map( A => n650, ZN => n6053);
   U914 : AOI22_X1 port map( A1 => Set_target(7), A2 => n630, B1 => n631, B2 =>
                           pc_target_14_7_port, ZN => n650);
   U915 : INV_X1 port map( A => n651, ZN => n6054);
   U916 : AOI22_X1 port map( A1 => Set_target(9), A2 => n630, B1 => n631, B2 =>
                           pc_target_14_9_port, ZN => n651);
   U917 : INV_X1 port map( A => n652, ZN => n6055);
   U918 : AOI22_X1 port map( A1 => Set_target(11), A2 => n630, B1 => n631, B2 
                           => pc_target_14_11_port, ZN => n652);
   U919 : INV_X1 port map( A => n653, ZN => n6056);
   U920 : AOI22_X1 port map( A1 => Set_target(13), A2 => n630, B1 => n631, B2 
                           => pc_target_14_13_port, ZN => n653);
   U921 : INV_X1 port map( A => n654, ZN => n6057);
   U922 : AOI22_X1 port map( A1 => Set_target(15), A2 => n630, B1 => n631, B2 
                           => pc_target_14_15_port, ZN => n654);
   U923 : INV_X1 port map( A => n655, ZN => n6058);
   U924 : AOI22_X1 port map( A1 => Set_target(17), A2 => n630, B1 => n631, B2 
                           => pc_target_14_17_port, ZN => n655);
   U925 : INV_X1 port map( A => n656, ZN => n6059);
   U926 : AOI22_X1 port map( A1 => Set_target(19), A2 => n630, B1 => n631, B2 
                           => pc_target_14_19_port, ZN => n656);
   U927 : INV_X1 port map( A => n657, ZN => n6060);
   U928 : AOI22_X1 port map( A1 => Set_target(21), A2 => n630, B1 => n631, B2 
                           => pc_target_14_21_port, ZN => n657);
   U929 : INV_X1 port map( A => n658, ZN => n6061);
   U930 : AOI22_X1 port map( A1 => Set_target(23), A2 => n630, B1 => n631, B2 
                           => pc_target_14_23_port, ZN => n658);
   U931 : INV_X1 port map( A => n659, ZN => n6062);
   U932 : AOI22_X1 port map( A1 => Set_target(25), A2 => n630, B1 => n631, B2 
                           => pc_target_14_25_port, ZN => n659);
   U933 : INV_X1 port map( A => n660, ZN => n6063);
   U934 : AOI22_X1 port map( A1 => Set_target(27), A2 => n630, B1 => n631, B2 
                           => pc_target_14_27_port, ZN => n660);
   U935 : INV_X1 port map( A => n661, ZN => n6064);
   U936 : AOI22_X1 port map( A1 => Set_target(29), A2 => n630, B1 => n631, B2 
                           => pc_target_14_29_port, ZN => n661);
   U937 : INV_X1 port map( A => n662, ZN => n6065);
   U938 : AOI22_X1 port map( A1 => Set_target(31), A2 => n630, B1 => n631, B2 
                           => pc_target_14_31_port, ZN => n662);
   U941 : OAI22_X1 port map( A1 => n75, A2 => n663, B1 => n664, B2 => n665, ZN 
                           => n6066);
   U942 : OAI22_X1 port map( A1 => n79, A2 => n663, B1 => n664, B2 => n666, ZN 
                           => n6067);
   U943 : OAI22_X1 port map( A1 => n81, A2 => n663, B1 => n664, B2 => n667, ZN 
                           => n6068);
   U944 : OAI22_X1 port map( A1 => n83, A2 => n663, B1 => n664, B2 => n668, ZN 
                           => n6069);
   U945 : OAI22_X1 port map( A1 => n85, A2 => n663, B1 => n664, B2 => n669, ZN 
                           => n6070);
   U946 : OAI22_X1 port map( A1 => n87, A2 => n663, B1 => n664, B2 => n670, ZN 
                           => n6071);
   U947 : OAI22_X1 port map( A1 => n89, A2 => n663, B1 => n664, B2 => n671, ZN 
                           => n6072);
   U948 : OAI22_X1 port map( A1 => n91, A2 => n663, B1 => n664, B2 => n672, ZN 
                           => n6073);
   U949 : OAI22_X1 port map( A1 => n93, A2 => n663, B1 => n664, B2 => n673, ZN 
                           => n6074);
   U950 : OAI22_X1 port map( A1 => n95, A2 => n663, B1 => n664, B2 => n674, ZN 
                           => n6075);
   U951 : OAI22_X1 port map( A1 => n97_port, A2 => n663, B1 => n664, B2 => n675
                           , ZN => n6076);
   U952 : OAI22_X1 port map( A1 => n99_port, A2 => n663, B1 => n664, B2 => n676
                           , ZN => n6077);
   U953 : OAI22_X1 port map( A1 => n101_port, A2 => n663, B1 => n664, B2 => 
                           n677, ZN => n6078);
   U954 : OAI22_X1 port map( A1 => n103_port, A2 => n663, B1 => n664, B2 => 
                           n678, ZN => n6079);
   U955 : OAI22_X1 port map( A1 => n105_port, A2 => n663, B1 => n664, B2 => 
                           n679, ZN => n6080);
   U956 : OAI22_X1 port map( A1 => n107_port, A2 => n663, B1 => n664, B2 => 
                           n680, ZN => n6081);
   U957 : OAI22_X1 port map( A1 => n109_port, A2 => n663, B1 => n664, B2 => 
                           n681, ZN => n6082);
   U958 : OAI22_X1 port map( A1 => n111_port, A2 => n663, B1 => n664, B2 => 
                           n682, ZN => n6083);
   U959 : OAI22_X1 port map( A1 => n113_port, A2 => n663, B1 => n664, B2 => 
                           n683, ZN => n6084);
   U960 : OAI22_X1 port map( A1 => n115_port, A2 => n663, B1 => n664, B2 => 
                           n684, ZN => n6085);
   U961 : OAI22_X1 port map( A1 => n117_port, A2 => n663, B1 => n664, B2 => 
                           n685, ZN => n6086);
   U962 : OAI22_X1 port map( A1 => n119_port, A2 => n663, B1 => n664, B2 => 
                           n686, ZN => n6087);
   U963 : OAI22_X1 port map( A1 => n121_port, A2 => n663, B1 => n664, B2 => 
                           n687, ZN => n6088);
   U964 : OAI22_X1 port map( A1 => n123_port, A2 => n663, B1 => n664, B2 => 
                           n688, ZN => n6089);
   U965 : OAI22_X1 port map( A1 => n125_port, A2 => n663, B1 => n664, B2 => 
                           n689, ZN => n6090);
   U966 : OAI22_X1 port map( A1 => n127_port, A2 => n663, B1 => n664, B2 => 
                           n690, ZN => n6091);
   U967 : OAI22_X1 port map( A1 => n129, A2 => n663, B1 => n664, B2 => n691, ZN
                           => n6092);
   U968 : OAI22_X1 port map( A1 => n131, A2 => n663, B1 => n664, B2 => n692, ZN
                           => n6093);
   U969 : OAI22_X1 port map( A1 => n133, A2 => n663, B1 => n664, B2 => n693, ZN
                           => n6094);
   U970 : OAI22_X1 port map( A1 => n135, A2 => n663, B1 => n664, B2 => n694, ZN
                           => n6095);
   U971 : OAI22_X1 port map( A1 => n137, A2 => n663, B1 => n664, B2 => n695, ZN
                           => n6096);
   U972 : OAI22_X1 port map( A1 => n139, A2 => n663, B1 => n664, B2 => n696, ZN
                           => n6097);
   U975 : OAI22_X1 port map( A1 => n75, A2 => n697, B1 => n698, B2 => n699, ZN 
                           => n6098);
   U976 : OAI22_X1 port map( A1 => n79, A2 => n697, B1 => n698, B2 => n700, ZN 
                           => n6099);
   U977 : OAI22_X1 port map( A1 => n81, A2 => n697, B1 => n698, B2 => n701, ZN 
                           => n6100);
   U978 : OAI22_X1 port map( A1 => n83, A2 => n697, B1 => n698, B2 => n702, ZN 
                           => n6101);
   U979 : OAI22_X1 port map( A1 => n85, A2 => n697, B1 => n698, B2 => n703, ZN 
                           => n6102);
   U980 : OAI22_X1 port map( A1 => n87, A2 => n697, B1 => n698, B2 => n704, ZN 
                           => n6103);
   U981 : OAI22_X1 port map( A1 => n89, A2 => n697, B1 => n698, B2 => n705, ZN 
                           => n6104);
   U982 : OAI22_X1 port map( A1 => n91, A2 => n697, B1 => n698, B2 => n706, ZN 
                           => n6105);
   U983 : OAI22_X1 port map( A1 => n93, A2 => n697, B1 => n698, B2 => n707, ZN 
                           => n6106);
   U984 : OAI22_X1 port map( A1 => n95, A2 => n697, B1 => n698, B2 => n708, ZN 
                           => n6107);
   U985 : OAI22_X1 port map( A1 => n97_port, A2 => n697, B1 => n698, B2 => n709
                           , ZN => n6108);
   U986 : OAI22_X1 port map( A1 => n99_port, A2 => n697, B1 => n698, B2 => n710
                           , ZN => n6109);
   U987 : OAI22_X1 port map( A1 => n101_port, A2 => n697, B1 => n698, B2 => 
                           n711, ZN => n6110);
   U988 : OAI22_X1 port map( A1 => n103_port, A2 => n697, B1 => n698, B2 => 
                           n712, ZN => n6111);
   U989 : OAI22_X1 port map( A1 => n105_port, A2 => n697, B1 => n698, B2 => 
                           n713, ZN => n6112);
   U990 : OAI22_X1 port map( A1 => n107_port, A2 => n697, B1 => n698, B2 => 
                           n714, ZN => n6113);
   U991 : OAI22_X1 port map( A1 => n109_port, A2 => n697, B1 => n698, B2 => 
                           n715, ZN => n6114);
   U992 : OAI22_X1 port map( A1 => n111_port, A2 => n697, B1 => n698, B2 => 
                           n716, ZN => n6115);
   U993 : OAI22_X1 port map( A1 => n113_port, A2 => n697, B1 => n698, B2 => 
                           n717, ZN => n6116);
   U994 : OAI22_X1 port map( A1 => n115_port, A2 => n697, B1 => n698, B2 => 
                           n718, ZN => n6117);
   U995 : OAI22_X1 port map( A1 => n117_port, A2 => n697, B1 => n698, B2 => 
                           n719, ZN => n6118);
   U996 : OAI22_X1 port map( A1 => n119_port, A2 => n697, B1 => n698, B2 => 
                           n720, ZN => n6119);
   U997 : OAI22_X1 port map( A1 => n121_port, A2 => n697, B1 => n698, B2 => 
                           n721, ZN => n6120);
   U998 : OAI22_X1 port map( A1 => n123_port, A2 => n697, B1 => n698, B2 => 
                           n722, ZN => n6121);
   U999 : OAI22_X1 port map( A1 => n125_port, A2 => n697, B1 => n698, B2 => 
                           n723, ZN => n6122);
   U1000 : OAI22_X1 port map( A1 => n127_port, A2 => n697, B1 => n698, B2 => 
                           n724, ZN => n6123);
   U1001 : OAI22_X1 port map( A1 => n129, A2 => n697, B1 => n698, B2 => n725, 
                           ZN => n6124);
   U1002 : OAI22_X1 port map( A1 => n131, A2 => n697, B1 => n698, B2 => n726, 
                           ZN => n6125);
   U1003 : OAI22_X1 port map( A1 => n133, A2 => n697, B1 => n698, B2 => n727, 
                           ZN => n6126);
   U1004 : OAI22_X1 port map( A1 => n135, A2 => n697, B1 => n698, B2 => n728, 
                           ZN => n6127);
   U1005 : OAI22_X1 port map( A1 => n137, A2 => n697, B1 => n698, B2 => n729, 
                           ZN => n6128);
   U1006 : OAI22_X1 port map( A1 => n139, A2 => n697, B1 => n698, B2 => n730, 
                           ZN => n6129);
   U1010 : INV_X1 port map( A => n732, ZN => n6130);
   U1011 : AOI22_X1 port map( A1 => Set_target(30), A2 => n733, B1 => n734, B2 
                           => pc_target_11_30_port, ZN => n732);
   U1012 : INV_X1 port map( A => n735, ZN => n6131);
   U1013 : AOI22_X1 port map( A1 => Set_target(28), A2 => n733, B1 => n734, B2 
                           => pc_target_11_28_port, ZN => n735);
   U1014 : INV_X1 port map( A => n736, ZN => n6132);
   U1015 : AOI22_X1 port map( A1 => Set_target(26), A2 => n733, B1 => n734, B2 
                           => pc_target_11_26_port, ZN => n736);
   U1016 : INV_X1 port map( A => n737, ZN => n6133);
   U1017 : AOI22_X1 port map( A1 => Set_target(24), A2 => n733, B1 => n734, B2 
                           => pc_target_11_24_port, ZN => n737);
   U1018 : INV_X1 port map( A => n738, ZN => n6134);
   U1019 : AOI22_X1 port map( A1 => Set_target(22), A2 => n733, B1 => n734, B2 
                           => pc_target_11_22_port, ZN => n738);
   U1020 : INV_X1 port map( A => n739, ZN => n6135);
   U1021 : AOI22_X1 port map( A1 => Set_target(20), A2 => n733, B1 => n734, B2 
                           => pc_target_11_20_port, ZN => n739);
   U1022 : INV_X1 port map( A => n740, ZN => n6136);
   U1023 : AOI22_X1 port map( A1 => Set_target(18), A2 => n733, B1 => n734, B2 
                           => pc_target_11_18_port, ZN => n740);
   U1024 : INV_X1 port map( A => n741, ZN => n6137);
   U1025 : AOI22_X1 port map( A1 => Set_target(16), A2 => n733, B1 => n734, B2 
                           => pc_target_11_16_port, ZN => n741);
   U1026 : INV_X1 port map( A => n742, ZN => n6138);
   U1027 : AOI22_X1 port map( A1 => Set_target(14), A2 => n733, B1 => n734, B2 
                           => pc_target_11_14_port, ZN => n742);
   U1028 : INV_X1 port map( A => n743, ZN => n6139);
   U1029 : AOI22_X1 port map( A1 => Set_target(12), A2 => n733, B1 => n734, B2 
                           => pc_target_11_12_port, ZN => n743);
   U1030 : INV_X1 port map( A => n744, ZN => n6140);
   U1031 : AOI22_X1 port map( A1 => Set_target(10), A2 => n733, B1 => n734, B2 
                           => pc_target_11_10_port, ZN => n744);
   U1032 : INV_X1 port map( A => n745, ZN => n6141);
   U1033 : AOI22_X1 port map( A1 => Set_target(8), A2 => n733, B1 => n734, B2 
                           => pc_target_11_8_port, ZN => n745);
   U1034 : INV_X1 port map( A => n746, ZN => n6142);
   U1035 : AOI22_X1 port map( A1 => Set_target(6), A2 => n733, B1 => n734, B2 
                           => pc_target_11_6_port, ZN => n746);
   U1036 : INV_X1 port map( A => n747, ZN => n6143);
   U1037 : AOI22_X1 port map( A1 => Set_target(4), A2 => n733, B1 => n734, B2 
                           => pc_target_11_4_port, ZN => n747);
   U1038 : INV_X1 port map( A => n748, ZN => n6144);
   U1039 : AOI22_X1 port map( A1 => Set_target(2), A2 => n733, B1 => n734, B2 
                           => pc_target_11_2_port, ZN => n748);
   U1040 : INV_X1 port map( A => n749, ZN => n6145);
   U1041 : AOI22_X1 port map( A1 => Set_target(0), A2 => n733, B1 => n734, B2 
                           => pc_target_11_0_port, ZN => n749);
   U1042 : INV_X1 port map( A => n750, ZN => n6146);
   U1043 : AOI22_X1 port map( A1 => Set_target(1), A2 => n733, B1 => n734, B2 
                           => pc_target_11_1_port, ZN => n750);
   U1044 : INV_X1 port map( A => n751, ZN => n6147);
   U1045 : AOI22_X1 port map( A1 => Set_target(3), A2 => n733, B1 => n734, B2 
                           => pc_target_11_3_port, ZN => n751);
   U1046 : INV_X1 port map( A => n752, ZN => n6148);
   U1047 : AOI22_X1 port map( A1 => Set_target(5), A2 => n733, B1 => n734, B2 
                           => pc_target_11_5_port, ZN => n752);
   U1048 : INV_X1 port map( A => n753, ZN => n6149);
   U1049 : AOI22_X1 port map( A1 => Set_target(7), A2 => n733, B1 => n734, B2 
                           => pc_target_11_7_port, ZN => n753);
   U1050 : INV_X1 port map( A => n754, ZN => n6150);
   U1051 : AOI22_X1 port map( A1 => Set_target(9), A2 => n733, B1 => n734, B2 
                           => pc_target_11_9_port, ZN => n754);
   U1052 : INV_X1 port map( A => n755, ZN => n6151);
   U1053 : AOI22_X1 port map( A1 => Set_target(11), A2 => n733, B1 => n734, B2 
                           => pc_target_11_11_port, ZN => n755);
   U1054 : INV_X1 port map( A => n756, ZN => n6152);
   U1055 : AOI22_X1 port map( A1 => Set_target(13), A2 => n733, B1 => n734, B2 
                           => pc_target_11_13_port, ZN => n756);
   U1056 : INV_X1 port map( A => n757, ZN => n6153);
   U1057 : AOI22_X1 port map( A1 => Set_target(15), A2 => n733, B1 => n734, B2 
                           => pc_target_11_15_port, ZN => n757);
   U1058 : INV_X1 port map( A => n758, ZN => n6154);
   U1059 : AOI22_X1 port map( A1 => Set_target(17), A2 => n733, B1 => n734, B2 
                           => pc_target_11_17_port, ZN => n758);
   U1060 : INV_X1 port map( A => n759, ZN => n6155);
   U1061 : AOI22_X1 port map( A1 => Set_target(19), A2 => n733, B1 => n734, B2 
                           => pc_target_11_19_port, ZN => n759);
   U1062 : INV_X1 port map( A => n760, ZN => n6156);
   U1063 : AOI22_X1 port map( A1 => Set_target(21), A2 => n733, B1 => n734, B2 
                           => pc_target_11_21_port, ZN => n760);
   U1064 : INV_X1 port map( A => n761, ZN => n6157);
   U1065 : AOI22_X1 port map( A1 => Set_target(23), A2 => n733, B1 => n734, B2 
                           => pc_target_11_23_port, ZN => n761);
   U1066 : INV_X1 port map( A => n762, ZN => n6158);
   U1067 : AOI22_X1 port map( A1 => Set_target(25), A2 => n733, B1 => n734, B2 
                           => pc_target_11_25_port, ZN => n762);
   U1068 : INV_X1 port map( A => n763, ZN => n6159);
   U1069 : AOI22_X1 port map( A1 => Set_target(27), A2 => n733, B1 => n734, B2 
                           => pc_target_11_27_port, ZN => n763);
   U1070 : INV_X1 port map( A => n764, ZN => n6160);
   U1071 : AOI22_X1 port map( A1 => Set_target(29), A2 => n733, B1 => n734, B2 
                           => pc_target_11_29_port, ZN => n764);
   U1072 : INV_X1 port map( A => n765, ZN => n6161);
   U1073 : AOI22_X1 port map( A1 => Set_target(31), A2 => n733, B1 => n734, B2 
                           => pc_target_11_31_port, ZN => n765);
   U1076 : INV_X1 port map( A => n767, ZN => n6162);
   U1077 : AOI22_X1 port map( A1 => Set_target(30), A2 => n3446, B1 => n769, B2
                           => pc_target_10_30_port, ZN => n767);
   U1078 : INV_X1 port map( A => n770, ZN => n6163);
   U1079 : AOI22_X1 port map( A1 => Set_target(28), A2 => n3446, B1 => n769, B2
                           => pc_target_10_28_port, ZN => n770);
   U1080 : INV_X1 port map( A => n771, ZN => n6164);
   U1081 : AOI22_X1 port map( A1 => Set_target(26), A2 => n3446, B1 => n769, B2
                           => pc_target_10_26_port, ZN => n771);
   U1082 : INV_X1 port map( A => n772, ZN => n6165);
   U1083 : AOI22_X1 port map( A1 => Set_target(24), A2 => n3446, B1 => n769, B2
                           => pc_target_10_24_port, ZN => n772);
   U1084 : INV_X1 port map( A => n773, ZN => n6166);
   U1085 : AOI22_X1 port map( A1 => Set_target(22), A2 => n3446, B1 => n769, B2
                           => pc_target_10_22_port, ZN => n773);
   U1086 : INV_X1 port map( A => n774, ZN => n6167);
   U1087 : AOI22_X1 port map( A1 => Set_target(20), A2 => n3446, B1 => n769, B2
                           => pc_target_10_20_port, ZN => n774);
   U1088 : INV_X1 port map( A => n775, ZN => n6168);
   U1089 : AOI22_X1 port map( A1 => Set_target(18), A2 => n3446, B1 => n769, B2
                           => pc_target_10_18_port, ZN => n775);
   U1090 : INV_X1 port map( A => n776, ZN => n6169);
   U1091 : AOI22_X1 port map( A1 => Set_target(16), A2 => n3446, B1 => n769, B2
                           => pc_target_10_16_port, ZN => n776);
   U1092 : INV_X1 port map( A => n777, ZN => n6170);
   U1093 : AOI22_X1 port map( A1 => Set_target(14), A2 => n3446, B1 => n769, B2
                           => pc_target_10_14_port, ZN => n777);
   U1094 : INV_X1 port map( A => n778, ZN => n6171);
   U1095 : AOI22_X1 port map( A1 => Set_target(12), A2 => n3446, B1 => n769, B2
                           => pc_target_10_12_port, ZN => n778);
   U1096 : INV_X1 port map( A => n779, ZN => n6172);
   U1097 : AOI22_X1 port map( A1 => Set_target(10), A2 => n3446, B1 => n769, B2
                           => pc_target_10_10_port, ZN => n779);
   U1098 : INV_X1 port map( A => n780, ZN => n6173);
   U1099 : AOI22_X1 port map( A1 => Set_target(8), A2 => n3446, B1 => n769, B2 
                           => pc_target_10_8_port, ZN => n780);
   U1100 : INV_X1 port map( A => n781, ZN => n6174);
   U1101 : AOI22_X1 port map( A1 => Set_target(6), A2 => n3446, B1 => n769, B2 
                           => pc_target_10_6_port, ZN => n781);
   U1102 : INV_X1 port map( A => n782, ZN => n6175);
   U1103 : AOI22_X1 port map( A1 => Set_target(4), A2 => n3446, B1 => n769, B2 
                           => pc_target_10_4_port, ZN => n782);
   U1104 : INV_X1 port map( A => n783, ZN => n6176);
   U1105 : AOI22_X1 port map( A1 => Set_target(2), A2 => n3446, B1 => n769, B2 
                           => pc_target_10_2_port, ZN => n783);
   U1106 : INV_X1 port map( A => n784, ZN => n6177);
   U1107 : AOI22_X1 port map( A1 => Set_target(0), A2 => n3446, B1 => n769, B2 
                           => pc_target_10_0_port, ZN => n784);
   U1108 : INV_X1 port map( A => n785, ZN => n6178);
   U1109 : AOI22_X1 port map( A1 => Set_target(1), A2 => n3446, B1 => n769, B2 
                           => pc_target_10_1_port, ZN => n785);
   U1110 : INV_X1 port map( A => n786, ZN => n6179);
   U1111 : AOI22_X1 port map( A1 => Set_target(3), A2 => n3446, B1 => n769, B2 
                           => pc_target_10_3_port, ZN => n786);
   U1112 : INV_X1 port map( A => n787, ZN => n6180);
   U1113 : AOI22_X1 port map( A1 => Set_target(5), A2 => n3446, B1 => n769, B2 
                           => pc_target_10_5_port, ZN => n787);
   U1114 : INV_X1 port map( A => n788, ZN => n6181);
   U1115 : AOI22_X1 port map( A1 => Set_target(7), A2 => n3446, B1 => n769, B2 
                           => pc_target_10_7_port, ZN => n788);
   U1116 : INV_X1 port map( A => n789, ZN => n6182);
   U1117 : AOI22_X1 port map( A1 => Set_target(9), A2 => n3446, B1 => n769, B2 
                           => pc_target_10_9_port, ZN => n789);
   U1118 : INV_X1 port map( A => n790, ZN => n6183);
   U1119 : AOI22_X1 port map( A1 => Set_target(11), A2 => n3446, B1 => n769, B2
                           => pc_target_10_11_port, ZN => n790);
   U1120 : INV_X1 port map( A => n791, ZN => n6184);
   U1121 : AOI22_X1 port map( A1 => Set_target(13), A2 => n3446, B1 => n769, B2
                           => pc_target_10_13_port, ZN => n791);
   U1122 : INV_X1 port map( A => n792, ZN => n6185);
   U1123 : AOI22_X1 port map( A1 => Set_target(15), A2 => n3446, B1 => n769, B2
                           => pc_target_10_15_port, ZN => n792);
   U1124 : INV_X1 port map( A => n793, ZN => n6186);
   U1125 : AOI22_X1 port map( A1 => Set_target(17), A2 => n3446, B1 => n769, B2
                           => pc_target_10_17_port, ZN => n793);
   U1126 : INV_X1 port map( A => n794, ZN => n6187);
   U1127 : AOI22_X1 port map( A1 => Set_target(19), A2 => n3446, B1 => n769, B2
                           => pc_target_10_19_port, ZN => n794);
   U1128 : INV_X1 port map( A => n795, ZN => n6188);
   U1129 : AOI22_X1 port map( A1 => Set_target(21), A2 => n3446, B1 => n769, B2
                           => pc_target_10_21_port, ZN => n795);
   U1130 : INV_X1 port map( A => n796, ZN => n6189);
   U1131 : AOI22_X1 port map( A1 => Set_target(23), A2 => n3446, B1 => n769, B2
                           => pc_target_10_23_port, ZN => n796);
   U1132 : INV_X1 port map( A => n797, ZN => n6190);
   U1133 : AOI22_X1 port map( A1 => Set_target(25), A2 => n3446, B1 => n769, B2
                           => pc_target_10_25_port, ZN => n797);
   U1134 : INV_X1 port map( A => n798, ZN => n6191);
   U1135 : AOI22_X1 port map( A1 => Set_target(27), A2 => n3446, B1 => n769, B2
                           => pc_target_10_27_port, ZN => n798);
   U1136 : INV_X1 port map( A => n799, ZN => n6192);
   U1137 : AOI22_X1 port map( A1 => Set_target(29), A2 => n3446, B1 => n769, B2
                           => pc_target_10_29_port, ZN => n799);
   U1138 : INV_X1 port map( A => n800, ZN => n6193);
   U1139 : AOI22_X1 port map( A1 => Set_target(31), A2 => n3446, B1 => n769, B2
                           => pc_target_10_31_port, ZN => n800);
   U1142 : OAI22_X1 port map( A1 => n75, A2 => n801, B1 => n3442, B2 => n803, 
                           ZN => n6194);
   U1143 : OAI22_X1 port map( A1 => n79, A2 => n801, B1 => n3442, B2 => n804, 
                           ZN => n6195);
   U1144 : OAI22_X1 port map( A1 => n81, A2 => n801, B1 => n3442, B2 => n805, 
                           ZN => n6196);
   U1145 : OAI22_X1 port map( A1 => n83, A2 => n801, B1 => n3442, B2 => n806, 
                           ZN => n6197);
   U1146 : OAI22_X1 port map( A1 => n85, A2 => n801, B1 => n3442, B2 => n807, 
                           ZN => n6198);
   U1147 : OAI22_X1 port map( A1 => n87, A2 => n801, B1 => n3442, B2 => n808, 
                           ZN => n6199);
   U1148 : OAI22_X1 port map( A1 => n89, A2 => n801, B1 => n3442, B2 => n809, 
                           ZN => n6200);
   U1149 : OAI22_X1 port map( A1 => n91, A2 => n801, B1 => n3442, B2 => n810, 
                           ZN => n6201);
   U1150 : OAI22_X1 port map( A1 => n93, A2 => n801, B1 => n3442, B2 => n811, 
                           ZN => n6202);
   U1151 : OAI22_X1 port map( A1 => n95, A2 => n801, B1 => n3442, B2 => n812, 
                           ZN => n6203);
   U1152 : OAI22_X1 port map( A1 => n97_port, A2 => n801, B1 => n3442, B2 => 
                           n813, ZN => n6204);
   U1153 : OAI22_X1 port map( A1 => n99_port, A2 => n801, B1 => n3442, B2 => 
                           n814, ZN => n6205);
   U1154 : OAI22_X1 port map( A1 => n101_port, A2 => n801, B1 => n3442, B2 => 
                           n815, ZN => n6206);
   U1155 : OAI22_X1 port map( A1 => n103_port, A2 => n801, B1 => n3442, B2 => 
                           n816, ZN => n6207);
   U1156 : OAI22_X1 port map( A1 => n105_port, A2 => n801, B1 => n3442, B2 => 
                           n817, ZN => n6208);
   U1157 : OAI22_X1 port map( A1 => n107_port, A2 => n801, B1 => n3442, B2 => 
                           n818, ZN => n6209);
   U1158 : OAI22_X1 port map( A1 => n109_port, A2 => n801, B1 => n3442, B2 => 
                           n819, ZN => n6210);
   U1159 : OAI22_X1 port map( A1 => n111_port, A2 => n801, B1 => n3442, B2 => 
                           n820, ZN => n6211);
   U1160 : OAI22_X1 port map( A1 => n113_port, A2 => n801, B1 => n3442, B2 => 
                           n821, ZN => n6212);
   U1161 : OAI22_X1 port map( A1 => n115_port, A2 => n801, B1 => n3442, B2 => 
                           n822, ZN => n6213);
   U1162 : OAI22_X1 port map( A1 => n117_port, A2 => n801, B1 => n3442, B2 => 
                           n823, ZN => n6214);
   U1163 : OAI22_X1 port map( A1 => n119_port, A2 => n801, B1 => n3442, B2 => 
                           n824, ZN => n6215);
   U1164 : OAI22_X1 port map( A1 => n121_port, A2 => n801, B1 => n3442, B2 => 
                           n825, ZN => n6216);
   U1165 : OAI22_X1 port map( A1 => n123_port, A2 => n801, B1 => n3442, B2 => 
                           n826, ZN => n6217);
   U1166 : OAI22_X1 port map( A1 => n125_port, A2 => n801, B1 => n3442, B2 => 
                           n827, ZN => n6218);
   U1167 : OAI22_X1 port map( A1 => n127_port, A2 => n801, B1 => n3442, B2 => 
                           n828, ZN => n6219);
   U1168 : OAI22_X1 port map( A1 => n129, A2 => n801, B1 => n3442, B2 => n829, 
                           ZN => n6220);
   U1169 : OAI22_X1 port map( A1 => n131, A2 => n801, B1 => n3442, B2 => n830, 
                           ZN => n6221);
   U1170 : OAI22_X1 port map( A1 => n133, A2 => n801, B1 => n3442, B2 => n831, 
                           ZN => n6222);
   U1171 : OAI22_X1 port map( A1 => n135, A2 => n801, B1 => n3442, B2 => n832, 
                           ZN => n6223);
   U1172 : OAI22_X1 port map( A1 => n137, A2 => n801, B1 => n3442, B2 => n833, 
                           ZN => n6224);
   U1173 : OAI22_X1 port map( A1 => n139, A2 => n801, B1 => n3442, B2 => n834, 
                           ZN => n6225);
   U1176 : OAI22_X1 port map( A1 => n75, A2 => n835, B1 => n836, B2 => n837, ZN
                           => n6226);
   U1177 : OAI22_X1 port map( A1 => n79, A2 => n835, B1 => n836, B2 => n838, ZN
                           => n6227);
   U1178 : OAI22_X1 port map( A1 => n81, A2 => n835, B1 => n836, B2 => n839, ZN
                           => n6228);
   U1179 : OAI22_X1 port map( A1 => n83, A2 => n835, B1 => n836, B2 => n840, ZN
                           => n6229);
   U1180 : OAI22_X1 port map( A1 => n85, A2 => n835, B1 => n836, B2 => n841, ZN
                           => n6230);
   U1181 : OAI22_X1 port map( A1 => n87, A2 => n835, B1 => n836, B2 => n842, ZN
                           => n6231);
   U1182 : OAI22_X1 port map( A1 => n89, A2 => n835, B1 => n836, B2 => n843, ZN
                           => n6232);
   U1183 : OAI22_X1 port map( A1 => n91, A2 => n835, B1 => n836, B2 => n844, ZN
                           => n6233);
   U1184 : OAI22_X1 port map( A1 => n93, A2 => n835, B1 => n836, B2 => n845, ZN
                           => n6234);
   U1185 : OAI22_X1 port map( A1 => n95, A2 => n835, B1 => n836, B2 => n846, ZN
                           => n6235);
   U1186 : OAI22_X1 port map( A1 => n97_port, A2 => n835, B1 => n836, B2 => 
                           n847, ZN => n6236);
   U1187 : OAI22_X1 port map( A1 => n99_port, A2 => n835, B1 => n836, B2 => 
                           n848, ZN => n6237);
   U1188 : OAI22_X1 port map( A1 => n101_port, A2 => n835, B1 => n836, B2 => 
                           n849, ZN => n6238);
   U1189 : OAI22_X1 port map( A1 => n103_port, A2 => n835, B1 => n836, B2 => 
                           n850, ZN => n6239);
   U1190 : OAI22_X1 port map( A1 => n105_port, A2 => n835, B1 => n836, B2 => 
                           n851, ZN => n6240);
   U1191 : OAI22_X1 port map( A1 => n107_port, A2 => n835, B1 => n836, B2 => 
                           n852, ZN => n6241);
   U1192 : OAI22_X1 port map( A1 => n109_port, A2 => n835, B1 => n836, B2 => 
                           n853, ZN => n6242);
   U1193 : OAI22_X1 port map( A1 => n111_port, A2 => n835, B1 => n836, B2 => 
                           n854, ZN => n6243);
   U1194 : OAI22_X1 port map( A1 => n113_port, A2 => n835, B1 => n836, B2 => 
                           n855, ZN => n6244);
   U1195 : OAI22_X1 port map( A1 => n115_port, A2 => n835, B1 => n836, B2 => 
                           n856, ZN => n6245);
   U1196 : OAI22_X1 port map( A1 => n117_port, A2 => n835, B1 => n836, B2 => 
                           n857, ZN => n6246);
   U1197 : OAI22_X1 port map( A1 => n119_port, A2 => n835, B1 => n836, B2 => 
                           n858, ZN => n6247);
   U1198 : OAI22_X1 port map( A1 => n121_port, A2 => n835, B1 => n836, B2 => 
                           n859, ZN => n6248);
   U1199 : OAI22_X1 port map( A1 => n123_port, A2 => n835, B1 => n836, B2 => 
                           n860, ZN => n6249);
   U1200 : OAI22_X1 port map( A1 => n125_port, A2 => n835, B1 => n836, B2 => 
                           n861, ZN => n6250);
   U1201 : OAI22_X1 port map( A1 => n127_port, A2 => n835, B1 => n836, B2 => 
                           n862, ZN => n6251);
   U1202 : OAI22_X1 port map( A1 => n129, A2 => n835, B1 => n836, B2 => n863, 
                           ZN => n6252);
   U1203 : OAI22_X1 port map( A1 => n131, A2 => n835, B1 => n836, B2 => n864, 
                           ZN => n6253);
   U1204 : OAI22_X1 port map( A1 => n133, A2 => n835, B1 => n836, B2 => n865, 
                           ZN => n6254);
   U1205 : OAI22_X1 port map( A1 => n135, A2 => n835, B1 => n836, B2 => n866, 
                           ZN => n6255);
   U1206 : OAI22_X1 port map( A1 => n137, A2 => n835, B1 => n836, B2 => n867, 
                           ZN => n6256);
   U1207 : OAI22_X1 port map( A1 => n139, A2 => n835, B1 => n836, B2 => n868, 
                           ZN => n6257);
   U1211 : INV_X1 port map( A => n869, ZN => n6258);
   U1212 : AOI22_X1 port map( A1 => Set_target(30), A2 => n870, B1 => n1656, B2
                           => pc_target_7_30_port, ZN => n869);
   U1213 : INV_X1 port map( A => n872, ZN => n6259);
   U1214 : AOI22_X1 port map( A1 => Set_target(28), A2 => n870, B1 => n1656, B2
                           => pc_target_7_28_port, ZN => n872);
   U1215 : INV_X1 port map( A => n873, ZN => n6260);
   U1216 : AOI22_X1 port map( A1 => Set_target(26), A2 => n870, B1 => n1611, B2
                           => pc_target_7_26_port, ZN => n873);
   U1217 : INV_X1 port map( A => n874, ZN => n6261);
   U1218 : AOI22_X1 port map( A1 => Set_target(24), A2 => n870, B1 => n1656, B2
                           => pc_target_7_24_port, ZN => n874);
   U1219 : INV_X1 port map( A => n875, ZN => n6262);
   U1220 : AOI22_X1 port map( A1 => Set_target(22), A2 => n870, B1 => n1656, B2
                           => pc_target_7_22_port, ZN => n875);
   U1221 : INV_X1 port map( A => n876, ZN => n6263);
   U1222 : AOI22_X1 port map( A1 => Set_target(20), A2 => n870, B1 => n1656, B2
                           => pc_target_7_20_port, ZN => n876);
   U1223 : INV_X1 port map( A => n877, ZN => n6264);
   U1224 : AOI22_X1 port map( A1 => Set_target(18), A2 => n870, B1 => n1656, B2
                           => pc_target_7_18_port, ZN => n877);
   U1225 : INV_X1 port map( A => n878, ZN => n6265);
   U1226 : AOI22_X1 port map( A1 => Set_target(16), A2 => n870, B1 => n1656, B2
                           => pc_target_7_16_port, ZN => n878);
   U1227 : INV_X1 port map( A => n879, ZN => n6266);
   U1228 : AOI22_X1 port map( A1 => Set_target(14), A2 => n870, B1 => n1611, B2
                           => pc_target_7_14_port, ZN => n879);
   U1229 : INV_X1 port map( A => n880, ZN => n6267);
   U1230 : AOI22_X1 port map( A1 => Set_target(12), A2 => n870, B1 => n1656, B2
                           => pc_target_7_12_port, ZN => n880);
   U1231 : INV_X1 port map( A => n881, ZN => n6268);
   U1232 : AOI22_X1 port map( A1 => Set_target(10), A2 => n870, B1 => n1656, B2
                           => pc_target_7_10_port, ZN => n881);
   U1233 : INV_X1 port map( A => n882, ZN => n6269);
   U1234 : AOI22_X1 port map( A1 => Set_target(8), A2 => n870, B1 => n1656, B2 
                           => pc_target_7_8_port, ZN => n882);
   U1235 : INV_X1 port map( A => n883, ZN => n6270);
   U1236 : AOI22_X1 port map( A1 => Set_target(6), A2 => n870, B1 => n1656, B2 
                           => pc_target_7_6_port, ZN => n883);
   U1237 : INV_X1 port map( A => n884, ZN => n6271);
   U1238 : AOI22_X1 port map( A1 => Set_target(4), A2 => n870, B1 => n1656, B2 
                           => pc_target_7_4_port, ZN => n884);
   U1239 : INV_X1 port map( A => n885, ZN => n6272);
   U1240 : AOI22_X1 port map( A1 => Set_target(2), A2 => n870, B1 => n1656, B2 
                           => pc_target_7_2_port, ZN => n885);
   U1241 : INV_X1 port map( A => n886, ZN => n6273);
   U1242 : AOI22_X1 port map( A1 => Set_target(0), A2 => n870, B1 => n1656, B2 
                           => pc_target_7_0_port, ZN => n886);
   U1243 : INV_X1 port map( A => n887, ZN => n6274);
   U1244 : AOI22_X1 port map( A1 => Set_target(1), A2 => n870, B1 => n1656, B2 
                           => pc_target_7_1_port, ZN => n887);
   U1245 : INV_X1 port map( A => n888, ZN => n6275);
   U1246 : AOI22_X1 port map( A1 => Set_target(3), A2 => n870, B1 => n1656, B2 
                           => pc_target_7_3_port, ZN => n888);
   U1247 : INV_X1 port map( A => n889, ZN => n6276);
   U1248 : AOI22_X1 port map( A1 => Set_target(5), A2 => n870, B1 => n1656, B2 
                           => pc_target_7_5_port, ZN => n889);
   U1249 : INV_X1 port map( A => n890, ZN => n6277);
   U1250 : AOI22_X1 port map( A1 => Set_target(7), A2 => n870, B1 => n1656, B2 
                           => pc_target_7_7_port, ZN => n890);
   U1251 : INV_X1 port map( A => n891, ZN => n6278);
   U1252 : AOI22_X1 port map( A1 => Set_target(9), A2 => n870, B1 => n1656, B2 
                           => pc_target_7_9_port, ZN => n891);
   U1253 : INV_X1 port map( A => n892, ZN => n6279);
   U1254 : AOI22_X1 port map( A1 => Set_target(11), A2 => n870, B1 => n1611, B2
                           => pc_target_7_11_port, ZN => n892);
   U1255 : INV_X1 port map( A => n893, ZN => n6280);
   U1256 : AOI22_X1 port map( A1 => Set_target(13), A2 => n870, B1 => n1656, B2
                           => pc_target_7_13_port, ZN => n893);
   U1257 : INV_X1 port map( A => n894, ZN => n6281);
   U1258 : AOI22_X1 port map( A1 => Set_target(15), A2 => n870, B1 => n1656, B2
                           => pc_target_7_15_port, ZN => n894);
   U1259 : INV_X1 port map( A => n895, ZN => n6282);
   U1260 : AOI22_X1 port map( A1 => Set_target(17), A2 => n870, B1 => n1656, B2
                           => pc_target_7_17_port, ZN => n895);
   U1261 : INV_X1 port map( A => n896, ZN => n6283);
   U1262 : AOI22_X1 port map( A1 => Set_target(19), A2 => n870, B1 => n1611, B2
                           => pc_target_7_19_port, ZN => n896);
   U1263 : INV_X1 port map( A => n897, ZN => n6284);
   U1264 : AOI22_X1 port map( A1 => Set_target(21), A2 => n870, B1 => n1656, B2
                           => pc_target_7_21_port, ZN => n897);
   U1265 : INV_X1 port map( A => n898, ZN => n6285);
   U1266 : AOI22_X1 port map( A1 => Set_target(23), A2 => n870, B1 => n1611, B2
                           => pc_target_7_23_port, ZN => n898);
   U1267 : INV_X1 port map( A => n899, ZN => n6286);
   U1268 : AOI22_X1 port map( A1 => Set_target(25), A2 => n870, B1 => n1656, B2
                           => pc_target_7_25_port, ZN => n899);
   U1269 : INV_X1 port map( A => n900, ZN => n6287);
   U1270 : AOI22_X1 port map( A1 => Set_target(27), A2 => n870, B1 => n1656, B2
                           => pc_target_7_27_port, ZN => n900);
   U1271 : INV_X1 port map( A => n901, ZN => n6288);
   U1272 : AOI22_X1 port map( A1 => Set_target(29), A2 => n870, B1 => n1656, B2
                           => pc_target_7_29_port, ZN => n901);
   U1273 : INV_X1 port map( A => n902, ZN => n6289);
   U1274 : AOI22_X1 port map( A1 => Set_target(31), A2 => n870, B1 => n1611, B2
                           => pc_target_7_31_port, ZN => n902);
   U1277 : INV_X1 port map( A => n904, ZN => n6290);
   U1278 : AOI22_X1 port map( A1 => Set_target(30), A2 => n905, B1 => n906, B2 
                           => pc_target_6_30_port, ZN => n904);
   U1279 : INV_X1 port map( A => n907, ZN => n6291);
   U1280 : AOI22_X1 port map( A1 => Set_target(28), A2 => n905, B1 => n906, B2 
                           => pc_target_6_28_port, ZN => n907);
   U1281 : INV_X1 port map( A => n908, ZN => n6292);
   U1282 : AOI22_X1 port map( A1 => Set_target(26), A2 => n905, B1 => n906, B2 
                           => pc_target_6_26_port, ZN => n908);
   U1283 : INV_X1 port map( A => n909, ZN => n6293);
   U1284 : AOI22_X1 port map( A1 => Set_target(24), A2 => n905, B1 => n906, B2 
                           => pc_target_6_24_port, ZN => n909);
   U1285 : INV_X1 port map( A => n910, ZN => n6294);
   U1286 : AOI22_X1 port map( A1 => Set_target(22), A2 => n905, B1 => n906, B2 
                           => pc_target_6_22_port, ZN => n910);
   U1287 : INV_X1 port map( A => n911, ZN => n6295);
   U1288 : AOI22_X1 port map( A1 => Set_target(20), A2 => n905, B1 => n906, B2 
                           => pc_target_6_20_port, ZN => n911);
   U1289 : INV_X1 port map( A => n912, ZN => n6296);
   U1290 : AOI22_X1 port map( A1 => Set_target(18), A2 => n905, B1 => n906, B2 
                           => pc_target_6_18_port, ZN => n912);
   U1291 : INV_X1 port map( A => n913, ZN => n6297);
   U1292 : AOI22_X1 port map( A1 => Set_target(16), A2 => n905, B1 => n906, B2 
                           => pc_target_6_16_port, ZN => n913);
   U1293 : INV_X1 port map( A => n914, ZN => n6298);
   U1294 : AOI22_X1 port map( A1 => Set_target(14), A2 => n905, B1 => n906, B2 
                           => pc_target_6_14_port, ZN => n914);
   U1295 : INV_X1 port map( A => n915, ZN => n6299);
   U1296 : AOI22_X1 port map( A1 => Set_target(12), A2 => n905, B1 => n906, B2 
                           => pc_target_6_12_port, ZN => n915);
   U1297 : INV_X1 port map( A => n916, ZN => n6300);
   U1298 : AOI22_X1 port map( A1 => Set_target(10), A2 => n905, B1 => n906, B2 
                           => pc_target_6_10_port, ZN => n916);
   U1299 : INV_X1 port map( A => n917, ZN => n6301);
   U1300 : AOI22_X1 port map( A1 => Set_target(8), A2 => n905, B1 => n906, B2 
                           => pc_target_6_8_port, ZN => n917);
   U1301 : INV_X1 port map( A => n918, ZN => n6302);
   U1302 : AOI22_X1 port map( A1 => Set_target(6), A2 => n905, B1 => n906, B2 
                           => pc_target_6_6_port, ZN => n918);
   U1303 : INV_X1 port map( A => n919, ZN => n6303);
   U1304 : AOI22_X1 port map( A1 => Set_target(4), A2 => n905, B1 => n906, B2 
                           => pc_target_6_4_port, ZN => n919);
   U1305 : INV_X1 port map( A => n920, ZN => n6304);
   U1306 : AOI22_X1 port map( A1 => Set_target(2), A2 => n905, B1 => n906, B2 
                           => pc_target_6_2_port, ZN => n920);
   U1307 : INV_X1 port map( A => n921, ZN => n6305);
   U1308 : AOI22_X1 port map( A1 => Set_target(0), A2 => n905, B1 => n906, B2 
                           => pc_target_6_0_port, ZN => n921);
   U1309 : INV_X1 port map( A => n922, ZN => n6306);
   U1310 : AOI22_X1 port map( A1 => Set_target(1), A2 => n905, B1 => n906, B2 
                           => pc_target_6_1_port, ZN => n922);
   U1311 : INV_X1 port map( A => n923, ZN => n6307);
   U1312 : AOI22_X1 port map( A1 => Set_target(3), A2 => n905, B1 => n906, B2 
                           => pc_target_6_3_port, ZN => n923);
   U1313 : INV_X1 port map( A => n924, ZN => n6308);
   U1314 : AOI22_X1 port map( A1 => Set_target(5), A2 => n905, B1 => n906, B2 
                           => pc_target_6_5_port, ZN => n924);
   U1315 : INV_X1 port map( A => n925, ZN => n6309);
   U1316 : AOI22_X1 port map( A1 => Set_target(7), A2 => n905, B1 => n906, B2 
                           => pc_target_6_7_port, ZN => n925);
   U1317 : INV_X1 port map( A => n926, ZN => n6310);
   U1318 : AOI22_X1 port map( A1 => Set_target(9), A2 => n905, B1 => n906, B2 
                           => pc_target_6_9_port, ZN => n926);
   U1319 : INV_X1 port map( A => n927, ZN => n6311);
   U1320 : AOI22_X1 port map( A1 => Set_target(11), A2 => n905, B1 => n906, B2 
                           => pc_target_6_11_port, ZN => n927);
   U1321 : INV_X1 port map( A => n928, ZN => n6312);
   U1322 : AOI22_X1 port map( A1 => Set_target(13), A2 => n905, B1 => n906, B2 
                           => pc_target_6_13_port, ZN => n928);
   U1323 : INV_X1 port map( A => n929, ZN => n6313);
   U1324 : AOI22_X1 port map( A1 => Set_target(15), A2 => n905, B1 => n906, B2 
                           => pc_target_6_15_port, ZN => n929);
   U1325 : INV_X1 port map( A => n930, ZN => n6314);
   U1326 : AOI22_X1 port map( A1 => Set_target(17), A2 => n905, B1 => n906, B2 
                           => pc_target_6_17_port, ZN => n930);
   U1327 : INV_X1 port map( A => n931, ZN => n6315);
   U1328 : AOI22_X1 port map( A1 => Set_target(19), A2 => n905, B1 => n906, B2 
                           => pc_target_6_19_port, ZN => n931);
   U1329 : INV_X1 port map( A => n932, ZN => n6316);
   U1330 : AOI22_X1 port map( A1 => Set_target(21), A2 => n905, B1 => n906, B2 
                           => pc_target_6_21_port, ZN => n932);
   U1331 : INV_X1 port map( A => n933, ZN => n6317);
   U1332 : AOI22_X1 port map( A1 => Set_target(23), A2 => n905, B1 => n906, B2 
                           => pc_target_6_23_port, ZN => n933);
   U1333 : INV_X1 port map( A => n934, ZN => n6318);
   U1334 : AOI22_X1 port map( A1 => Set_target(25), A2 => n905, B1 => n906, B2 
                           => pc_target_6_25_port, ZN => n934);
   U1335 : INV_X1 port map( A => n935, ZN => n6319);
   U1336 : AOI22_X1 port map( A1 => Set_target(27), A2 => n905, B1 => n906, B2 
                           => pc_target_6_27_port, ZN => n935);
   U1337 : INV_X1 port map( A => n936, ZN => n6320);
   U1338 : AOI22_X1 port map( A1 => Set_target(29), A2 => n905, B1 => n906, B2 
                           => pc_target_6_29_port, ZN => n936);
   U1339 : INV_X1 port map( A => n937, ZN => n6321);
   U1340 : AOI22_X1 port map( A1 => Set_target(31), A2 => n905, B1 => n906, B2 
                           => pc_target_6_31_port, ZN => n937);
   U1343 : OAI22_X1 port map( A1 => n75, A2 => n938, B1 => n939, B2 => n940, ZN
                           => n6322);
   U1344 : OAI22_X1 port map( A1 => n79, A2 => n938, B1 => n939, B2 => n941, ZN
                           => n6323);
   U1345 : OAI22_X1 port map( A1 => n81, A2 => n938, B1 => n939, B2 => n942, ZN
                           => n6324);
   U1346 : OAI22_X1 port map( A1 => n83, A2 => n938, B1 => n939, B2 => n943, ZN
                           => n6325);
   U1347 : OAI22_X1 port map( A1 => n85, A2 => n938, B1 => n939, B2 => n944, ZN
                           => n6326);
   U1348 : OAI22_X1 port map( A1 => n87, A2 => n938, B1 => n939, B2 => n945, ZN
                           => n6327);
   U1349 : OAI22_X1 port map( A1 => n89, A2 => n938, B1 => n939, B2 => n946, ZN
                           => n6328);
   U1350 : OAI22_X1 port map( A1 => n91, A2 => n938, B1 => n939, B2 => n947, ZN
                           => n6329);
   U1351 : OAI22_X1 port map( A1 => n93, A2 => n938, B1 => n939, B2 => n948, ZN
                           => n6330);
   U1352 : OAI22_X1 port map( A1 => n95, A2 => n938, B1 => n939, B2 => n949, ZN
                           => n6331);
   U1353 : OAI22_X1 port map( A1 => n97_port, A2 => n938, B1 => n939, B2 => 
                           n950, ZN => n6332);
   U1354 : OAI22_X1 port map( A1 => n99_port, A2 => n938, B1 => n939, B2 => 
                           n951, ZN => n6333);
   U1355 : OAI22_X1 port map( A1 => n101_port, A2 => n938, B1 => n939, B2 => 
                           n952, ZN => n6334);
   U1356 : OAI22_X1 port map( A1 => n103_port, A2 => n938, B1 => n939, B2 => 
                           n953, ZN => n6335);
   U1357 : OAI22_X1 port map( A1 => n105_port, A2 => n938, B1 => n939, B2 => 
                           n954, ZN => n6336);
   U1358 : OAI22_X1 port map( A1 => n107_port, A2 => n938, B1 => n939, B2 => 
                           n955, ZN => n6337);
   U1359 : OAI22_X1 port map( A1 => n109_port, A2 => n938, B1 => n939, B2 => 
                           n956, ZN => n6338);
   U1360 : OAI22_X1 port map( A1 => n111_port, A2 => n938, B1 => n939, B2 => 
                           n957, ZN => n6339);
   U1361 : OAI22_X1 port map( A1 => n113_port, A2 => n938, B1 => n939, B2 => 
                           n958, ZN => n6340);
   U1362 : OAI22_X1 port map( A1 => n115_port, A2 => n938, B1 => n939, B2 => 
                           n959, ZN => n6341);
   U1363 : OAI22_X1 port map( A1 => n117_port, A2 => n938, B1 => n939, B2 => 
                           n960, ZN => n6342);
   U1364 : OAI22_X1 port map( A1 => n119_port, A2 => n938, B1 => n939, B2 => 
                           n961, ZN => n6343);
   U1365 : OAI22_X1 port map( A1 => n121_port, A2 => n938, B1 => n939, B2 => 
                           n962, ZN => n6344);
   U1366 : OAI22_X1 port map( A1 => n123_port, A2 => n938, B1 => n939, B2 => 
                           n963, ZN => n6345);
   U1367 : OAI22_X1 port map( A1 => n125_port, A2 => n938, B1 => n939, B2 => 
                           n964, ZN => n6346);
   U1368 : OAI22_X1 port map( A1 => n127_port, A2 => n938, B1 => n939, B2 => 
                           n965, ZN => n6347);
   U1369 : OAI22_X1 port map( A1 => n129, A2 => n938, B1 => n939, B2 => n966, 
                           ZN => n6348);
   U1370 : OAI22_X1 port map( A1 => n131, A2 => n938, B1 => n939, B2 => n967, 
                           ZN => n6349);
   U1371 : OAI22_X1 port map( A1 => n133, A2 => n938, B1 => n939, B2 => n968, 
                           ZN => n6350);
   U1372 : OAI22_X1 port map( A1 => n135, A2 => n938, B1 => n939, B2 => n969, 
                           ZN => n6351);
   U1373 : OAI22_X1 port map( A1 => n137, A2 => n938, B1 => n939, B2 => n970, 
                           ZN => n6352);
   U1374 : OAI22_X1 port map( A1 => n139, A2 => n938, B1 => n939, B2 => n971, 
                           ZN => n6353);
   U1377 : OAI22_X1 port map( A1 => n75, A2 => n972, B1 => n3443, B2 => n974, 
                           ZN => n6354);
   U1378 : OAI22_X1 port map( A1 => n79, A2 => n972, B1 => n3443, B2 => n975, 
                           ZN => n6355);
   U1379 : OAI22_X1 port map( A1 => n81, A2 => n972, B1 => n3443, B2 => n976, 
                           ZN => n6356);
   U1380 : OAI22_X1 port map( A1 => n83, A2 => n972, B1 => n3443, B2 => n977, 
                           ZN => n6357);
   U1381 : OAI22_X1 port map( A1 => n85, A2 => n972, B1 => n3443, B2 => n978, 
                           ZN => n6358);
   U1382 : OAI22_X1 port map( A1 => n87, A2 => n972, B1 => n3443, B2 => n979, 
                           ZN => n6359);
   U1383 : OAI22_X1 port map( A1 => n89, A2 => n972, B1 => n3443, B2 => n980, 
                           ZN => n6360);
   U1384 : OAI22_X1 port map( A1 => n91, A2 => n972, B1 => n3443, B2 => n981, 
                           ZN => n6361);
   U1385 : OAI22_X1 port map( A1 => n93, A2 => n972, B1 => n3443, B2 => n982, 
                           ZN => n6362);
   U1386 : OAI22_X1 port map( A1 => n95, A2 => n972, B1 => n3443, B2 => n983, 
                           ZN => n6363);
   U1387 : OAI22_X1 port map( A1 => n97_port, A2 => n972, B1 => n3443, B2 => 
                           n984, ZN => n6364);
   U1388 : OAI22_X1 port map( A1 => n99_port, A2 => n972, B1 => n3443, B2 => 
                           n985, ZN => n6365);
   U1389 : OAI22_X1 port map( A1 => n101_port, A2 => n972, B1 => n3443, B2 => 
                           n986, ZN => n6366);
   U1390 : OAI22_X1 port map( A1 => n103_port, A2 => n972, B1 => n3443, B2 => 
                           n987, ZN => n6367);
   U1391 : OAI22_X1 port map( A1 => n105_port, A2 => n972, B1 => n3443, B2 => 
                           n988, ZN => n6368);
   U1392 : OAI22_X1 port map( A1 => n107_port, A2 => n972, B1 => n3443, B2 => 
                           n989, ZN => n6369);
   U1393 : OAI22_X1 port map( A1 => n109_port, A2 => n972, B1 => n3443, B2 => 
                           n990, ZN => n6370);
   U1394 : OAI22_X1 port map( A1 => n111_port, A2 => n972, B1 => n3443, B2 => 
                           n991, ZN => n6371);
   U1395 : OAI22_X1 port map( A1 => n113_port, A2 => n972, B1 => n3443, B2 => 
                           n992, ZN => n6372);
   U1396 : OAI22_X1 port map( A1 => n115_port, A2 => n972, B1 => n3443, B2 => 
                           n993, ZN => n6373);
   U1397 : OAI22_X1 port map( A1 => n117_port, A2 => n972, B1 => n3443, B2 => 
                           n994, ZN => n6374);
   U1398 : OAI22_X1 port map( A1 => n119_port, A2 => n972, B1 => n3443, B2 => 
                           n995, ZN => n6375);
   U1399 : OAI22_X1 port map( A1 => n121_port, A2 => n972, B1 => n3443, B2 => 
                           n996, ZN => n6376);
   U1400 : OAI22_X1 port map( A1 => n123_port, A2 => n972, B1 => n3443, B2 => 
                           n997, ZN => n6377);
   U1401 : OAI22_X1 port map( A1 => n125_port, A2 => n972, B1 => n3443, B2 => 
                           n998, ZN => n6378);
   U1402 : OAI22_X1 port map( A1 => n127_port, A2 => n972, B1 => n3443, B2 => 
                           n999, ZN => n6379);
   U1403 : OAI22_X1 port map( A1 => n129, A2 => n972, B1 => n3443, B2 => n1000,
                           ZN => n6380);
   U1404 : OAI22_X1 port map( A1 => n131, A2 => n972, B1 => n3443, B2 => n1001,
                           ZN => n6381);
   U1405 : OAI22_X1 port map( A1 => n133, A2 => n972, B1 => n3443, B2 => n1002,
                           ZN => n6382);
   U1406 : OAI22_X1 port map( A1 => n135, A2 => n972, B1 => n3443, B2 => n1003,
                           ZN => n6383);
   U1407 : OAI22_X1 port map( A1 => n137, A2 => n972, B1 => n3443, B2 => n1004,
                           ZN => n6384);
   U1408 : OAI22_X1 port map( A1 => n139, A2 => n972, B1 => n3443, B2 => n1005,
                           ZN => n6385);
   U1412 : INV_X1 port map( A => n1006, ZN => n6386);
   U1413 : AOI22_X1 port map( A1 => Set_target(30), A2 => n1007, B1 => n1008, 
                           B2 => pc_target_3_30_port, ZN => n1006);
   U1414 : INV_X1 port map( A => n1009, ZN => n6387);
   U1415 : AOI22_X1 port map( A1 => Set_target(28), A2 => n1007, B1 => n1008, 
                           B2 => pc_target_3_28_port, ZN => n1009);
   U1416 : INV_X1 port map( A => n1010, ZN => n6388);
   U1417 : AOI22_X1 port map( A1 => Set_target(26), A2 => n1007, B1 => n1008, 
                           B2 => pc_target_3_26_port, ZN => n1010);
   U1418 : INV_X1 port map( A => n1011, ZN => n6389);
   U1419 : AOI22_X1 port map( A1 => Set_target(24), A2 => n1007, B1 => n1008, 
                           B2 => pc_target_3_24_port, ZN => n1011);
   U1420 : INV_X1 port map( A => n1012, ZN => n6390);
   U1421 : AOI22_X1 port map( A1 => Set_target(22), A2 => n1007, B1 => n1008, 
                           B2 => pc_target_3_22_port, ZN => n1012);
   U1422 : INV_X1 port map( A => n1013, ZN => n6391);
   U1423 : AOI22_X1 port map( A1 => Set_target(20), A2 => n1007, B1 => n1008, 
                           B2 => pc_target_3_20_port, ZN => n1013);
   U1424 : INV_X1 port map( A => n1014, ZN => n6392);
   U1425 : AOI22_X1 port map( A1 => Set_target(18), A2 => n1007, B1 => n1008, 
                           B2 => pc_target_3_18_port, ZN => n1014);
   U1426 : INV_X1 port map( A => n1015, ZN => n6393);
   U1427 : AOI22_X1 port map( A1 => Set_target(16), A2 => n1007, B1 => n1008, 
                           B2 => pc_target_3_16_port, ZN => n1015);
   U1428 : INV_X1 port map( A => n1016, ZN => n6394);
   U1429 : AOI22_X1 port map( A1 => Set_target(14), A2 => n1007, B1 => n1008, 
                           B2 => pc_target_3_14_port, ZN => n1016);
   U1430 : INV_X1 port map( A => n1017, ZN => n6395);
   U1431 : AOI22_X1 port map( A1 => Set_target(12), A2 => n1007, B1 => n1008, 
                           B2 => pc_target_3_12_port, ZN => n1017);
   U1432 : INV_X1 port map( A => n1018, ZN => n6396);
   U1433 : AOI22_X1 port map( A1 => Set_target(10), A2 => n1007, B1 => n1008, 
                           B2 => pc_target_3_10_port, ZN => n1018);
   U1434 : INV_X1 port map( A => n1019, ZN => n6397);
   U1435 : AOI22_X1 port map( A1 => Set_target(8), A2 => n1007, B1 => n1008, B2
                           => pc_target_3_8_port, ZN => n1019);
   U1436 : INV_X1 port map( A => n1020, ZN => n6398);
   U1437 : AOI22_X1 port map( A1 => Set_target(6), A2 => n1007, B1 => n1008, B2
                           => pc_target_3_6_port, ZN => n1020);
   U1438 : INV_X1 port map( A => n1021, ZN => n6399);
   U1439 : AOI22_X1 port map( A1 => Set_target(4), A2 => n1007, B1 => n1008, B2
                           => pc_target_3_4_port, ZN => n1021);
   U1440 : INV_X1 port map( A => n1022, ZN => n6400);
   U1441 : AOI22_X1 port map( A1 => Set_target(2), A2 => n1007, B1 => n1008, B2
                           => pc_target_3_2_port, ZN => n1022);
   U1442 : INV_X1 port map( A => n1023, ZN => n6401);
   U1443 : AOI22_X1 port map( A1 => Set_target(0), A2 => n1007, B1 => n1008, B2
                           => pc_target_3_0_port, ZN => n1023);
   U1444 : INV_X1 port map( A => n1024, ZN => n6402);
   U1445 : AOI22_X1 port map( A1 => Set_target(1), A2 => n1007, B1 => n1008, B2
                           => pc_target_3_1_port, ZN => n1024);
   U1446 : INV_X1 port map( A => n1025, ZN => n6403);
   U1447 : AOI22_X1 port map( A1 => Set_target(3), A2 => n1007, B1 => n1008, B2
                           => pc_target_3_3_port, ZN => n1025);
   U1448 : INV_X1 port map( A => n1026, ZN => n6404);
   U1449 : AOI22_X1 port map( A1 => Set_target(5), A2 => n1007, B1 => n1008, B2
                           => pc_target_3_5_port, ZN => n1026);
   U1450 : INV_X1 port map( A => n1027, ZN => n6405);
   U1451 : AOI22_X1 port map( A1 => Set_target(7), A2 => n1007, B1 => n1008, B2
                           => pc_target_3_7_port, ZN => n1027);
   U1452 : INV_X1 port map( A => n1028, ZN => n6406);
   U1453 : AOI22_X1 port map( A1 => Set_target(9), A2 => n1007, B1 => n1008, B2
                           => pc_target_3_9_port, ZN => n1028);
   U1454 : INV_X1 port map( A => n1029, ZN => n6407);
   U1455 : AOI22_X1 port map( A1 => Set_target(11), A2 => n1007, B1 => n1008, 
                           B2 => pc_target_3_11_port, ZN => n1029);
   U1456 : INV_X1 port map( A => n1030, ZN => n6408);
   U1457 : AOI22_X1 port map( A1 => Set_target(13), A2 => n1007, B1 => n1008, 
                           B2 => pc_target_3_13_port, ZN => n1030);
   U1458 : INV_X1 port map( A => n1031, ZN => n6409);
   U1459 : AOI22_X1 port map( A1 => Set_target(15), A2 => n1007, B1 => n1008, 
                           B2 => pc_target_3_15_port, ZN => n1031);
   U1460 : INV_X1 port map( A => n1032, ZN => n6410);
   U1461 : AOI22_X1 port map( A1 => Set_target(17), A2 => n1007, B1 => n1008, 
                           B2 => pc_target_3_17_port, ZN => n1032);
   U1462 : INV_X1 port map( A => n1033, ZN => n6411);
   U1463 : AOI22_X1 port map( A1 => Set_target(19), A2 => n1007, B1 => n1008, 
                           B2 => pc_target_3_19_port, ZN => n1033);
   U1464 : INV_X1 port map( A => n1034, ZN => n6412);
   U1465 : AOI22_X1 port map( A1 => Set_target(21), A2 => n1007, B1 => n1008, 
                           B2 => pc_target_3_21_port, ZN => n1034);
   U1466 : INV_X1 port map( A => n1035, ZN => n6413);
   U1467 : AOI22_X1 port map( A1 => Set_target(23), A2 => n1007, B1 => n1008, 
                           B2 => pc_target_3_23_port, ZN => n1035);
   U1468 : INV_X1 port map( A => n1036, ZN => n6414);
   U1469 : AOI22_X1 port map( A1 => Set_target(25), A2 => n1007, B1 => n1008, 
                           B2 => pc_target_3_25_port, ZN => n1036);
   U1470 : INV_X1 port map( A => n1037, ZN => n6415);
   U1471 : AOI22_X1 port map( A1 => Set_target(27), A2 => n1007, B1 => n1008, 
                           B2 => pc_target_3_27_port, ZN => n1037);
   U1472 : INV_X1 port map( A => n1038, ZN => n6416);
   U1473 : AOI22_X1 port map( A1 => Set_target(29), A2 => n1007, B1 => n1008, 
                           B2 => pc_target_3_29_port, ZN => n1038);
   U1474 : INV_X1 port map( A => n1039, ZN => n6417);
   U1475 : AOI22_X1 port map( A1 => Set_target(31), A2 => n1007, B1 => n1008, 
                           B2 => pc_target_3_31_port, ZN => n1039);
   U1478 : INV_X1 port map( A => n1041, ZN => n6418);
   U1479 : AOI22_X1 port map( A1 => Set_target(30), A2 => n1042, B1 => n1043, 
                           B2 => pc_target_2_30_port, ZN => n1041);
   U1480 : INV_X1 port map( A => n1044, ZN => n6419);
   U1481 : AOI22_X1 port map( A1 => Set_target(28), A2 => n1042, B1 => n1043, 
                           B2 => pc_target_2_28_port, ZN => n1044);
   U1482 : INV_X1 port map( A => n1045, ZN => n6420);
   U1483 : AOI22_X1 port map( A1 => Set_target(26), A2 => n1042, B1 => n1043, 
                           B2 => pc_target_2_26_port, ZN => n1045);
   U1484 : INV_X1 port map( A => n1046, ZN => n6421);
   U1485 : AOI22_X1 port map( A1 => Set_target(24), A2 => n1042, B1 => n1043, 
                           B2 => pc_target_2_24_port, ZN => n1046);
   U1486 : INV_X1 port map( A => n1047, ZN => n6422);
   U1487 : AOI22_X1 port map( A1 => Set_target(22), A2 => n1042, B1 => n1043, 
                           B2 => pc_target_2_22_port, ZN => n1047);
   U1488 : INV_X1 port map( A => n1048, ZN => n6423);
   U1489 : AOI22_X1 port map( A1 => Set_target(20), A2 => n1042, B1 => n1043, 
                           B2 => pc_target_2_20_port, ZN => n1048);
   U1490 : INV_X1 port map( A => n1049, ZN => n6424);
   U1491 : AOI22_X1 port map( A1 => Set_target(18), A2 => n1042, B1 => n1043, 
                           B2 => pc_target_2_18_port, ZN => n1049);
   U1492 : INV_X1 port map( A => n1050, ZN => n6425);
   U1493 : AOI22_X1 port map( A1 => Set_target(16), A2 => n1042, B1 => n1043, 
                           B2 => pc_target_2_16_port, ZN => n1050);
   U1494 : INV_X1 port map( A => n1051, ZN => n6426);
   U1495 : AOI22_X1 port map( A1 => Set_target(14), A2 => n1042, B1 => n1043, 
                           B2 => pc_target_2_14_port, ZN => n1051);
   U1496 : INV_X1 port map( A => n1052, ZN => n6427);
   U1497 : AOI22_X1 port map( A1 => Set_target(12), A2 => n1042, B1 => n1043, 
                           B2 => pc_target_2_12_port, ZN => n1052);
   U1498 : INV_X1 port map( A => n1053, ZN => n6428);
   U1499 : AOI22_X1 port map( A1 => Set_target(10), A2 => n1042, B1 => n1043, 
                           B2 => pc_target_2_10_port, ZN => n1053);
   U1500 : INV_X1 port map( A => n1054, ZN => n6429);
   U1501 : AOI22_X1 port map( A1 => Set_target(8), A2 => n1042, B1 => n1043, B2
                           => pc_target_2_8_port, ZN => n1054);
   U1502 : INV_X1 port map( A => n1055, ZN => n6430);
   U1503 : AOI22_X1 port map( A1 => Set_target(6), A2 => n1042, B1 => n1043, B2
                           => pc_target_2_6_port, ZN => n1055);
   U1504 : INV_X1 port map( A => n1056, ZN => n6431);
   U1505 : AOI22_X1 port map( A1 => Set_target(4), A2 => n1042, B1 => n1043, B2
                           => pc_target_2_4_port, ZN => n1056);
   U1506 : INV_X1 port map( A => n1057, ZN => n6432);
   U1507 : AOI22_X1 port map( A1 => Set_target(2), A2 => n1042, B1 => n1043, B2
                           => pc_target_2_2_port, ZN => n1057);
   U1508 : INV_X1 port map( A => n1058, ZN => n6433);
   U1509 : AOI22_X1 port map( A1 => Set_target(0), A2 => n1042, B1 => n1043, B2
                           => pc_target_2_0_port, ZN => n1058);
   U1510 : INV_X1 port map( A => n1059, ZN => n6434);
   U1511 : AOI22_X1 port map( A1 => Set_target(1), A2 => n1042, B1 => n1043, B2
                           => pc_target_2_1_port, ZN => n1059);
   U1512 : INV_X1 port map( A => n1060, ZN => n6435);
   U1513 : AOI22_X1 port map( A1 => Set_target(3), A2 => n1042, B1 => n1043, B2
                           => pc_target_2_3_port, ZN => n1060);
   U1514 : INV_X1 port map( A => n1061, ZN => n6436);
   U1515 : AOI22_X1 port map( A1 => Set_target(5), A2 => n1042, B1 => n1043, B2
                           => pc_target_2_5_port, ZN => n1061);
   U1516 : INV_X1 port map( A => n1062, ZN => n6437);
   U1517 : AOI22_X1 port map( A1 => Set_target(7), A2 => n1042, B1 => n1043, B2
                           => pc_target_2_7_port, ZN => n1062);
   U1518 : INV_X1 port map( A => n1063, ZN => n6438);
   U1519 : AOI22_X1 port map( A1 => Set_target(9), A2 => n1042, B1 => n1043, B2
                           => pc_target_2_9_port, ZN => n1063);
   U1520 : INV_X1 port map( A => n1064, ZN => n6439);
   U1521 : AOI22_X1 port map( A1 => Set_target(11), A2 => n1042, B1 => n1043, 
                           B2 => pc_target_2_11_port, ZN => n1064);
   U1522 : INV_X1 port map( A => n1065, ZN => n6440);
   U1523 : AOI22_X1 port map( A1 => Set_target(13), A2 => n1042, B1 => n1043, 
                           B2 => pc_target_2_13_port, ZN => n1065);
   U1524 : INV_X1 port map( A => n1066, ZN => n6441);
   U1525 : AOI22_X1 port map( A1 => Set_target(15), A2 => n1042, B1 => n1043, 
                           B2 => pc_target_2_15_port, ZN => n1066);
   U1526 : INV_X1 port map( A => n1067, ZN => n6442);
   U1527 : AOI22_X1 port map( A1 => Set_target(17), A2 => n1042, B1 => n1043, 
                           B2 => pc_target_2_17_port, ZN => n1067);
   U1528 : INV_X1 port map( A => n1068, ZN => n6443);
   U1529 : AOI22_X1 port map( A1 => Set_target(19), A2 => n1042, B1 => n1043, 
                           B2 => pc_target_2_19_port, ZN => n1068);
   U1530 : INV_X1 port map( A => n1069, ZN => n6444);
   U1531 : AOI22_X1 port map( A1 => Set_target(21), A2 => n1042, B1 => n1043, 
                           B2 => pc_target_2_21_port, ZN => n1069);
   U1532 : INV_X1 port map( A => n1070, ZN => n6445);
   U1533 : AOI22_X1 port map( A1 => Set_target(23), A2 => n1042, B1 => n1043, 
                           B2 => pc_target_2_23_port, ZN => n1070);
   U1534 : INV_X1 port map( A => n1071, ZN => n6446);
   U1535 : AOI22_X1 port map( A1 => Set_target(25), A2 => n1042, B1 => n1043, 
                           B2 => pc_target_2_25_port, ZN => n1071);
   U1536 : INV_X1 port map( A => n1072, ZN => n6447);
   U1537 : AOI22_X1 port map( A1 => Set_target(27), A2 => n1042, B1 => n1043, 
                           B2 => pc_target_2_27_port, ZN => n1072);
   U1538 : INV_X1 port map( A => n1073, ZN => n6448);
   U1539 : AOI22_X1 port map( A1 => Set_target(29), A2 => n1042, B1 => n1043, 
                           B2 => pc_target_2_29_port, ZN => n1073);
   U1540 : INV_X1 port map( A => n1074, ZN => n6449);
   U1541 : AOI22_X1 port map( A1 => Set_target(31), A2 => n1042, B1 => n1043, 
                           B2 => pc_target_2_31_port, ZN => n1074);
   U1544 : OAI22_X1 port map( A1 => n75, A2 => n1075, B1 => n1076, B2 => n1077,
                           ZN => n6450);
   U1545 : OAI22_X1 port map( A1 => n79, A2 => n1075, B1 => n1076, B2 => n1078,
                           ZN => n6451);
   U1546 : OAI22_X1 port map( A1 => n81, A2 => n1075, B1 => n1076, B2 => n1079,
                           ZN => n6452);
   U1547 : OAI22_X1 port map( A1 => n83, A2 => n1075, B1 => n1076, B2 => n1080,
                           ZN => n6453);
   U1548 : OAI22_X1 port map( A1 => n85, A2 => n1075, B1 => n1076, B2 => n1081,
                           ZN => n6454);
   U1549 : OAI22_X1 port map( A1 => n87, A2 => n1075, B1 => n1076, B2 => n1082,
                           ZN => n6455);
   U1550 : OAI22_X1 port map( A1 => n89, A2 => n1075, B1 => n1076, B2 => n1083,
                           ZN => n6456);
   U1551 : OAI22_X1 port map( A1 => n91, A2 => n1075, B1 => n1076, B2 => n1084,
                           ZN => n6457);
   U1552 : OAI22_X1 port map( A1 => n93, A2 => n1075, B1 => n1076, B2 => n1085,
                           ZN => n6458);
   U1553 : OAI22_X1 port map( A1 => n95, A2 => n1075, B1 => n1076, B2 => n1086,
                           ZN => n6459);
   U1554 : OAI22_X1 port map( A1 => n97_port, A2 => n1075, B1 => n1076, B2 => 
                           n1087, ZN => n6460);
   U1555 : OAI22_X1 port map( A1 => n99_port, A2 => n1075, B1 => n1076, B2 => 
                           n1088, ZN => n6461);
   U1556 : OAI22_X1 port map( A1 => n101_port, A2 => n1075, B1 => n1076, B2 => 
                           n1089, ZN => n6462);
   U1557 : OAI22_X1 port map( A1 => n103_port, A2 => n1075, B1 => n1076, B2 => 
                           n1090, ZN => n6463);
   U1558 : OAI22_X1 port map( A1 => n105_port, A2 => n1075, B1 => n1076, B2 => 
                           n1091, ZN => n6464);
   U1559 : OAI22_X1 port map( A1 => n107_port, A2 => n1075, B1 => n1076, B2 => 
                           n1092, ZN => n6465);
   U1560 : OAI22_X1 port map( A1 => n109_port, A2 => n1075, B1 => n1076, B2 => 
                           n1093, ZN => n6466);
   U1561 : OAI22_X1 port map( A1 => n111_port, A2 => n1075, B1 => n1076, B2 => 
                           n1094, ZN => n6467);
   U1562 : OAI22_X1 port map( A1 => n113_port, A2 => n1075, B1 => n1076, B2 => 
                           n1095, ZN => n6468);
   U1563 : OAI22_X1 port map( A1 => n115_port, A2 => n1075, B1 => n1076, B2 => 
                           n1096, ZN => n6469);
   U1564 : OAI22_X1 port map( A1 => n117_port, A2 => n1075, B1 => n1076, B2 => 
                           n1097, ZN => n6470);
   U1565 : OAI22_X1 port map( A1 => n119_port, A2 => n1075, B1 => n1076, B2 => 
                           n1098, ZN => n6471);
   U1566 : OAI22_X1 port map( A1 => n121_port, A2 => n1075, B1 => n1076, B2 => 
                           n1099, ZN => n6472);
   U1567 : OAI22_X1 port map( A1 => n123_port, A2 => n1075, B1 => n1076, B2 => 
                           n1100, ZN => n6473);
   U1568 : OAI22_X1 port map( A1 => n125_port, A2 => n1075, B1 => n1076, B2 => 
                           n1101, ZN => n6474);
   U1569 : OAI22_X1 port map( A1 => n127_port, A2 => n1075, B1 => n1076, B2 => 
                           n1102, ZN => n6475);
   U1570 : OAI22_X1 port map( A1 => n129, A2 => n1075, B1 => n1076, B2 => n1103
                           , ZN => n6476);
   U1571 : OAI22_X1 port map( A1 => n131, A2 => n1075, B1 => n1076, B2 => n1104
                           , ZN => n6477);
   U1572 : OAI22_X1 port map( A1 => n133, A2 => n1075, B1 => n1076, B2 => n1105
                           , ZN => n6478);
   U1573 : OAI22_X1 port map( A1 => n135, A2 => n1075, B1 => n1076, B2 => n1106
                           , ZN => n6479);
   U1574 : OAI22_X1 port map( A1 => n137, A2 => n1075, B1 => n1076, B2 => n1107
                           , ZN => n6480);
   U1575 : OAI22_X1 port map( A1 => n139, A2 => n1075, B1 => n1076, B2 => n1108
                           , ZN => n6481);
   U1578 : OAI22_X1 port map( A1 => n75, A2 => n1109, B1 => n1110, B2 => n1111,
                           ZN => n6482);
   U1580 : OAI22_X1 port map( A1 => n79, A2 => n1109, B1 => n1110, B2 => n1112,
                           ZN => n6483);
   U1582 : OAI22_X1 port map( A1 => n81, A2 => n1109, B1 => n1110, B2 => n1113,
                           ZN => n6484);
   U1584 : OAI22_X1 port map( A1 => n83, A2 => n1109, B1 => n1110, B2 => n1114,
                           ZN => n6485);
   U1586 : OAI22_X1 port map( A1 => n85, A2 => n1109, B1 => n1110, B2 => n1115,
                           ZN => n6486);
   U1588 : OAI22_X1 port map( A1 => n87, A2 => n1109, B1 => n1110, B2 => n1116,
                           ZN => n6487);
   U1590 : OAI22_X1 port map( A1 => n89, A2 => n1109, B1 => n1110, B2 => n1117,
                           ZN => n6488);
   U1592 : OAI22_X1 port map( A1 => n91, A2 => n1109, B1 => n1110, B2 => n1118,
                           ZN => n6489);
   U1594 : OAI22_X1 port map( A1 => n93, A2 => n1109, B1 => n1110, B2 => n1119,
                           ZN => n6490);
   U1596 : OAI22_X1 port map( A1 => n95, A2 => n1109, B1 => n1110, B2 => n1120,
                           ZN => n6491);
   U1598 : OAI22_X1 port map( A1 => n97_port, A2 => n1109, B1 => n1110, B2 => 
                           n1121, ZN => n6492);
   U1599 : INV_X1 port map( A => Set_target(10), ZN => n97_port);
   U1600 : OAI22_X1 port map( A1 => n99_port, A2 => n1109, B1 => n1110, B2 => 
                           n1122, ZN => n6493);
   U1601 : INV_X1 port map( A => Set_target(8), ZN => n99_port);
   U1602 : OAI22_X1 port map( A1 => n101_port, A2 => n1109, B1 => n1110, B2 => 
                           n1123, ZN => n6494);
   U1603 : INV_X1 port map( A => Set_target(6), ZN => n101_port);
   U1604 : OAI22_X1 port map( A1 => n103_port, A2 => n1109, B1 => n1110, B2 => 
                           n1124, ZN => n6495);
   U1605 : INV_X1 port map( A => Set_target(4), ZN => n103_port);
   U1606 : OAI22_X1 port map( A1 => n105_port, A2 => n1109, B1 => n1110, B2 => 
                           n1125, ZN => n6496);
   U1607 : INV_X1 port map( A => Set_target(2), ZN => n105_port);
   U1608 : OAI22_X1 port map( A1 => n107_port, A2 => n1109, B1 => n1110, B2 => 
                           n1126, ZN => n6497);
   U1609 : INV_X1 port map( A => Set_target(0), ZN => n107_port);
   U1610 : OAI22_X1 port map( A1 => n109_port, A2 => n1109, B1 => n1110, B2 => 
                           n1127, ZN => n6498);
   U1611 : INV_X1 port map( A => Set_target(1), ZN => n109_port);
   U1612 : OAI22_X1 port map( A1 => n111_port, A2 => n1109, B1 => n1110, B2 => 
                           n1128, ZN => n6499);
   U1613 : INV_X1 port map( A => Set_target(3), ZN => n111_port);
   U1614 : OAI22_X1 port map( A1 => n113_port, A2 => n1109, B1 => n1110, B2 => 
                           n1129, ZN => n6500);
   U1615 : INV_X1 port map( A => Set_target(5), ZN => n113_port);
   U1616 : OAI22_X1 port map( A1 => n115_port, A2 => n1109, B1 => n1110, B2 => 
                           n1130, ZN => n6501);
   U1617 : INV_X1 port map( A => Set_target(7), ZN => n115_port);
   U1618 : OAI22_X1 port map( A1 => n117_port, A2 => n1109, B1 => n1110, B2 => 
                           n1131, ZN => n6502);
   U1619 : INV_X1 port map( A => Set_target(9), ZN => n117_port);
   U1620 : OAI22_X1 port map( A1 => n119_port, A2 => n1109, B1 => n1110, B2 => 
                           n1132, ZN => n6503);
   U1622 : OAI22_X1 port map( A1 => n121_port, A2 => n1109, B1 => n1110, B2 => 
                           n1133, ZN => n6504);
   U1624 : OAI22_X1 port map( A1 => n123_port, A2 => n1109, B1 => n1110, B2 => 
                           n1134, ZN => n6505);
   U1626 : OAI22_X1 port map( A1 => n125_port, A2 => n1109, B1 => n1110, B2 => 
                           n1135, ZN => n6506);
   U1628 : OAI22_X1 port map( A1 => n127_port, A2 => n1109, B1 => n1110, B2 => 
                           n1136, ZN => n6507);
   U1630 : OAI22_X1 port map( A1 => n129, A2 => n1109, B1 => n1110, B2 => n1137
                           , ZN => n6508);
   U1632 : OAI22_X1 port map( A1 => n131, A2 => n1109, B1 => n1110, B2 => n1138
                           , ZN => n6509);
   U1634 : OAI22_X1 port map( A1 => n133, A2 => n1109, B1 => n1110, B2 => n1139
                           , ZN => n6510);
   U1636 : OAI22_X1 port map( A1 => n135, A2 => n1109, B1 => n1110, B2 => n1140
                           , ZN => n6511);
   U1638 : OAI22_X1 port map( A1 => n137, A2 => n1109, B1 => n1110, B2 => n1141
                           , ZN => n6512);
   U1640 : OAI22_X1 port map( A1 => n139, A2 => n1109, B1 => n1110, B2 => n1142
                           , ZN => n6513);
   U1646 : INV_X1 port map( A => Set_target(31), ZN => n139);
   U1647 : OAI22_X1 port map( A1 => n3808, A2 => n1146, B1 => n1147, B2 => 
                           n1148, ZN => n6514);
   U1649 : OAI22_X1 port map( A1 => n3808, A2 => n1149, B1 => n1148, B2 => 
                           n1150, ZN => n6515);
   U1651 : OAI22_X1 port map( A1 => n3809, A2 => n1151, B1 => n1148, B2 => 
                           n1152, ZN => n6516);
   U1653 : OAI22_X1 port map( A1 => n3809, A2 => n1153, B1 => n1148, B2 => 
                           n1154, ZN => n6517);
   U1655 : OAI22_X1 port map( A1 => n3808, A2 => n1155, B1 => n1148, B2 => 
                           n1156, ZN => n6518);
   U1657 : OAI22_X1 port map( A1 => n3808, A2 => n1157, B1 => n1148, B2 => 
                           n1158, ZN => n6519);
   U1659 : OAI22_X1 port map( A1 => n3809, A2 => n1159, B1 => n1148, B2 => 
                           n1160, ZN => n6520);
   U1661 : OAI22_X1 port map( A1 => n3809, A2 => n1161, B1 => n1148, B2 => 
                           n1162, ZN => n6521);
   U1663 : OAI22_X1 port map( A1 => n3809, A2 => n1163, B1 => n1148, B2 => 
                           n1164, ZN => n6522);
   U1665 : OAI22_X1 port map( A1 => n3808, A2 => n1165, B1 => n1148, B2 => 
                           n1166, ZN => n6523);
   U1667 : OAI22_X1 port map( A1 => n3809, A2 => n1167, B1 => n1148, B2 => 
                           n1168, ZN => n6524);
   U1669 : OAI22_X1 port map( A1 => n3809, A2 => n1169, B1 => n1148, B2 => 
                           n1170, ZN => n6525);
   U1671 : OAI22_X1 port map( A1 => n3809, A2 => n1171, B1 => n1148, B2 => 
                           n1172, ZN => n6526);
   U1673 : INV_X1 port map( A => n1173, ZN => n6527);
   U1674 : AOI22_X1 port map( A1 => n1148, A2 => pc_lut_31_4_port, B1 => n3521,
                           B2 => n3809, ZN => n1173);
   U1675 : INV_X1 port map( A => n1174, ZN => n6528);
   U1676 : AOI22_X1 port map( A1 => n1148, A2 => pc_lut_31_2_port, B1 => n3521,
                           B2 => n3807, ZN => n1174);
   U1677 : INV_X1 port map( A => n1175, ZN => n6529);
   U1678 : AOI22_X1 port map( A1 => n1148, A2 => pc_lut_31_0_port, B1 => n3521,
                           B2 => n3807, ZN => n1175);
   U1679 : INV_X1 port map( A => n1176, ZN => n6530);
   U1680 : AOI22_X1 port map( A1 => n1148, A2 => pc_lut_31_1_port, B1 => n3521,
                           B2 => n3807, ZN => n1176);
   U1681 : INV_X1 port map( A => n1177, ZN => n6531);
   U1682 : AOI22_X1 port map( A1 => n1148, A2 => pc_lut_31_3_port, B1 => n3521,
                           B2 => n3807, ZN => n1177);
   U1683 : OAI22_X1 port map( A1 => n3808, A2 => n1178, B1 => n1148, B2 => 
                           n1179, ZN => n6532);
   U1685 : OAI22_X1 port map( A1 => n3809, A2 => n1180, B1 => n1148, B2 => 
                           n1181, ZN => n6533);
   U1687 : OAI22_X1 port map( A1 => n3809, A2 => n1182, B1 => n1148, B2 => 
                           n1183, ZN => n6534);
   U1689 : OAI22_X1 port map( A1 => n3808, A2 => n1184, B1 => n1148, B2 => 
                           n1185, ZN => n6535);
   U1691 : OAI22_X1 port map( A1 => n3809, A2 => n1186, B1 => n1148, B2 => 
                           n1187, ZN => n6536);
   U1693 : OAI22_X1 port map( A1 => n3808, A2 => n1188, B1 => n1148, B2 => 
                           n1189, ZN => n6537);
   U1695 : OAI22_X1 port map( A1 => n3809, A2 => n1190, B1 => n1148, B2 => 
                           n1191, ZN => n6538);
   U1697 : OAI22_X1 port map( A1 => n3808, A2 => n1192, B1 => n1148, B2 => 
                           n1193, ZN => n6539);
   U1699 : OAI22_X1 port map( A1 => n3809, A2 => n1194, B1 => n1148, B2 => 
                           n1195, ZN => n6540);
   U1701 : OAI22_X1 port map( A1 => n3808, A2 => n1196, B1 => n1148, B2 => 
                           n1197, ZN => n6541);
   U1703 : OAI22_X1 port map( A1 => n3808, A2 => n1198, B1 => n1148, B2 => 
                           n1199, ZN => n6542);
   U1705 : OAI22_X1 port map( A1 => n3808, A2 => n1200, B1 => n1148, B2 => 
                           n1201, ZN => n6543);
   U1707 : OAI22_X1 port map( A1 => n3808, A2 => n1202, B1 => n1148, B2 => 
                           n1203, ZN => n6544);
   U1709 : OAI22_X1 port map( A1 => n3808, A2 => n1204, B1 => n1148, B2 => 
                           n1205, ZN => n6545);
   U1713 : OAI22_X1 port map( A1 => n3805, A2 => n1208, B1 => n1147, B2 => 
                           n1209, ZN => n6546);
   U1715 : OAI22_X1 port map( A1 => n3805, A2 => n1210, B1 => n1150, B2 => 
                           n1209, ZN => n6547);
   U1717 : OAI22_X1 port map( A1 => n3805, A2 => n1211, B1 => n1152, B2 => 
                           n1209, ZN => n6548);
   U1719 : OAI22_X1 port map( A1 => n3805, A2 => n1212, B1 => n1154, B2 => 
                           n1209, ZN => n6549);
   U1721 : OAI22_X1 port map( A1 => n3805, A2 => n1213, B1 => n1156, B2 => 
                           n1209, ZN => n6550);
   U1723 : OAI22_X1 port map( A1 => n3805, A2 => n1214, B1 => n1158, B2 => 
                           n1209, ZN => n6551);
   U1725 : OAI22_X1 port map( A1 => n3805, A2 => n1215, B1 => n1160, B2 => 
                           n1209, ZN => n6552);
   U1727 : OAI22_X1 port map( A1 => n3805, A2 => n1216, B1 => n1162, B2 => 
                           n1209, ZN => n6553);
   U1729 : OAI22_X1 port map( A1 => n3805, A2 => n1217, B1 => n1164, B2 => 
                           n1209, ZN => n6554);
   U1731 : OAI22_X1 port map( A1 => n3805, A2 => n1218, B1 => n1166, B2 => 
                           n1209, ZN => n6555);
   U1733 : OAI22_X1 port map( A1 => n3805, A2 => n1219, B1 => n1168, B2 => 
                           n1209, ZN => n6556);
   U1735 : OAI22_X1 port map( A1 => n3805, A2 => n1220, B1 => n1170, B2 => 
                           n1209, ZN => n6557);
   U1737 : OAI22_X1 port map( A1 => n3805, A2 => n1221, B1 => n1172, B2 => 
                           n1209, ZN => n6558);
   U1739 : INV_X1 port map( A => n1222, ZN => n6559);
   U1740 : AOI22_X1 port map( A1 => n1209, A2 => pc_lut_30_4_port, B1 => n3521,
                           B2 => n3805, ZN => n1222);
   U1741 : INV_X1 port map( A => n1223, ZN => n6560);
   U1742 : AOI22_X1 port map( A1 => n1209, A2 => pc_lut_30_2_port, B1 => n3521,
                           B2 => n3805, ZN => n1223);
   U1744 : INV_X1 port map( A => n1224, ZN => n6562);
   U1745 : AOI22_X1 port map( A1 => n1209, A2 => pc_lut_30_1_port, B1 => n3521,
                           B2 => n3805, ZN => n1224);
   U1746 : INV_X1 port map( A => n1225, ZN => n6563);
   U1747 : AOI22_X1 port map( A1 => n1209, A2 => pc_lut_30_3_port, B1 => n3521,
                           B2 => n3805, ZN => n1225);
   U1748 : OAI22_X1 port map( A1 => n3805, A2 => n1226, B1 => n1179, B2 => 
                           n1209, ZN => n6564);
   U1750 : OAI22_X1 port map( A1 => n3805, A2 => n1227, B1 => n1181, B2 => 
                           n1209, ZN => n6565);
   U1752 : OAI22_X1 port map( A1 => n3805, A2 => n1228, B1 => n1183, B2 => 
                           n1209, ZN => n6566);
   U1754 : OAI22_X1 port map( A1 => n3805, A2 => n1229, B1 => n1185, B2 => 
                           n1209, ZN => n6567);
   U1756 : OAI22_X1 port map( A1 => n3805, A2 => n1230, B1 => n1187, B2 => 
                           n1209, ZN => n6568);
   U1758 : OAI22_X1 port map( A1 => n3805, A2 => n1231, B1 => n1189, B2 => 
                           n1209, ZN => n6569);
   U1760 : OAI22_X1 port map( A1 => n3805, A2 => n1232, B1 => n1191, B2 => 
                           n1209, ZN => n6570);
   U1762 : OAI22_X1 port map( A1 => n3805, A2 => n1233, B1 => n1193, B2 => 
                           n1209, ZN => n6571);
   U1764 : OAI22_X1 port map( A1 => n3805, A2 => n1234, B1 => n1195, B2 => 
                           n1209, ZN => n6572);
   U1766 : OAI22_X1 port map( A1 => n3805, A2 => n1235, B1 => n1197, B2 => 
                           n1209, ZN => n6573);
   U1768 : OAI22_X1 port map( A1 => n3805, A2 => n1236, B1 => n1199, B2 => 
                           n1209, ZN => n6574);
   U1770 : OAI22_X1 port map( A1 => n3805, A2 => n1237, B1 => n1201, B2 => 
                           n1209, ZN => n6575);
   U1772 : OAI22_X1 port map( A1 => n3805, A2 => n1238, B1 => n1203, B2 => 
                           n1209, ZN => n6576);
   U1774 : OAI22_X1 port map( A1 => n3805, A2 => n1239, B1 => n1205, B2 => 
                           n1209, ZN => n6577);
   U1778 : OAI22_X1 port map( A1 => n3536, A2 => n1241, B1 => n1147, B2 => 
                           n1242, ZN => n6578);
   U1779 : OAI22_X1 port map( A1 => n3536, A2 => n1243, B1 => n1150, B2 => 
                           n1242, ZN => n6579);
   U1780 : OAI22_X1 port map( A1 => n3536, A2 => n1244, B1 => n1152, B2 => 
                           n1242, ZN => n6580);
   U1781 : OAI22_X1 port map( A1 => n3536, A2 => n1245, B1 => n1154, B2 => 
                           n1242, ZN => n6581);
   U1782 : OAI22_X1 port map( A1 => n3536, A2 => n1246, B1 => n1156, B2 => 
                           n1242, ZN => n6582);
   U1783 : OAI22_X1 port map( A1 => n3536, A2 => n1247, B1 => n1158, B2 => 
                           n1242, ZN => n6583);
   U1784 : OAI22_X1 port map( A1 => n3536, A2 => n1248, B1 => n1160, B2 => 
                           n1242, ZN => n6584);
   U1785 : OAI22_X1 port map( A1 => n3536, A2 => n1249, B1 => n1162, B2 => 
                           n1242, ZN => n6585);
   U1786 : OAI22_X1 port map( A1 => n3536, A2 => n1250, B1 => n1164, B2 => 
                           n1242, ZN => n6586);
   U1787 : OAI22_X1 port map( A1 => n3536, A2 => n1251, B1 => n1166, B2 => 
                           n1242, ZN => n6587);
   U1788 : OAI22_X1 port map( A1 => n3536, A2 => n1252, B1 => n1168, B2 => 
                           n1242, ZN => n6588);
   U1789 : OAI22_X1 port map( A1 => n3536, A2 => n1253, B1 => n1170, B2 => 
                           n1242, ZN => n6589);
   U1790 : OAI22_X1 port map( A1 => n3536, A2 => n1254, B1 => n1172, B2 => 
                           n1242, ZN => n6590);
   U1791 : OAI22_X1 port map( A1 => n3536, A2 => n1255, B1 => n1496, B2 => 
                           n1242, ZN => n6591);
   U1792 : OAI22_X1 port map( A1 => n3536, A2 => n1257, B1 => n1496, B2 => 
                           n1242, ZN => n6592);
   U1793 : OAI22_X1 port map( A1 => n3536, A2 => n1258, B1 => n1496, B2 => 
                           n1242, ZN => n6593);
   U1795 : OAI22_X1 port map( A1 => n3536, A2 => n1260, B1 => n1496, B2 => 
                           n1242, ZN => n6595);
   U1796 : OAI22_X1 port map( A1 => n3536, A2 => n1261, B1 => n1179, B2 => 
                           n1242, ZN => n6596);
   U1797 : OAI22_X1 port map( A1 => n3536, A2 => n1262, B1 => n1181, B2 => 
                           n1242, ZN => n6597);
   U1798 : OAI22_X1 port map( A1 => n3536, A2 => n1263, B1 => n1183, B2 => 
                           n1242, ZN => n6598);
   U1799 : OAI22_X1 port map( A1 => n3536, A2 => n1264, B1 => n1185, B2 => 
                           n1242, ZN => n6599);
   U1800 : OAI22_X1 port map( A1 => n3536, A2 => n1265, B1 => n1187, B2 => 
                           n1242, ZN => n6600);
   U1801 : OAI22_X1 port map( A1 => n3536, A2 => n1266, B1 => n1189, B2 => 
                           n1242, ZN => n6601);
   U1802 : OAI22_X1 port map( A1 => n3536, A2 => n1267, B1 => n1191, B2 => 
                           n1242, ZN => n6602);
   U1803 : OAI22_X1 port map( A1 => n3536, A2 => n1268, B1 => n1193, B2 => 
                           n1242, ZN => n6603);
   U1804 : OAI22_X1 port map( A1 => n3536, A2 => n1269, B1 => n1195, B2 => 
                           n1242, ZN => n6604);
   U1805 : OAI22_X1 port map( A1 => n3536, A2 => n1270, B1 => n1197, B2 => 
                           n1242, ZN => n6605);
   U1806 : OAI22_X1 port map( A1 => n3536, A2 => n1271, B1 => n1199, B2 => 
                           n1242, ZN => n6606);
   U1807 : OAI22_X1 port map( A1 => n3536, A2 => n1272, B1 => n1201, B2 => 
                           n1242, ZN => n6607);
   U1808 : OAI22_X1 port map( A1 => n3536, A2 => n1273, B1 => n1203, B2 => 
                           n1242, ZN => n6608);
   U1809 : OAI22_X1 port map( A1 => n3536, A2 => n1274, B1 => n1205, B2 => 
                           n1242, ZN => n6609);
   U1812 : OAI22_X1 port map( A1 => n3534, A2 => n1276, B1 => n1147, B2 => 
                           n1277, ZN => n6610);
   U1813 : OAI22_X1 port map( A1 => n3534, A2 => n1278, B1 => n1150, B2 => 
                           n1277, ZN => n6611);
   U1814 : OAI22_X1 port map( A1 => n3534, A2 => n1279, B1 => n1152, B2 => 
                           n1277, ZN => n6612);
   U1815 : OAI22_X1 port map( A1 => n3534, A2 => n1280, B1 => n1154, B2 => 
                           n1277, ZN => n6613);
   U1816 : OAI22_X1 port map( A1 => n3534, A2 => n1281, B1 => n1156, B2 => 
                           n1277, ZN => n6614);
   U1817 : OAI22_X1 port map( A1 => n3534, A2 => n1282, B1 => n1158, B2 => 
                           n1277, ZN => n6615);
   U1818 : OAI22_X1 port map( A1 => n3534, A2 => n1283, B1 => n1160, B2 => 
                           n1277, ZN => n6616);
   U1819 : OAI22_X1 port map( A1 => n3534, A2 => n1284, B1 => n1162, B2 => 
                           n1277, ZN => n6617);
   U1820 : OAI22_X1 port map( A1 => n3534, A2 => n1285, B1 => n1164, B2 => 
                           n1277, ZN => n6618);
   U1821 : OAI22_X1 port map( A1 => n3534, A2 => n1286, B1 => n1166, B2 => 
                           n1277, ZN => n6619);
   U1822 : OAI22_X1 port map( A1 => n3534, A2 => n1287, B1 => n1168, B2 => 
                           n1277, ZN => n6620);
   U1823 : OAI22_X1 port map( A1 => n3534, A2 => n1288, B1 => n1170, B2 => 
                           n1277, ZN => n6621);
   U1824 : OAI22_X1 port map( A1 => n3534, A2 => n1289, B1 => n1172, B2 => 
                           n1277, ZN => n6622);
   U1825 : OAI22_X1 port map( A1 => n3534, A2 => n1290, B1 => n1496, B2 => 
                           n1277, ZN => n6623);
   U1826 : OAI22_X1 port map( A1 => n3534, A2 => n1291, B1 => n1496, B2 => 
                           n1277, ZN => n6624);
   U1829 : OAI22_X1 port map( A1 => n3534, A2 => n1294, B1 => n1496, B2 => 
                           n1277, ZN => n6627);
   U1830 : OAI22_X1 port map( A1 => n3534, A2 => n1295, B1 => n1179, B2 => 
                           n1277, ZN => n6628);
   U1831 : OAI22_X1 port map( A1 => n3534, A2 => n1296, B1 => n1181, B2 => 
                           n1277, ZN => n6629);
   U1832 : OAI22_X1 port map( A1 => n3534, A2 => n1297, B1 => n1183, B2 => 
                           n1277, ZN => n6630);
   U1833 : OAI22_X1 port map( A1 => n3534, A2 => n1298, B1 => n1185, B2 => 
                           n1277, ZN => n6631);
   U1834 : OAI22_X1 port map( A1 => n3534, A2 => n1299, B1 => n1187, B2 => 
                           n1277, ZN => n6632);
   U1835 : OAI22_X1 port map( A1 => n3534, A2 => n1300, B1 => n1189, B2 => 
                           n1277, ZN => n6633);
   U1836 : OAI22_X1 port map( A1 => n3534, A2 => n1301, B1 => n1191, B2 => 
                           n1277, ZN => n6634);
   U1837 : OAI22_X1 port map( A1 => n3534, A2 => n1302, B1 => n1193, B2 => 
                           n1277, ZN => n6635);
   U1838 : OAI22_X1 port map( A1 => n3534, A2 => n1303, B1 => n1195, B2 => 
                           n1277, ZN => n6636);
   U1839 : OAI22_X1 port map( A1 => n3534, A2 => n1304, B1 => n1197, B2 => 
                           n1277, ZN => n6637);
   U1840 : OAI22_X1 port map( A1 => n3534, A2 => n1305, B1 => n1199, B2 => 
                           n1277, ZN => n6638);
   U1841 : OAI22_X1 port map( A1 => n3534, A2 => n1306, B1 => n1201, B2 => 
                           n1277, ZN => n6639);
   U1842 : OAI22_X1 port map( A1 => n3534, A2 => n1307, B1 => n1203, B2 => 
                           n1277, ZN => n6640);
   U1843 : OAI22_X1 port map( A1 => n3534, A2 => n1308, B1 => n1205, B2 => 
                           n1277, ZN => n6641);
   U1847 : OAI22_X1 port map( A1 => n3803, A2 => n1311, B1 => n1147, B2 => 
                           n1312, ZN => n6642);
   U1849 : OAI22_X1 port map( A1 => n3803, A2 => n1313, B1 => n1150, B2 => 
                           n1312, ZN => n6643);
   U1851 : OAI22_X1 port map( A1 => n3804, A2 => n1314, B1 => n1152, B2 => 
                           n1312, ZN => n6644);
   U1853 : OAI22_X1 port map( A1 => n3804, A2 => n1315, B1 => n1154, B2 => 
                           n1312, ZN => n6645);
   U1855 : OAI22_X1 port map( A1 => n3803, A2 => n1316, B1 => n1156, B2 => 
                           n1312, ZN => n6646);
   U1857 : OAI22_X1 port map( A1 => n3803, A2 => n1317, B1 => n1158, B2 => 
                           n1312, ZN => n6647);
   U1859 : OAI22_X1 port map( A1 => n3804, A2 => n1318, B1 => n1160, B2 => 
                           n1312, ZN => n6648);
   U1861 : OAI22_X1 port map( A1 => n3803, A2 => n1319, B1 => n1162, B2 => 
                           n1312, ZN => n6649);
   U1863 : OAI22_X1 port map( A1 => n3804, A2 => n1320, B1 => n1164, B2 => 
                           n1312, ZN => n6650);
   U1865 : OAI22_X1 port map( A1 => n3804, A2 => n1321, B1 => n1166, B2 => 
                           n1312, ZN => n6651);
   U1867 : OAI22_X1 port map( A1 => n3804, A2 => n1322, B1 => n1168, B2 => 
                           n1312, ZN => n6652);
   U1869 : OAI22_X1 port map( A1 => n3804, A2 => n1323, B1 => n1170, B2 => 
                           n1312, ZN => n6653);
   U1871 : OAI22_X1 port map( A1 => n3803, A2 => n1324, B1 => n1172, B2 => 
                           n1312, ZN => n6654);
   U1873 : INV_X1 port map( A => n1325, ZN => n6655);
   U1874 : AOI22_X1 port map( A1 => n1312, A2 => pc_lut_27_4_port, B1 => n3521,
                           B2 => n3804, ZN => n1325);
   U1876 : INV_X1 port map( A => n1326, ZN => n6657);
   U1877 : AOI22_X1 port map( A1 => n1312, A2 => pc_lut_27_0_port, B1 => n3521,
                           B2 => n3802, ZN => n1326);
   U1878 : INV_X1 port map( A => n1327, ZN => n6658);
   U1879 : AOI22_X1 port map( A1 => n1312, A2 => pc_lut_27_1_port, B1 => n3521,
                           B2 => n3802, ZN => n1327);
   U1880 : INV_X1 port map( A => n1328, ZN => n6659);
   U1881 : AOI22_X1 port map( A1 => n1312, A2 => pc_lut_27_3_port, B1 => n3521,
                           B2 => n3802, ZN => n1328);
   U1882 : OAI22_X1 port map( A1 => n3803, A2 => n1329, B1 => n1179, B2 => 
                           n1312, ZN => n6660);
   U1884 : OAI22_X1 port map( A1 => n3803, A2 => n1330, B1 => n1181, B2 => 
                           n1312, ZN => n6661);
   U1886 : OAI22_X1 port map( A1 => n3804, A2 => n1331, B1 => n1183, B2 => 
                           n1312, ZN => n6662);
   U1888 : OAI22_X1 port map( A1 => n3803, A2 => n1332, B1 => n1185, B2 => 
                           n1312, ZN => n6663);
   U1890 : OAI22_X1 port map( A1 => n3804, A2 => n1333, B1 => n1187, B2 => 
                           n1312, ZN => n6664);
   U1892 : OAI22_X1 port map( A1 => n3803, A2 => n1334, B1 => n1189, B2 => 
                           n1312, ZN => n6665);
   U1894 : OAI22_X1 port map( A1 => n3804, A2 => n1335, B1 => n1191, B2 => 
                           n1312, ZN => n6666);
   U1896 : OAI22_X1 port map( A1 => n3803, A2 => n1336, B1 => n1193, B2 => 
                           n1312, ZN => n6667);
   U1898 : OAI22_X1 port map( A1 => n3804, A2 => n1337, B1 => n1195, B2 => 
                           n1312, ZN => n6668);
   U1900 : OAI22_X1 port map( A1 => n3803, A2 => n1338, B1 => n1197, B2 => 
                           n1312, ZN => n6669);
   U1902 : OAI22_X1 port map( A1 => n3804, A2 => n1339, B1 => n1199, B2 => 
                           n1312, ZN => n6670);
   U1904 : OAI22_X1 port map( A1 => n3803, A2 => n1340, B1 => n1201, B2 => 
                           n1312, ZN => n6671);
   U1906 : OAI22_X1 port map( A1 => n3804, A2 => n1341, B1 => n1203, B2 => 
                           n1312, ZN => n6672);
   U1908 : OAI22_X1 port map( A1 => n3803, A2 => n1342, B1 => n1205, B2 => 
                           n1312, ZN => n6673);
   U1912 : OAI22_X1 port map( A1 => n3538, A2 => n1345, B1 => n1147, B2 => 
                           n1346, ZN => n6674);
   U1914 : OAI22_X1 port map( A1 => n3538, A2 => n1347, B1 => n1150, B2 => 
                           n1346, ZN => n6675);
   U1916 : OAI22_X1 port map( A1 => n3538, A2 => n1348, B1 => n1152, B2 => 
                           n1346, ZN => n6676);
   U1918 : OAI22_X1 port map( A1 => n3538, A2 => n1349, B1 => n1154, B2 => 
                           n1346, ZN => n6677);
   U1920 : OAI22_X1 port map( A1 => n3538, A2 => n1350, B1 => n1156, B2 => 
                           n1346, ZN => n6678);
   U1922 : OAI22_X1 port map( A1 => n3538, A2 => n1351, B1 => n1158, B2 => 
                           n1346, ZN => n6679);
   U1924 : OAI22_X1 port map( A1 => n3538, A2 => n1352, B1 => n1160, B2 => 
                           n1346, ZN => n6680);
   U1926 : OAI22_X1 port map( A1 => n3538, A2 => n1353, B1 => n1162, B2 => 
                           n1346, ZN => n6681);
   U1928 : OAI22_X1 port map( A1 => n3538, A2 => n1354, B1 => n1164, B2 => 
                           n1346, ZN => n6682);
   U1930 : OAI22_X1 port map( A1 => n3538, A2 => n1355, B1 => n1166, B2 => 
                           n1346, ZN => n6683);
   U1932 : OAI22_X1 port map( A1 => n3538, A2 => n1356, B1 => n1168, B2 => 
                           n1346, ZN => n6684);
   U1934 : OAI22_X1 port map( A1 => n3538, A2 => n1357, B1 => n1170, B2 => 
                           n1346, ZN => n6685);
   U1936 : OAI22_X1 port map( A1 => n3538, A2 => n1358, B1 => n1172, B2 => 
                           n1346, ZN => n6686);
   U1938 : INV_X1 port map( A => n1359, ZN => n6687);
   U1939 : AOI22_X1 port map( A1 => n1346, A2 => pc_lut_26_4_port, B1 => n3521,
                           B2 => n3538, ZN => n1359);
   U1942 : INV_X1 port map( A => n1360, ZN => n6690);
   U1943 : AOI22_X1 port map( A1 => n1346, A2 => pc_lut_26_1_port, B1 => n3521,
                           B2 => n3538, ZN => n1360);
   U1944 : INV_X1 port map( A => n1361, ZN => n6691);
   U1945 : AOI22_X1 port map( A1 => n1346, A2 => pc_lut_26_3_port, B1 => n3521,
                           B2 => n3538, ZN => n1361);
   U1946 : OAI22_X1 port map( A1 => n3538, A2 => n1362, B1 => n1179, B2 => 
                           n1346, ZN => n6692);
   U1948 : OAI22_X1 port map( A1 => n3538, A2 => n1363, B1 => n1181, B2 => 
                           n1346, ZN => n6693);
   U1950 : OAI22_X1 port map( A1 => n3538, A2 => n1364, B1 => n1183, B2 => 
                           n1346, ZN => n6694);
   U1952 : OAI22_X1 port map( A1 => n3538, A2 => n1365, B1 => n1185, B2 => 
                           n1346, ZN => n6695);
   U1954 : OAI22_X1 port map( A1 => n3538, A2 => n1366, B1 => n1187, B2 => 
                           n1346, ZN => n6696);
   U1956 : OAI22_X1 port map( A1 => n3538, A2 => n1367, B1 => n1189, B2 => 
                           n1346, ZN => n6697);
   U1958 : OAI22_X1 port map( A1 => n3538, A2 => n1368, B1 => n1191, B2 => 
                           n1346, ZN => n6698);
   U1960 : OAI22_X1 port map( A1 => n3538, A2 => n1369, B1 => n1193, B2 => 
                           n1346, ZN => n6699);
   U1962 : OAI22_X1 port map( A1 => n3538, A2 => n1370, B1 => n1195, B2 => 
                           n1346, ZN => n6700);
   U1964 : OAI22_X1 port map( A1 => n3538, A2 => n1371, B1 => n1197, B2 => 
                           n1346, ZN => n6701);
   U1966 : OAI22_X1 port map( A1 => n3538, A2 => n1372, B1 => n1199, B2 => 
                           n1346, ZN => n6702);
   U1968 : OAI22_X1 port map( A1 => n3538, A2 => n1373, B1 => n1201, B2 => 
                           n1346, ZN => n6703);
   U1970 : OAI22_X1 port map( A1 => n3538, A2 => n1374, B1 => n1203, B2 => 
                           n1346, ZN => n6704);
   U1972 : OAI22_X1 port map( A1 => n3538, A2 => n1375, B1 => n1205, B2 => 
                           n1346, ZN => n6705);
   U1976 : OAI22_X1 port map( A1 => n1376, A2 => n1377, B1 => n1147, B2 => 
                           n1378, ZN => n6706);
   U1977 : OAI22_X1 port map( A1 => n1376, A2 => n1379, B1 => n1150, B2 => 
                           n1378, ZN => n6707);
   U1978 : OAI22_X1 port map( A1 => n1376, A2 => n1380, B1 => n1152, B2 => 
                           n1378, ZN => n6708);
   U1979 : OAI22_X1 port map( A1 => n1376, A2 => n1381, B1 => n1154, B2 => 
                           n1378, ZN => n6709);
   U1980 : OAI22_X1 port map( A1 => n1376, A2 => n1382, B1 => n1156, B2 => 
                           n1378, ZN => n6710);
   U1981 : OAI22_X1 port map( A1 => n1376, A2 => n1383, B1 => n1158, B2 => 
                           n1378, ZN => n6711);
   U1982 : OAI22_X1 port map( A1 => n1376, A2 => n1384, B1 => n1160, B2 => 
                           n1378, ZN => n6712);
   U1983 : OAI22_X1 port map( A1 => n1376, A2 => n1385, B1 => n1162, B2 => 
                           n1378, ZN => n6713);
   U1984 : OAI22_X1 port map( A1 => n1376, A2 => n1386, B1 => n1164, B2 => 
                           n1378, ZN => n6714);
   U1985 : OAI22_X1 port map( A1 => n1376, A2 => n1387, B1 => n1166, B2 => 
                           n1378, ZN => n6715);
   U1986 : OAI22_X1 port map( A1 => n1376, A2 => n1388, B1 => n1168, B2 => 
                           n1378, ZN => n6716);
   U1987 : OAI22_X1 port map( A1 => n1376, A2 => n1389, B1 => n1170, B2 => 
                           n1378, ZN => n6717);
   U1988 : OAI22_X1 port map( A1 => n1376, A2 => n1390, B1 => n1172, B2 => 
                           n1378, ZN => n6718);
   U1989 : OAI22_X1 port map( A1 => n1376, A2 => n1391, B1 => n3529, B2 => 
                           n1378, ZN => n6719);
   U1991 : OAI22_X1 port map( A1 => n1376, A2 => n1393, B1 => n3529, B2 => 
                           n1378, ZN => n6721);
   U1993 : OAI22_X1 port map( A1 => n1376, A2 => n1395, B1 => n3529, B2 => 
                           n1378, ZN => n6723);
   U1994 : OAI22_X1 port map( A1 => n1376, A2 => n1396, B1 => n1179, B2 => 
                           n1378, ZN => n6724);
   U1995 : OAI22_X1 port map( A1 => n1376, A2 => n1397, B1 => n1181, B2 => 
                           n1378, ZN => n6725);
   U1996 : OAI22_X1 port map( A1 => n1376, A2 => n1398, B1 => n1183, B2 => 
                           n1378, ZN => n6726);
   U1997 : OAI22_X1 port map( A1 => n1376, A2 => n1399, B1 => n1185, B2 => 
                           n1378, ZN => n6727);
   U1998 : OAI22_X1 port map( A1 => n1376, A2 => n1400, B1 => n1187, B2 => 
                           n1378, ZN => n6728);
   U1999 : OAI22_X1 port map( A1 => n1376, A2 => n1401, B1 => n1189, B2 => 
                           n1378, ZN => n6729);
   U2000 : OAI22_X1 port map( A1 => n1376, A2 => n1402, B1 => n1191, B2 => 
                           n1378, ZN => n6730);
   U2001 : OAI22_X1 port map( A1 => n1376, A2 => n1403, B1 => n1193, B2 => 
                           n1378, ZN => n6731);
   U2002 : OAI22_X1 port map( A1 => n1376, A2 => n1404, B1 => n1195, B2 => 
                           n1378, ZN => n6732);
   U2003 : OAI22_X1 port map( A1 => n1376, A2 => n1405, B1 => n1197, B2 => 
                           n1378, ZN => n6733);
   U2004 : OAI22_X1 port map( A1 => n1376, A2 => n1406, B1 => n1199, B2 => 
                           n1378, ZN => n6734);
   U2005 : OAI22_X1 port map( A1 => n1376, A2 => n1407, B1 => n1201, B2 => 
                           n1378, ZN => n6735);
   U2006 : OAI22_X1 port map( A1 => n1376, A2 => n1408, B1 => n1203, B2 => 
                           n1378, ZN => n6736);
   U2007 : OAI22_X1 port map( A1 => n1376, A2 => n1409, B1 => n1205, B2 => 
                           n1378, ZN => n6737);
   U2010 : OAI22_X1 port map( A1 => n1410, A2 => n1411, B1 => n1147, B2 => 
                           n1412, ZN => n6738);
   U2011 : OAI22_X1 port map( A1 => n1410, A2 => n1413, B1 => n1150, B2 => 
                           n1412, ZN => n6739);
   U2012 : OAI22_X1 port map( A1 => n1410, A2 => n1414, B1 => n1152, B2 => 
                           n1412, ZN => n6740);
   U2013 : OAI22_X1 port map( A1 => n1410, A2 => n1415, B1 => n1154, B2 => 
                           n1412, ZN => n6741);
   U2014 : OAI22_X1 port map( A1 => n1410, A2 => n1416, B1 => n1156, B2 => 
                           n1412, ZN => n6742);
   U2015 : OAI22_X1 port map( A1 => n1410, A2 => n1417, B1 => n1158, B2 => 
                           n1412, ZN => n6743);
   U2016 : OAI22_X1 port map( A1 => n1410, A2 => n1418, B1 => n1160, B2 => 
                           n1412, ZN => n6744);
   U2017 : OAI22_X1 port map( A1 => n1410, A2 => n1419, B1 => n1162, B2 => 
                           n1412, ZN => n6745);
   U2018 : OAI22_X1 port map( A1 => n1410, A2 => n1420, B1 => n1164, B2 => 
                           n1412, ZN => n6746);
   U2019 : OAI22_X1 port map( A1 => n1410, A2 => n1421, B1 => n1166, B2 => 
                           n1412, ZN => n6747);
   U2020 : OAI22_X1 port map( A1 => n1410, A2 => n1422, B1 => n1168, B2 => 
                           n1412, ZN => n6748);
   U2021 : OAI22_X1 port map( A1 => n1410, A2 => n1423, B1 => n1170, B2 => 
                           n1412, ZN => n6749);
   U2022 : OAI22_X1 port map( A1 => n1410, A2 => n1424, B1 => n1172, B2 => 
                           n1412, ZN => n6750);
   U2023 : OAI22_X1 port map( A1 => n1410, A2 => n1425, B1 => n1496, B2 => 
                           n1412, ZN => n6751);
   U2027 : OAI22_X1 port map( A1 => n1410, A2 => n1429, B1 => n1496, B2 => 
                           n1412, ZN => n6755);
   U2028 : OAI22_X1 port map( A1 => n1410, A2 => n1430, B1 => n1179, B2 => 
                           n1412, ZN => n6756);
   U2029 : OAI22_X1 port map( A1 => n1410, A2 => n1431, B1 => n1181, B2 => 
                           n1412, ZN => n6757);
   U2030 : OAI22_X1 port map( A1 => n1410, A2 => n1432, B1 => n1183, B2 => 
                           n1412, ZN => n6758);
   U2031 : OAI22_X1 port map( A1 => n1410, A2 => n1433, B1 => n1185, B2 => 
                           n1412, ZN => n6759);
   U2032 : OAI22_X1 port map( A1 => n1410, A2 => n1434, B1 => n1187, B2 => 
                           n1412, ZN => n6760);
   U2033 : OAI22_X1 port map( A1 => n1410, A2 => n1435, B1 => n1189, B2 => 
                           n1412, ZN => n6761);
   U2034 : OAI22_X1 port map( A1 => n1410, A2 => n1436, B1 => n1191, B2 => 
                           n1412, ZN => n6762);
   U2035 : OAI22_X1 port map( A1 => n1410, A2 => n1437, B1 => n1193, B2 => 
                           n1412, ZN => n6763);
   U2036 : OAI22_X1 port map( A1 => n1410, A2 => n1438, B1 => n1195, B2 => 
                           n1412, ZN => n6764);
   U2037 : OAI22_X1 port map( A1 => n1410, A2 => n1439, B1 => n1197, B2 => 
                           n1412, ZN => n6765);
   U2038 : OAI22_X1 port map( A1 => n1410, A2 => n1440, B1 => n1199, B2 => 
                           n1412, ZN => n6766);
   U2039 : OAI22_X1 port map( A1 => n1410, A2 => n1441, B1 => n1201, B2 => 
                           n1412, ZN => n6767);
   U2040 : OAI22_X1 port map( A1 => n1410, A2 => n1442, B1 => n1203, B2 => 
                           n1412, ZN => n6768);
   U2041 : OAI22_X1 port map( A1 => n1410, A2 => n1443, B1 => n1205, B2 => 
                           n1412, ZN => n6769);
   U2045 : OAI22_X1 port map( A1 => n1444, A2 => n1445, B1 => n1147, B2 => 
                           n1427, ZN => n6770);
   U2046 : OAI22_X1 port map( A1 => n1444, A2 => n1447, B1 => n1150, B2 => 
                           n1428, ZN => n6771);
   U2047 : OAI22_X1 port map( A1 => n1444, A2 => n1448, B1 => n1152, B2 => 
                           n1428, ZN => n6772);
   U2048 : OAI22_X1 port map( A1 => n1444, A2 => n1449, B1 => n1154, B2 => 
                           n1428, ZN => n6773);
   U2049 : OAI22_X1 port map( A1 => n1444, A2 => n1450, B1 => n1156, B2 => 
                           n1428, ZN => n6774);
   U2050 : OAI22_X1 port map( A1 => n1444, A2 => n1451, B1 => n1158, B2 => 
                           n1427, ZN => n6775);
   U2051 : OAI22_X1 port map( A1 => n1444, A2 => n1452, B1 => n1160, B2 => 
                           n1428, ZN => n6776);
   U2052 : OAI22_X1 port map( A1 => n1444, A2 => n1453, B1 => n1162, B2 => 
                           n1427, ZN => n6777);
   U2053 : OAI22_X1 port map( A1 => n1444, A2 => n1454, B1 => n1164, B2 => 
                           n1428, ZN => n6778);
   U2054 : OAI22_X1 port map( A1 => n1444, A2 => n1455, B1 => n1166, B2 => 
                           n1427, ZN => n6779);
   U2055 : OAI22_X1 port map( A1 => n1444, A2 => n1456, B1 => n1168, B2 => 
                           n1428, ZN => n6780);
   U2056 : OAI22_X1 port map( A1 => n1444, A2 => n1457, B1 => n1170, B2 => 
                           n1428, ZN => n6781);
   U2057 : OAI22_X1 port map( A1 => n1444, A2 => n1458, B1 => n1172, B2 => 
                           n1428, ZN => n6782);
   U2058 : OAI22_X1 port map( A1 => n1444, A2 => n1459, B1 => n3529, B2 => 
                           n1428, ZN => n6783);
   U2059 : OAI22_X1 port map( A1 => n1444, A2 => n1460, B1 => n3529, B2 => 
                           n1428, ZN => n6784);
   U2060 : OAI22_X1 port map( A1 => n1444, A2 => n1461, B1 => n3529, B2 => 
                           n1428, ZN => n6785);
   U2061 : OAI22_X1 port map( A1 => n1444, A2 => n1462, B1 => n3529, B2 => 
                           n1428, ZN => n6786);
   U2063 : OAI22_X1 port map( A1 => n1444, A2 => n1464, B1 => n1179, B2 => 
                           n1428, ZN => n6788);
   U2064 : OAI22_X1 port map( A1 => n1444, A2 => n1465, B1 => n1181, B2 => 
                           n1428, ZN => n6789);
   U2065 : OAI22_X1 port map( A1 => n1444, A2 => n1466, B1 => n1183, B2 => 
                           n1428, ZN => n6790);
   U2066 : OAI22_X1 port map( A1 => n1444, A2 => n1467, B1 => n1185, B2 => 
                           n1428, ZN => n6791);
   U2067 : OAI22_X1 port map( A1 => n1444, A2 => n1468, B1 => n1187, B2 => 
                           n1428, ZN => n6792);
   U2068 : OAI22_X1 port map( A1 => n1444, A2 => n1469, B1 => n1189, B2 => 
                           n1428, ZN => n6793);
   U2069 : OAI22_X1 port map( A1 => n1444, A2 => n1470, B1 => n1191, B2 => 
                           n1428, ZN => n6794);
   U2070 : OAI22_X1 port map( A1 => n1444, A2 => n1471, B1 => n1193, B2 => 
                           n1428, ZN => n6795);
   U2071 : OAI22_X1 port map( A1 => n1444, A2 => n1472, B1 => n1195, B2 => 
                           n1427, ZN => n6796);
   U2072 : OAI22_X1 port map( A1 => n1444, A2 => n1473, B1 => n1197, B2 => 
                           n1428, ZN => n6797);
   U2073 : OAI22_X1 port map( A1 => n1444, A2 => n1474, B1 => n1199, B2 => 
                           n1428, ZN => n6798);
   U2074 : OAI22_X1 port map( A1 => n1444, A2 => n1475, B1 => n1201, B2 => 
                           n1428, ZN => n6799);
   U2075 : OAI22_X1 port map( A1 => n1444, A2 => n1476, B1 => n1203, B2 => 
                           n1428, ZN => n6800);
   U2076 : OAI22_X1 port map( A1 => n1444, A2 => n1477, B1 => n1205, B2 => 
                           n1428, ZN => n6801);
   U2079 : OAI22_X1 port map( A1 => n1479, A2 => n1480, B1 => n1147, B2 => 
                           n1394, ZN => n6802);
   U2080 : OAI22_X1 port map( A1 => n1479, A2 => n1482, B1 => n1150, B2 => 
                           n1394, ZN => n6803);
   U2081 : OAI22_X1 port map( A1 => n1479, A2 => n1483, B1 => n1152, B2 => 
                           n1392, ZN => n6804);
   U2082 : OAI22_X1 port map( A1 => n1479, A2 => n1484, B1 => n1154, B2 => 
                           n1394, ZN => n6805);
   U2083 : OAI22_X1 port map( A1 => n1479, A2 => n1485, B1 => n1156, B2 => 
                           n1394, ZN => n6806);
   U2084 : OAI22_X1 port map( A1 => n1479, A2 => n1486, B1 => n1158, B2 => 
                           n1392, ZN => n6807);
   U2085 : OAI22_X1 port map( A1 => n1479, A2 => n1487, B1 => n1160, B2 => 
                           n1394, ZN => n6808);
   U2086 : OAI22_X1 port map( A1 => n1479, A2 => n1488, B1 => n1162, B2 => 
                           n1392, ZN => n6809);
   U2087 : OAI22_X1 port map( A1 => n1479, A2 => n1489, B1 => n1164, B2 => 
                           n1394, ZN => n6810);
   U2088 : OAI22_X1 port map( A1 => n1479, A2 => n1490, B1 => n1166, B2 => 
                           n1394, ZN => n6811);
   U2089 : OAI22_X1 port map( A1 => n1479, A2 => n1491, B1 => n1168, B2 => 
                           n1394, ZN => n6812);
   U2090 : OAI22_X1 port map( A1 => n1479, A2 => n1492, B1 => n1170, B2 => 
                           n1394, ZN => n6813);
   U2091 : OAI22_X1 port map( A1 => n1479, A2 => n1493, B1 => n1172, B2 => 
                           n1394, ZN => n6814);
   U2092 : OAI22_X1 port map( A1 => n1479, A2 => n1494, B1 => n3529, B2 => 
                           n1394, ZN => n6815);
   U2093 : OAI22_X1 port map( A1 => n1479, A2 => n1495, B1 => n3529, B2 => 
                           n1394, ZN => n6816);
   U2095 : OAI22_X1 port map( A1 => n1479, A2 => n1497, B1 => n3529, B2 => 
                           n1392, ZN => n6818);
   U2097 : OAI22_X1 port map( A1 => n1479, A2 => n1499, B1 => n1179, B2 => 
                           n1394, ZN => n6820);
   U2098 : OAI22_X1 port map( A1 => n1479, A2 => n1500, B1 => n1181, B2 => 
                           n1394, ZN => n6821);
   U2099 : OAI22_X1 port map( A1 => n1479, A2 => n1501, B1 => n1183, B2 => 
                           n1394, ZN => n6822);
   U2100 : OAI22_X1 port map( A1 => n1479, A2 => n1502, B1 => n1185, B2 => 
                           n1394, ZN => n6823);
   U2101 : OAI22_X1 port map( A1 => n1479, A2 => n1503, B1 => n1187, B2 => 
                           n1394, ZN => n6824);
   U2102 : OAI22_X1 port map( A1 => n1479, A2 => n1504, B1 => n1189, B2 => 
                           n1394, ZN => n6825);
   U2103 : OAI22_X1 port map( A1 => n1479, A2 => n1505, B1 => n1191, B2 => 
                           n1394, ZN => n6826);
   U2104 : OAI22_X1 port map( A1 => n1479, A2 => n1506, B1 => n1193, B2 => 
                           n1394, ZN => n6827);
   U2105 : OAI22_X1 port map( A1 => n1479, A2 => n1507, B1 => n1195, B2 => 
                           n1394, ZN => n6828);
   U2106 : OAI22_X1 port map( A1 => n1479, A2 => n1508, B1 => n1197, B2 => 
                           n1394, ZN => n6829);
   U2107 : OAI22_X1 port map( A1 => n1479, A2 => n1509, B1 => n1199, B2 => 
                           n1394, ZN => n6830);
   U2108 : OAI22_X1 port map( A1 => n1479, A2 => n1510, B1 => n1201, B2 => 
                           n1394, ZN => n6831);
   U2109 : OAI22_X1 port map( A1 => n1479, A2 => n1511, B1 => n1203, B2 => 
                           n1394, ZN => n6832);
   U2110 : OAI22_X1 port map( A1 => n1479, A2 => n1512, B1 => n1205, B2 => 
                           n1394, ZN => n6833);
   U2113 : OAI22_X1 port map( A1 => n3810, A2 => n1514, B1 => n1147, B2 => 
                           n1515, ZN => n6834);
   U2115 : OAI22_X1 port map( A1 => n3810, A2 => n1516, B1 => n1150, B2 => 
                           n1515, ZN => n6835);
   U2117 : OAI22_X1 port map( A1 => n3810, A2 => n1517, B1 => n1152, B2 => 
                           n1515, ZN => n6836);
   U2119 : OAI22_X1 port map( A1 => n3810, A2 => n1518, B1 => n1154, B2 => 
                           n1515, ZN => n6837);
   U2121 : OAI22_X1 port map( A1 => n3810, A2 => n1519, B1 => n1156, B2 => 
                           n1515, ZN => n6838);
   U2123 : OAI22_X1 port map( A1 => n3810, A2 => n1520, B1 => n1158, B2 => 
                           n1515, ZN => n6839);
   U2125 : OAI22_X1 port map( A1 => n3810, A2 => n1521, B1 => n1160, B2 => 
                           n1515, ZN => n6840);
   U2127 : OAI22_X1 port map( A1 => n3810, A2 => n1522, B1 => n1162, B2 => 
                           n1515, ZN => n6841);
   U2129 : OAI22_X1 port map( A1 => n3810, A2 => n1523, B1 => n1164, B2 => 
                           n1515, ZN => n6842);
   U2131 : OAI22_X1 port map( A1 => n3810, A2 => n1524, B1 => n1166, B2 => 
                           n1515, ZN => n6843);
   U2133 : OAI22_X1 port map( A1 => n3810, A2 => n1525, B1 => n1168, B2 => 
                           n1515, ZN => n6844);
   U2135 : OAI22_X1 port map( A1 => n3810, A2 => n1526, B1 => n1170, B2 => 
                           n1515, ZN => n6845);
   U2137 : OAI22_X1 port map( A1 => n3810, A2 => n1527, B1 => n1172, B2 => 
                           n1515, ZN => n6846);
   U2139 : INV_X1 port map( A => n1528, ZN => n6847);
   U2140 : AOI22_X1 port map( A1 => n1515, A2 => pc_lut_21_4_port, B1 => n3521,
                           B2 => n3810, ZN => n1528);
   U2141 : INV_X1 port map( A => n1529, ZN => n6848);
   U2142 : AOI22_X1 port map( A1 => n1515, A2 => pc_lut_21_2_port, B1 => n3521,
                           B2 => n3810, ZN => n1529);
   U2143 : INV_X1 port map( A => n1530, ZN => n6849);
   U2144 : AOI22_X1 port map( A1 => n1515, A2 => pc_lut_21_0_port, B1 => n3521,
                           B2 => n3810, ZN => n1530);
   U2147 : OAI22_X1 port map( A1 => n3810, A2 => n1531, B1 => n1179, B2 => 
                           n1515, ZN => n6852);
   U2149 : OAI22_X1 port map( A1 => n3810, A2 => n1532, B1 => n1181, B2 => 
                           n1515, ZN => n6853);
   U2151 : OAI22_X1 port map( A1 => n3810, A2 => n1533, B1 => n1183, B2 => 
                           n1515, ZN => n6854);
   U2153 : OAI22_X1 port map( A1 => n3810, A2 => n1534, B1 => n1185, B2 => 
                           n1515, ZN => n6855);
   U2155 : OAI22_X1 port map( A1 => n3810, A2 => n1535, B1 => n1187, B2 => 
                           n1515, ZN => n6856);
   U2157 : OAI22_X1 port map( A1 => n3810, A2 => n1536, B1 => n1189, B2 => 
                           n1515, ZN => n6857);
   U2159 : OAI22_X1 port map( A1 => n3810, A2 => n1537, B1 => n1191, B2 => 
                           n1515, ZN => n6858);
   U2161 : OAI22_X1 port map( A1 => n3810, A2 => n1538, B1 => n1193, B2 => 
                           n1515, ZN => n6859);
   U2163 : OAI22_X1 port map( A1 => n3810, A2 => n1539, B1 => n1195, B2 => 
                           n1515, ZN => n6860);
   U2165 : OAI22_X1 port map( A1 => n3810, A2 => n1540, B1 => n1197, B2 => 
                           n1515, ZN => n6861);
   U2167 : OAI22_X1 port map( A1 => n3810, A2 => n1541, B1 => n1199, B2 => 
                           n1515, ZN => n6862);
   U2169 : OAI22_X1 port map( A1 => n3810, A2 => n1542, B1 => n1201, B2 => 
                           n1515, ZN => n6863);
   U2171 : OAI22_X1 port map( A1 => n3810, A2 => n1543, B1 => n1203, B2 => 
                           n1515, ZN => n6864);
   U2173 : OAI22_X1 port map( A1 => n3810, A2 => n1544, B1 => n1205, B2 => 
                           n1515, ZN => n6865);
   U2177 : OAI22_X1 port map( A1 => n3800, A2 => n1546, B1 => n1147, B2 => 
                           n1547, ZN => n6866);
   U2179 : OAI22_X1 port map( A1 => n3800, A2 => n1548, B1 => n1150, B2 => 
                           n1547, ZN => n6867);
   U2181 : OAI22_X1 port map( A1 => n3800, A2 => n1549, B1 => n1152, B2 => 
                           n1547, ZN => n6868);
   U2183 : OAI22_X1 port map( A1 => n3800, A2 => n1550, B1 => n1154, B2 => 
                           n1547, ZN => n6869);
   U2185 : OAI22_X1 port map( A1 => n3800, A2 => n1551, B1 => n1156, B2 => 
                           n1547, ZN => n6870);
   U2187 : OAI22_X1 port map( A1 => n3800, A2 => n1552, B1 => n1158, B2 => 
                           n1547, ZN => n6871);
   U2189 : OAI22_X1 port map( A1 => n3800, A2 => n1553, B1 => n1160, B2 => 
                           n1547, ZN => n6872);
   U2191 : OAI22_X1 port map( A1 => n3800, A2 => n1554, B1 => n1162, B2 => 
                           n1547, ZN => n6873);
   U2193 : OAI22_X1 port map( A1 => n3800, A2 => n1555, B1 => n1164, B2 => 
                           n1547, ZN => n6874);
   U2195 : OAI22_X1 port map( A1 => n3800, A2 => n1556, B1 => n1166, B2 => 
                           n1547, ZN => n6875);
   U2197 : OAI22_X1 port map( A1 => n3800, A2 => n1557, B1 => n1168, B2 => 
                           n1547, ZN => n6876);
   U2199 : OAI22_X1 port map( A1 => n3800, A2 => n1558, B1 => n1170, B2 => 
                           n1547, ZN => n6877);
   U2201 : OAI22_X1 port map( A1 => n3800, A2 => n1559, B1 => n1172, B2 => 
                           n1547, ZN => n6878);
   U2203 : INV_X1 port map( A => n1560, ZN => n6879);
   U2204 : AOI22_X1 port map( A1 => n1547, A2 => pc_lut_20_4_port, B1 => n3521,
                           B2 => n3800, ZN => n1560);
   U2205 : INV_X1 port map( A => n1561, ZN => n6880);
   U2206 : AOI22_X1 port map( A1 => n1547, A2 => pc_lut_20_2_port, B1 => n3521,
                           B2 => n3800, ZN => n1561);
   U2210 : OAI22_X1 port map( A1 => n3800, A2 => n1562, B1 => n1179, B2 => 
                           n1547, ZN => n6884);
   U2212 : OAI22_X1 port map( A1 => n3800, A2 => n1563, B1 => n1181, B2 => 
                           n1547, ZN => n6885);
   U2214 : OAI22_X1 port map( A1 => n3800, A2 => n1564, B1 => n1183, B2 => 
                           n1547, ZN => n6886);
   U2216 : OAI22_X1 port map( A1 => n3800, A2 => n1565, B1 => n1185, B2 => 
                           n1547, ZN => n6887);
   U2218 : OAI22_X1 port map( A1 => n3800, A2 => n1566, B1 => n1187, B2 => 
                           n1547, ZN => n6888);
   U2220 : OAI22_X1 port map( A1 => n3800, A2 => n1567, B1 => n1189, B2 => 
                           n1547, ZN => n6889);
   U2222 : OAI22_X1 port map( A1 => n3800, A2 => n1568, B1 => n1191, B2 => 
                           n1547, ZN => n6890);
   U2224 : OAI22_X1 port map( A1 => n3800, A2 => n1569, B1 => n1193, B2 => 
                           n1547, ZN => n6891);
   U2226 : OAI22_X1 port map( A1 => n3800, A2 => n1570, B1 => n1195, B2 => 
                           n1547, ZN => n6892);
   U2228 : OAI22_X1 port map( A1 => n3800, A2 => n1571, B1 => n1197, B2 => 
                           n1547, ZN => n6893);
   U2230 : OAI22_X1 port map( A1 => n3800, A2 => n1572, B1 => n1199, B2 => 
                           n1547, ZN => n6894);
   U2232 : OAI22_X1 port map( A1 => n3800, A2 => n1573, B1 => n1201, B2 => 
                           n1547, ZN => n6895);
   U2234 : OAI22_X1 port map( A1 => n3800, A2 => n1574, B1 => n1203, B2 => 
                           n1547, ZN => n6896);
   U2236 : OAI22_X1 port map( A1 => n3800, A2 => n1575, B1 => n1205, B2 => 
                           n1547, ZN => n6897);
   U2240 : AND2_X1 port map( A1 => n1309, A2 => n454, ZN => n1478);
   U2241 : OAI22_X1 port map( A1 => n1576, A2 => n1577, B1 => n1147, B2 => 
                           n3532, ZN => n6898);
   U2243 : OAI22_X1 port map( A1 => n1576, A2 => n1579, B1 => n1150, B2 => 
                           n3532, ZN => n6899);
   U2245 : OAI22_X1 port map( A1 => n1576, A2 => n1580, B1 => n1152, B2 => 
                           n3532, ZN => n6900);
   U2247 : OAI22_X1 port map( A1 => n1576, A2 => n1581, B1 => n1154, B2 => 
                           n3532, ZN => n6901);
   U2249 : OAI22_X1 port map( A1 => n1576, A2 => n1582, B1 => n1156, B2 => 
                           n3533, ZN => n6902);
   U2251 : OAI22_X1 port map( A1 => n1576, A2 => n1583, B1 => n1158, B2 => 
                           n3533, ZN => n6903);
   U2253 : OAI22_X1 port map( A1 => n1576, A2 => n1584, B1 => n1160, B2 => 
                           n3532, ZN => n6904);
   U2255 : OAI22_X1 port map( A1 => n1576, A2 => n1585, B1 => n1162, B2 => 
                           n3533, ZN => n6905);
   U2257 : OAI22_X1 port map( A1 => n1576, A2 => n1586, B1 => n1164, B2 => 
                           n3533, ZN => n6906);
   U2259 : OAI22_X1 port map( A1 => n1576, A2 => n1587, B1 => n1166, B2 => 
                           n3533, ZN => n6907);
   U2261 : OAI22_X1 port map( A1 => n1576, A2 => n1588, B1 => n1168, B2 => 
                           n3532, ZN => n6908);
   U2263 : OAI22_X1 port map( A1 => n1576, A2 => n1589, B1 => n1170, B2 => 
                           n3532, ZN => n6909);
   U2265 : OAI22_X1 port map( A1 => n1576, A2 => n1590, B1 => n1172, B2 => 
                           n3532, ZN => n6910);
   U2267 : INV_X1 port map( A => n1591, ZN => n6911);
   U2268 : AOI22_X1 port map( A1 => n3533, A2 => pc_lut_19_4_port, B1 => n3521,
                           B2 => n1576, ZN => n1591);
   U2270 : INV_X1 port map( A => n1592, ZN => n6913);
   U2271 : AOI22_X1 port map( A1 => n3532, A2 => pc_lut_19_0_port, B1 => n3521,
                           B2 => n1576, ZN => n1592);
   U2272 : INV_X1 port map( A => n1593, ZN => n6914);
   U2273 : AOI22_X1 port map( A1 => n3533, A2 => pc_lut_19_1_port, B1 => n3521,
                           B2 => n1576, ZN => n1593);
   U2275 : OAI22_X1 port map( A1 => n1576, A2 => n1594, B1 => n1179, B2 => 
                           n3532, ZN => n6916);
   U2277 : OAI22_X1 port map( A1 => n1576, A2 => n1595, B1 => n1181, B2 => 
                           n3533, ZN => n6917);
   U2279 : OAI22_X1 port map( A1 => n1576, A2 => n1596, B1 => n1183, B2 => 
                           n3532, ZN => n6918);
   U2281 : OAI22_X1 port map( A1 => n1576, A2 => n1597, B1 => n1185, B2 => 
                           n3533, ZN => n6919);
   U2283 : OAI22_X1 port map( A1 => n1576, A2 => n1598, B1 => n1187, B2 => 
                           n3532, ZN => n6920);
   U2285 : OAI22_X1 port map( A1 => n1576, A2 => n1599, B1 => n1189, B2 => 
                           n3533, ZN => n6921);
   U2287 : OAI22_X1 port map( A1 => n1576, A2 => n1600, B1 => n1191, B2 => 
                           n3533, ZN => n6922);
   U2289 : OAI22_X1 port map( A1 => n1576, A2 => n1601, B1 => n1193, B2 => 
                           n3533, ZN => n6923);
   U2291 : OAI22_X1 port map( A1 => n1576, A2 => n1602, B1 => n1195, B2 => 
                           n3532, ZN => n6924);
   U2293 : OAI22_X1 port map( A1 => n1576, A2 => n1603, B1 => n1197, B2 => 
                           n3533, ZN => n6925);
   U2295 : OAI22_X1 port map( A1 => n1576, A2 => n1604, B1 => n1199, B2 => 
                           n3532, ZN => n6926);
   U2297 : OAI22_X1 port map( A1 => n1576, A2 => n1605, B1 => n1201, B2 => 
                           n3533, ZN => n6927);
   U2299 : OAI22_X1 port map( A1 => n1576, A2 => n1606, B1 => n1203, B2 => 
                           n3532, ZN => n6928);
   U2301 : OAI22_X1 port map( A1 => n1576, A2 => n1607, B1 => n1205, B2 => 
                           n3533, ZN => n6929);
   U2304 : NAND2_X1 port map( A1 => n1608, A2 => n38, ZN => n1578);
   U2305 : OAI22_X1 port map( A1 => n1609, A2 => n1610, B1 => n1147, B2 => n558
                           , ZN => n6930);
   U2307 : OAI22_X1 port map( A1 => n1609, A2 => n1612, B1 => n1150, B2 => n768
                           , ZN => n6931);
   U2309 : OAI22_X1 port map( A1 => n1609, A2 => n1613, B1 => n1152, B2 => n768
                           , ZN => n6932);
   U2311 : OAI22_X1 port map( A1 => n1609, A2 => n1614, B1 => n1154, B2 => n768
                           , ZN => n6933);
   U2313 : OAI22_X1 port map( A1 => n1609, A2 => n1615, B1 => n1156, B2 => n768
                           , ZN => n6934);
   U2315 : OAI22_X1 port map( A1 => n1609, A2 => n1616, B1 => n1158, B2 => n768
                           , ZN => n6935);
   U2317 : OAI22_X1 port map( A1 => n1609, A2 => n1617, B1 => n1160, B2 => n768
                           , ZN => n6936);
   U2319 : OAI22_X1 port map( A1 => n1609, A2 => n1618, B1 => n1162, B2 => n768
                           , ZN => n6937);
   U2321 : OAI22_X1 port map( A1 => n1609, A2 => n1619, B1 => n1164, B2 => n768
                           , ZN => n6938);
   U2323 : OAI22_X1 port map( A1 => n1609, A2 => n1620, B1 => n1166, B2 => n768
                           , ZN => n6939);
   U2325 : OAI22_X1 port map( A1 => n1609, A2 => n1621, B1 => n1168, B2 => n768
                           , ZN => n6940);
   U2327 : OAI22_X1 port map( A1 => n1609, A2 => n1622, B1 => n1170, B2 => n768
                           , ZN => n6941);
   U2329 : OAI22_X1 port map( A1 => n1609, A2 => n1623, B1 => n1172, B2 => n768
                           , ZN => n6942);
   U2331 : INV_X1 port map( A => n1624, ZN => n6943);
   U2332 : AOI22_X1 port map( A1 => n558, A2 => pc_lut_18_4_port, B1 => n3521, 
                           B2 => n1609, ZN => n1624);
   U2335 : INV_X1 port map( A => n1625, ZN => n6946);
   U2336 : AOI22_X1 port map( A1 => n558, A2 => pc_lut_18_1_port, B1 => n3521, 
                           B2 => n1609, ZN => n1625);
   U2338 : OAI22_X1 port map( A1 => n1609, A2 => n1626, B1 => n1179, B2 => n768
                           , ZN => n6948);
   U2340 : OAI22_X1 port map( A1 => n1609, A2 => n1627, B1 => n1181, B2 => n768
                           , ZN => n6949);
   U2342 : OAI22_X1 port map( A1 => n1609, A2 => n1628, B1 => n1183, B2 => n768
                           , ZN => n6950);
   U2344 : OAI22_X1 port map( A1 => n1609, A2 => n1629, B1 => n1185, B2 => n768
                           , ZN => n6951);
   U2346 : OAI22_X1 port map( A1 => n1609, A2 => n1630, B1 => n1187, B2 => n768
                           , ZN => n6952);
   U2348 : OAI22_X1 port map( A1 => n1609, A2 => n1631, B1 => n1189, B2 => n768
                           , ZN => n6953);
   U2350 : OAI22_X1 port map( A1 => n1609, A2 => n1632, B1 => n1191, B2 => n768
                           , ZN => n6954);
   U2352 : OAI22_X1 port map( A1 => n1609, A2 => n1633, B1 => n1193, B2 => n768
                           , ZN => n6955);
   U2354 : OAI22_X1 port map( A1 => n1609, A2 => n1634, B1 => n1195, B2 => n768
                           , ZN => n6956);
   U2356 : OAI22_X1 port map( A1 => n1609, A2 => n1635, B1 => n1197, B2 => n768
                           , ZN => n6957);
   U2358 : OAI22_X1 port map( A1 => n1609, A2 => n1636, B1 => n1199, B2 => n768
                           , ZN => n6958);
   U2360 : OAI22_X1 port map( A1 => n1609, A2 => n1637, B1 => n1201, B2 => n768
                           , ZN => n6959);
   U2362 : OAI22_X1 port map( A1 => n1609, A2 => n1638, B1 => n1203, B2 => n768
                           , ZN => n6960);
   U2364 : OAI22_X1 port map( A1 => n1609, A2 => n1639, B1 => n1205, B2 => n768
                           , ZN => n6961);
   U2368 : OAI22_X1 port map( A1 => n1640, A2 => n1641, B1 => n1147, B2 => 
                           n1642, ZN => n6962);
   U2369 : OAI22_X1 port map( A1 => n1640, A2 => n1643, B1 => n1150, B2 => 
                           n1642, ZN => n6963);
   U2370 : OAI22_X1 port map( A1 => n1640, A2 => n1644, B1 => n1152, B2 => 
                           n1642, ZN => n6964);
   U2371 : OAI22_X1 port map( A1 => n1640, A2 => n1645, B1 => n1154, B2 => 
                           n1642, ZN => n6965);
   U2372 : OAI22_X1 port map( A1 => n1640, A2 => n1646, B1 => n1156, B2 => 
                           n1642, ZN => n6966);
   U2373 : OAI22_X1 port map( A1 => n1640, A2 => n1647, B1 => n1158, B2 => 
                           n1642, ZN => n6967);
   U2374 : OAI22_X1 port map( A1 => n1640, A2 => n1648, B1 => n1160, B2 => 
                           n1642, ZN => n6968);
   U2375 : OAI22_X1 port map( A1 => n1640, A2 => n1649, B1 => n1162, B2 => 
                           n1642, ZN => n6969);
   U2376 : OAI22_X1 port map( A1 => n1640, A2 => n1650, B1 => n1164, B2 => 
                           n1642, ZN => n6970);
   U2377 : OAI22_X1 port map( A1 => n1640, A2 => n1651, B1 => n1166, B2 => 
                           n1642, ZN => n6971);
   U2378 : OAI22_X1 port map( A1 => n1640, A2 => n1652, B1 => n1168, B2 => 
                           n1642, ZN => n6972);
   U2379 : OAI22_X1 port map( A1 => n1640, A2 => n1653, B1 => n1170, B2 => 
                           n1642, ZN => n6973);
   U2380 : OAI22_X1 port map( A1 => n1640, A2 => n1654, B1 => n1172, B2 => 
                           n1642, ZN => n6974);
   U2381 : OAI22_X1 port map( A1 => n1640, A2 => n1655, B1 => n1496, B2 => 
                           n1642, ZN => n6975);
   U2383 : OAI22_X1 port map( A1 => n1640, A2 => n1657, B1 => n1496, B2 => 
                           n1642, ZN => n6977);
   U2386 : OAI22_X1 port map( A1 => n1640, A2 => n1660, B1 => n1179, B2 => 
                           n1642, ZN => n6980);
   U2387 : OAI22_X1 port map( A1 => n1640, A2 => n1661, B1 => n1181, B2 => 
                           n1642, ZN => n6981);
   U2388 : OAI22_X1 port map( A1 => n1640, A2 => n1662, B1 => n1183, B2 => 
                           n1642, ZN => n6982);
   U2389 : OAI22_X1 port map( A1 => n1640, A2 => n1663, B1 => n1185, B2 => 
                           n1642, ZN => n6983);
   U2390 : OAI22_X1 port map( A1 => n1640, A2 => n1664, B1 => n1187, B2 => 
                           n1642, ZN => n6984);
   U2391 : OAI22_X1 port map( A1 => n1640, A2 => n1665, B1 => n1189, B2 => 
                           n1642, ZN => n6985);
   U2392 : OAI22_X1 port map( A1 => n1640, A2 => n1666, B1 => n1191, B2 => 
                           n1642, ZN => n6986);
   U2393 : OAI22_X1 port map( A1 => n1640, A2 => n1667, B1 => n1193, B2 => 
                           n1642, ZN => n6987);
   U2394 : OAI22_X1 port map( A1 => n1640, A2 => n1668, B1 => n1195, B2 => 
                           n1642, ZN => n6988);
   U2395 : OAI22_X1 port map( A1 => n1640, A2 => n1669, B1 => n1197, B2 => 
                           n1642, ZN => n6989);
   U2396 : OAI22_X1 port map( A1 => n1640, A2 => n1670, B1 => n1199, B2 => 
                           n1642, ZN => n6990);
   U2397 : OAI22_X1 port map( A1 => n1640, A2 => n1671, B1 => n1201, B2 => 
                           n1642, ZN => n6991);
   U2398 : OAI22_X1 port map( A1 => n1640, A2 => n1672, B1 => n1203, B2 => 
                           n1642, ZN => n6992);
   U2399 : OAI22_X1 port map( A1 => n1640, A2 => n1673, B1 => n1205, B2 => 
                           n1642, ZN => n6993);
   U2402 : OAI22_X1 port map( A1 => n1674, A2 => n1675, B1 => n1147, B2 => 
                           n1676, ZN => n6994);
   U2403 : OAI22_X1 port map( A1 => n1674, A2 => n1677, B1 => n1150, B2 => 
                           n1676, ZN => n6995);
   U2404 : OAI22_X1 port map( A1 => n1674, A2 => n1678, B1 => n1152, B2 => 
                           n1676, ZN => n6996);
   U2405 : OAI22_X1 port map( A1 => n1674, A2 => n1679, B1 => n1154, B2 => 
                           n1676, ZN => n6997);
   U2406 : OAI22_X1 port map( A1 => n1674, A2 => n1680, B1 => n1156, B2 => 
                           n1676, ZN => n6998);
   U2407 : OAI22_X1 port map( A1 => n1674, A2 => n1681, B1 => n1158, B2 => 
                           n1676, ZN => n6999);
   U2408 : OAI22_X1 port map( A1 => n1674, A2 => n1682, B1 => n1160, B2 => 
                           n1676, ZN => n7000);
   U2409 : OAI22_X1 port map( A1 => n1674, A2 => n1683, B1 => n1162, B2 => 
                           n1676, ZN => n7001);
   U2410 : OAI22_X1 port map( A1 => n1674, A2 => n1684, B1 => n1164, B2 => 
                           n1676, ZN => n7002);
   U2411 : OAI22_X1 port map( A1 => n1674, A2 => n1685, B1 => n1166, B2 => 
                           n1676, ZN => n7003);
   U2412 : OAI22_X1 port map( A1 => n1674, A2 => n1686, B1 => n1168, B2 => 
                           n1676, ZN => n7004);
   U2413 : OAI22_X1 port map( A1 => n1674, A2 => n1687, B1 => n1170, B2 => 
                           n1676, ZN => n7005);
   U2414 : OAI22_X1 port map( A1 => n1674, A2 => n1688, B1 => n1172, B2 => 
                           n1676, ZN => n7006);
   U2415 : OAI22_X1 port map( A1 => n1674, A2 => n1689, B1 => n1496, B2 => 
                           n1676, ZN => n7007);
   U2420 : OAI22_X1 port map( A1 => n1674, A2 => n1694, B1 => n1179, B2 => 
                           n1676, ZN => n7012);
   U2421 : OAI22_X1 port map( A1 => n1674, A2 => n1695, B1 => n1181, B2 => 
                           n1676, ZN => n7013);
   U2422 : OAI22_X1 port map( A1 => n1674, A2 => n1696, B1 => n1183, B2 => 
                           n1676, ZN => n7014);
   U2423 : OAI22_X1 port map( A1 => n1674, A2 => n1697, B1 => n1185, B2 => 
                           n1676, ZN => n7015);
   U2424 : OAI22_X1 port map( A1 => n1674, A2 => n1698, B1 => n1187, B2 => 
                           n1676, ZN => n7016);
   U2425 : OAI22_X1 port map( A1 => n1674, A2 => n1699, B1 => n1189, B2 => 
                           n1676, ZN => n7017);
   U2426 : OAI22_X1 port map( A1 => n1674, A2 => n1700, B1 => n1191, B2 => 
                           n1676, ZN => n7018);
   U2427 : OAI22_X1 port map( A1 => n1674, A2 => n1701, B1 => n1193, B2 => 
                           n1676, ZN => n7019);
   U2428 : OAI22_X1 port map( A1 => n1674, A2 => n1702, B1 => n1195, B2 => 
                           n1676, ZN => n7020);
   U2429 : OAI22_X1 port map( A1 => n1674, A2 => n1703, B1 => n1197, B2 => 
                           n1676, ZN => n7021);
   U2430 : OAI22_X1 port map( A1 => n1674, A2 => n1704, B1 => n1199, B2 => 
                           n1676, ZN => n7022);
   U2431 : OAI22_X1 port map( A1 => n1674, A2 => n1705, B1 => n1201, B2 => 
                           n1676, ZN => n7023);
   U2432 : OAI22_X1 port map( A1 => n1674, A2 => n1706, B1 => n1203, B2 => 
                           n1676, ZN => n7024);
   U2433 : OAI22_X1 port map( A1 => n1674, A2 => n1707, B1 => n1205, B2 => 
                           n1676, ZN => n7025);
   U2437 : NOR2_X1 port map( A1 => n3793, A2 => n1143, ZN => n1309);
   U2438 : INV_X1 port map( A => PC_write(4), ZN => n1143);
   U2439 : OAI22_X1 port map( A1 => n3537, A2 => n1710, B1 => n1147, B2 => 
                           n1711, ZN => n7026);
   U2441 : OAI22_X1 port map( A1 => n3537, A2 => n1712, B1 => n1150, B2 => 
                           n1711, ZN => n7027);
   U2443 : OAI22_X1 port map( A1 => n3537, A2 => n1713, B1 => n1152, B2 => 
                           n1711, ZN => n7028);
   U2445 : OAI22_X1 port map( A1 => n3537, A2 => n1714, B1 => n1154, B2 => 
                           n1711, ZN => n7029);
   U2447 : OAI22_X1 port map( A1 => n3537, A2 => n1715, B1 => n1156, B2 => 
                           n1711, ZN => n7030);
   U2449 : OAI22_X1 port map( A1 => n3537, A2 => n1716, B1 => n1158, B2 => 
                           n1711, ZN => n7031);
   U2451 : OAI22_X1 port map( A1 => n3537, A2 => n1717, B1 => n1160, B2 => 
                           n1711, ZN => n7032);
   U2453 : OAI22_X1 port map( A1 => n3537, A2 => n1718, B1 => n1162, B2 => 
                           n1711, ZN => n7033);
   U2455 : OAI22_X1 port map( A1 => n3537, A2 => n1719, B1 => n1164, B2 => 
                           n1711, ZN => n7034);
   U2457 : OAI22_X1 port map( A1 => n3537, A2 => n1720, B1 => n1166, B2 => 
                           n1711, ZN => n7035);
   U2459 : OAI22_X1 port map( A1 => n3537, A2 => n1721, B1 => n1168, B2 => 
                           n1711, ZN => n7036);
   U2461 : OAI22_X1 port map( A1 => n3537, A2 => n1722, B1 => n1170, B2 => 
                           n1711, ZN => n7037);
   U2463 : OAI22_X1 port map( A1 => n3537, A2 => n1723, B1 => n1172, B2 => 
                           n1711, ZN => n7038);
   U2466 : INV_X1 port map( A => n1724, ZN => n7040);
   U2467 : AOI22_X1 port map( A1 => n1711, A2 => pc_lut_15_2_port, B1 => n3521,
                           B2 => n3537, ZN => n1724);
   U2468 : INV_X1 port map( A => n1725, ZN => n7041);
   U2469 : AOI22_X1 port map( A1 => n1711, A2 => pc_lut_15_0_port, B1 => n3521,
                           B2 => n3537, ZN => n1725);
   U2470 : INV_X1 port map( A => n1726, ZN => n7042);
   U2471 : AOI22_X1 port map( A1 => n1711, A2 => pc_lut_15_1_port, B1 => n3521,
                           B2 => n3537, ZN => n1726);
   U2472 : INV_X1 port map( A => n1727, ZN => n7043);
   U2473 : AOI22_X1 port map( A1 => n1711, A2 => pc_lut_15_3_port, B1 => n3521,
                           B2 => n3537, ZN => n1727);
   U2474 : OAI22_X1 port map( A1 => n3537, A2 => n1728, B1 => n1179, B2 => 
                           n1711, ZN => n7044);
   U2476 : OAI22_X1 port map( A1 => n3537, A2 => n1729, B1 => n1181, B2 => 
                           n1711, ZN => n7045);
   U2478 : OAI22_X1 port map( A1 => n3537, A2 => n1730, B1 => n1183, B2 => 
                           n1711, ZN => n7046);
   U2480 : OAI22_X1 port map( A1 => n3537, A2 => n1731, B1 => n1185, B2 => 
                           n1711, ZN => n7047);
   U2482 : OAI22_X1 port map( A1 => n3537, A2 => n1732, B1 => n1187, B2 => 
                           n1711, ZN => n7048);
   U2484 : OAI22_X1 port map( A1 => n3537, A2 => n1733, B1 => n1189, B2 => 
                           n1711, ZN => n7049);
   U2486 : OAI22_X1 port map( A1 => n3537, A2 => n1734, B1 => n1191, B2 => 
                           n1711, ZN => n7050);
   U2488 : OAI22_X1 port map( A1 => n3537, A2 => n1735, B1 => n1193, B2 => 
                           n1711, ZN => n7051);
   U2490 : OAI22_X1 port map( A1 => n3537, A2 => n1736, B1 => n1195, B2 => 
                           n1711, ZN => n7052);
   U2492 : OAI22_X1 port map( A1 => n3537, A2 => n1737, B1 => n1197, B2 => 
                           n1711, ZN => n7053);
   U2494 : OAI22_X1 port map( A1 => n3537, A2 => n1738, B1 => n1199, B2 => 
                           n1711, ZN => n7054);
   U2496 : OAI22_X1 port map( A1 => n3537, A2 => n1739, B1 => n1201, B2 => 
                           n1711, ZN => n7055);
   U2498 : OAI22_X1 port map( A1 => n3537, A2 => n1740, B1 => n1203, B2 => 
                           n1711, ZN => n7056);
   U2500 : OAI22_X1 port map( A1 => n3537, A2 => n1741, B1 => n1205, B2 => 
                           n1711, ZN => n7057);
   U2504 : OAI22_X1 port map( A1 => n3535, A2 => n1744, B1 => n1147, B2 => 
                           n1745, ZN => n7058);
   U2506 : OAI22_X1 port map( A1 => n3535, A2 => n1746, B1 => n1150, B2 => 
                           n1745, ZN => n7059);
   U2508 : OAI22_X1 port map( A1 => n3535, A2 => n1747, B1 => n1152, B2 => 
                           n1745, ZN => n7060);
   U2510 : OAI22_X1 port map( A1 => n3535, A2 => n1748, B1 => n1154, B2 => 
                           n1745, ZN => n7061);
   U2512 : OAI22_X1 port map( A1 => n3535, A2 => n1749, B1 => n1156, B2 => 
                           n1745, ZN => n7062);
   U2514 : OAI22_X1 port map( A1 => n3535, A2 => n1750, B1 => n1158, B2 => 
                           n1745, ZN => n7063);
   U2516 : OAI22_X1 port map( A1 => n3535, A2 => n1751, B1 => n1160, B2 => 
                           n1745, ZN => n7064);
   U2518 : OAI22_X1 port map( A1 => n3535, A2 => n1752, B1 => n1162, B2 => 
                           n1745, ZN => n7065);
   U2520 : OAI22_X1 port map( A1 => n3535, A2 => n1753, B1 => n1164, B2 => 
                           n1745, ZN => n7066);
   U2522 : OAI22_X1 port map( A1 => n3535, A2 => n1754, B1 => n1166, B2 => 
                           n1745, ZN => n7067);
   U2524 : OAI22_X1 port map( A1 => n3535, A2 => n1755, B1 => n1168, B2 => 
                           n1745, ZN => n7068);
   U2526 : OAI22_X1 port map( A1 => n3535, A2 => n1756, B1 => n1170, B2 => 
                           n1745, ZN => n7069);
   U2528 : OAI22_X1 port map( A1 => n3535, A2 => n1757, B1 => n1172, B2 => 
                           n1745, ZN => n7070);
   U2531 : INV_X1 port map( A => n1758, ZN => n7072);
   U2532 : AOI22_X1 port map( A1 => n1745, A2 => pc_lut_14_2_port, B1 => n3521,
                           B2 => n3535, ZN => n1758);
   U2534 : INV_X1 port map( A => n1759, ZN => n7074);
   U2535 : AOI22_X1 port map( A1 => n1745, A2 => pc_lut_14_1_port, B1 => n3521,
                           B2 => n3535, ZN => n1759);
   U2536 : INV_X1 port map( A => n1760, ZN => n7075);
   U2537 : AOI22_X1 port map( A1 => n1745, A2 => pc_lut_14_3_port, B1 => n3521,
                           B2 => n3535, ZN => n1760);
   U2538 : OAI22_X1 port map( A1 => n3535, A2 => n1761, B1 => n1179, B2 => 
                           n1745, ZN => n7076);
   U2540 : OAI22_X1 port map( A1 => n3535, A2 => n1762, B1 => n1181, B2 => 
                           n1745, ZN => n7077);
   U2542 : OAI22_X1 port map( A1 => n3535, A2 => n1763, B1 => n1183, B2 => 
                           n1745, ZN => n7078);
   U2544 : OAI22_X1 port map( A1 => n3535, A2 => n1764, B1 => n1185, B2 => 
                           n1745, ZN => n7079);
   U2546 : OAI22_X1 port map( A1 => n3535, A2 => n1765, B1 => n1187, B2 => 
                           n1745, ZN => n7080);
   U2548 : OAI22_X1 port map( A1 => n3535, A2 => n1766, B1 => n1189, B2 => 
                           n1745, ZN => n7081);
   U2550 : OAI22_X1 port map( A1 => n3535, A2 => n1767, B1 => n1191, B2 => 
                           n1745, ZN => n7082);
   U2552 : OAI22_X1 port map( A1 => n3535, A2 => n1768, B1 => n1193, B2 => 
                           n1745, ZN => n7083);
   U2554 : OAI22_X1 port map( A1 => n3535, A2 => n1769, B1 => n1195, B2 => 
                           n1745, ZN => n7084);
   U2556 : OAI22_X1 port map( A1 => n3535, A2 => n1770, B1 => n1197, B2 => 
                           n1745, ZN => n7085);
   U2558 : OAI22_X1 port map( A1 => n3535, A2 => n1771, B1 => n1199, B2 => 
                           n1745, ZN => n7086);
   U2560 : OAI22_X1 port map( A1 => n3535, A2 => n1772, B1 => n1201, B2 => 
                           n1745, ZN => n7087);
   U2562 : OAI22_X1 port map( A1 => n3535, A2 => n1773, B1 => n1203, B2 => 
                           n1745, ZN => n7088);
   U2564 : OAI22_X1 port map( A1 => n3535, A2 => n1774, B1 => n1205, B2 => 
                           n1745, ZN => n7089);
   U2568 : OAI22_X1 port map( A1 => n1775, A2 => n1776, B1 => n1147, B2 => 
                           n1777, ZN => n7090);
   U2569 : OAI22_X1 port map( A1 => n1775, A2 => n1778, B1 => n1150, B2 => 
                           n1777, ZN => n7091);
   U2570 : OAI22_X1 port map( A1 => n1775, A2 => n1779, B1 => n1152, B2 => 
                           n1777, ZN => n7092);
   U2571 : OAI22_X1 port map( A1 => n1775, A2 => n1780, B1 => n1154, B2 => 
                           n1777, ZN => n7093);
   U2572 : OAI22_X1 port map( A1 => n1775, A2 => n1781, B1 => n1156, B2 => 
                           n1777, ZN => n7094);
   U2573 : OAI22_X1 port map( A1 => n1775, A2 => n1782, B1 => n1158, B2 => 
                           n1777, ZN => n7095);
   U2574 : OAI22_X1 port map( A1 => n1775, A2 => n1783, B1 => n1160, B2 => 
                           n1777, ZN => n7096);
   U2575 : OAI22_X1 port map( A1 => n1775, A2 => n1784, B1 => n1162, B2 => 
                           n1777, ZN => n7097);
   U2576 : OAI22_X1 port map( A1 => n1775, A2 => n1785, B1 => n1164, B2 => 
                           n1777, ZN => n7098);
   U2577 : OAI22_X1 port map( A1 => n1775, A2 => n1786, B1 => n1166, B2 => 
                           n1777, ZN => n7099);
   U2578 : OAI22_X1 port map( A1 => n1775, A2 => n1787, B1 => n1168, B2 => 
                           n1777, ZN => n7100);
   U2579 : OAI22_X1 port map( A1 => n1775, A2 => n1788, B1 => n1170, B2 => 
                           n1777, ZN => n7101);
   U2580 : OAI22_X1 port map( A1 => n1775, A2 => n1789, B1 => n1172, B2 => 
                           n1777, ZN => n7102);
   U2582 : OAI22_X1 port map( A1 => n1775, A2 => n1791, B1 => n3529, B2 => 
                           n1777, ZN => n7104);
   U2583 : OAI22_X1 port map( A1 => n1775, A2 => n1792, B1 => n3529, B2 => 
                           n1777, ZN => n7105);
   U2585 : OAI22_X1 port map( A1 => n1775, A2 => n1794, B1 => n3529, B2 => 
                           n1777, ZN => n7107);
   U2586 : OAI22_X1 port map( A1 => n1775, A2 => n1795, B1 => n1179, B2 => 
                           n1777, ZN => n7108);
   U2587 : OAI22_X1 port map( A1 => n1775, A2 => n1796, B1 => n1181, B2 => 
                           n1777, ZN => n7109);
   U2588 : OAI22_X1 port map( A1 => n1775, A2 => n1797, B1 => n1183, B2 => 
                           n1777, ZN => n7110);
   U2589 : OAI22_X1 port map( A1 => n1775, A2 => n1798, B1 => n1185, B2 => 
                           n1777, ZN => n7111);
   U2590 : OAI22_X1 port map( A1 => n1775, A2 => n1799, B1 => n1187, B2 => 
                           n1777, ZN => n7112);
   U2591 : OAI22_X1 port map( A1 => n1775, A2 => n1800, B1 => n1189, B2 => 
                           n1777, ZN => n7113);
   U2592 : OAI22_X1 port map( A1 => n1775, A2 => n1801, B1 => n1191, B2 => 
                           n1777, ZN => n7114);
   U2593 : OAI22_X1 port map( A1 => n1775, A2 => n1802, B1 => n1193, B2 => 
                           n1777, ZN => n7115);
   U2594 : OAI22_X1 port map( A1 => n1775, A2 => n1803, B1 => n1195, B2 => 
                           n1777, ZN => n7116);
   U2595 : OAI22_X1 port map( A1 => n1775, A2 => n1804, B1 => n1197, B2 => 
                           n1777, ZN => n7117);
   U2596 : OAI22_X1 port map( A1 => n1775, A2 => n1805, B1 => n1199, B2 => 
                           n1777, ZN => n7118);
   U2597 : OAI22_X1 port map( A1 => n1775, A2 => n1806, B1 => n1201, B2 => 
                           n1777, ZN => n7119);
   U2598 : OAI22_X1 port map( A1 => n1775, A2 => n1807, B1 => n1203, B2 => 
                           n1777, ZN => n7120);
   U2599 : OAI22_X1 port map( A1 => n1775, A2 => n1808, B1 => n1205, B2 => 
                           n1777, ZN => n7121);
   U2602 : OAI22_X1 port map( A1 => n1809, A2 => n1810, B1 => n1147, B2 => 
                           n1811, ZN => n7122);
   U2603 : OAI22_X1 port map( A1 => n1809, A2 => n1812, B1 => n1150, B2 => 
                           n1811, ZN => n7123);
   U2604 : OAI22_X1 port map( A1 => n1809, A2 => n1813, B1 => n1152, B2 => 
                           n1811, ZN => n7124);
   U2605 : OAI22_X1 port map( A1 => n1809, A2 => n1814, B1 => n1154, B2 => 
                           n1811, ZN => n7125);
   U2606 : OAI22_X1 port map( A1 => n1809, A2 => n1815, B1 => n1156, B2 => 
                           n1811, ZN => n7126);
   U2607 : OAI22_X1 port map( A1 => n1809, A2 => n1816, B1 => n1158, B2 => 
                           n1811, ZN => n7127);
   U2608 : OAI22_X1 port map( A1 => n1809, A2 => n1817, B1 => n1160, B2 => 
                           n1811, ZN => n7128);
   U2609 : OAI22_X1 port map( A1 => n1809, A2 => n1818, B1 => n1162, B2 => 
                           n1811, ZN => n7129);
   U2610 : OAI22_X1 port map( A1 => n1809, A2 => n1819, B1 => n1164, B2 => 
                           n1811, ZN => n7130);
   U2611 : OAI22_X1 port map( A1 => n1809, A2 => n1820, B1 => n1166, B2 => 
                           n1811, ZN => n7131);
   U2612 : OAI22_X1 port map( A1 => n1809, A2 => n1821, B1 => n1168, B2 => 
                           n1811, ZN => n7132);
   U2613 : OAI22_X1 port map( A1 => n1809, A2 => n1822, B1 => n1170, B2 => 
                           n1811, ZN => n7133);
   U2614 : OAI22_X1 port map( A1 => n1809, A2 => n1823, B1 => n1172, B2 => 
                           n1811, ZN => n7134);
   U2616 : OAI22_X1 port map( A1 => n1809, A2 => n1825, B1 => n1496, B2 => 
                           n1811, ZN => n7136);
   U2619 : OAI22_X1 port map( A1 => n1809, A2 => n1828, B1 => n1496, B2 => 
                           n1811, ZN => n7139);
   U2620 : OAI22_X1 port map( A1 => n1809, A2 => n1829, B1 => n1179, B2 => 
                           n1811, ZN => n7140);
   U2621 : OAI22_X1 port map( A1 => n1809, A2 => n1830, B1 => n1181, B2 => 
                           n1811, ZN => n7141);
   U2622 : OAI22_X1 port map( A1 => n1809, A2 => n1831, B1 => n1183, B2 => 
                           n1811, ZN => n7142);
   U2623 : OAI22_X1 port map( A1 => n1809, A2 => n1832, B1 => n1185, B2 => 
                           n1811, ZN => n7143);
   U2624 : OAI22_X1 port map( A1 => n1809, A2 => n1833, B1 => n1187, B2 => 
                           n1811, ZN => n7144);
   U2625 : OAI22_X1 port map( A1 => n1809, A2 => n1834, B1 => n1189, B2 => 
                           n1811, ZN => n7145);
   U2626 : OAI22_X1 port map( A1 => n1809, A2 => n1835, B1 => n1191, B2 => 
                           n1811, ZN => n7146);
   U2627 : OAI22_X1 port map( A1 => n1809, A2 => n1836, B1 => n1193, B2 => 
                           n1811, ZN => n7147);
   U2628 : OAI22_X1 port map( A1 => n1809, A2 => n1837, B1 => n1195, B2 => 
                           n1811, ZN => n7148);
   U2629 : OAI22_X1 port map( A1 => n1809, A2 => n1838, B1 => n1197, B2 => 
                           n1811, ZN => n7149);
   U2630 : OAI22_X1 port map( A1 => n1809, A2 => n1839, B1 => n1199, B2 => 
                           n1811, ZN => n7150);
   U2631 : OAI22_X1 port map( A1 => n1809, A2 => n1840, B1 => n1201, B2 => 
                           n1811, ZN => n7151);
   U2632 : OAI22_X1 port map( A1 => n1809, A2 => n1841, B1 => n1203, B2 => 
                           n1811, ZN => n7152);
   U2633 : OAI22_X1 port map( A1 => n1809, A2 => n1842, B1 => n1205, B2 => 
                           n1811, ZN => n7153);
   U2637 : NOR2_X1 port map( A1 => n1844, A2 => n1845, ZN => n178);
   U2638 : OAI22_X1 port map( A1 => n1846, A2 => n1847, B1 => n1147, B2 => 
                           n3527, ZN => n7154);
   U2640 : OAI22_X1 port map( A1 => n1846, A2 => n1849, B1 => n1150, B2 => 
                           n3527, ZN => n7155);
   U2642 : OAI22_X1 port map( A1 => n1846, A2 => n1850, B1 => n1152, B2 => 
                           n3527, ZN => n7156);
   U2644 : OAI22_X1 port map( A1 => n1846, A2 => n1851, B1 => n1154, B2 => 
                           n3527, ZN => n7157);
   U2646 : OAI22_X1 port map( A1 => n1846, A2 => n1852, B1 => n1156, B2 => 
                           n3527, ZN => n7158);
   U2648 : OAI22_X1 port map( A1 => n1846, A2 => n1853, B1 => n1158, B2 => 
                           n3527, ZN => n7159);
   U2650 : OAI22_X1 port map( A1 => n1846, A2 => n1854, B1 => n1160, B2 => 
                           n3527, ZN => n7160);
   U2652 : OAI22_X1 port map( A1 => n1846, A2 => n1855, B1 => n1162, B2 => 
                           n3527, ZN => n7161);
   U2654 : OAI22_X1 port map( A1 => n1846, A2 => n1856, B1 => n1164, B2 => 
                           n3527, ZN => n7162);
   U2656 : OAI22_X1 port map( A1 => n1846, A2 => n1857, B1 => n1166, B2 => 
                           n3527, ZN => n7163);
   U2658 : OAI22_X1 port map( A1 => n1846, A2 => n1858, B1 => n1168, B2 => 
                           n3527, ZN => n7164);
   U2660 : OAI22_X1 port map( A1 => n1846, A2 => n1859, B1 => n1170, B2 => 
                           n3527, ZN => n7165);
   U2662 : OAI22_X1 port map( A1 => n1846, A2 => n1860, B1 => n1172, B2 => 
                           n3527, ZN => n7166);
   U2666 : INV_X1 port map( A => n1861, ZN => n7169);
   U2667 : AOI22_X1 port map( A1 => n3527, A2 => pc_lut_11_0_port, B1 => n3521,
                           B2 => n1846, ZN => n1861);
   U2668 : INV_X1 port map( A => n1862, ZN => n7170);
   U2669 : AOI22_X1 port map( A1 => n3527, A2 => pc_lut_11_1_port, B1 => n3521,
                           B2 => n1846, ZN => n1862);
   U2670 : INV_X1 port map( A => n1863, ZN => n7171);
   U2671 : AOI22_X1 port map( A1 => n3527, A2 => pc_lut_11_3_port, B1 => n3521,
                           B2 => n1846, ZN => n1863);
   U2672 : OAI22_X1 port map( A1 => n1846, A2 => n1864, B1 => n1179, B2 => 
                           n3527, ZN => n7172);
   U2674 : OAI22_X1 port map( A1 => n1846, A2 => n1865, B1 => n1181, B2 => 
                           n3527, ZN => n7173);
   U2676 : OAI22_X1 port map( A1 => n1846, A2 => n1866, B1 => n1183, B2 => 
                           n3527, ZN => n7174);
   U2678 : OAI22_X1 port map( A1 => n1846, A2 => n1867, B1 => n1185, B2 => 
                           n3527, ZN => n7175);
   U2680 : OAI22_X1 port map( A1 => n1846, A2 => n1868, B1 => n1187, B2 => 
                           n3527, ZN => n7176);
   U2682 : OAI22_X1 port map( A1 => n1846, A2 => n1869, B1 => n1189, B2 => 
                           n3527, ZN => n7177);
   U2684 : OAI22_X1 port map( A1 => n1846, A2 => n1870, B1 => n1191, B2 => 
                           n3527, ZN => n7178);
   U2686 : OAI22_X1 port map( A1 => n1846, A2 => n1871, B1 => n1193, B2 => 
                           n3527, ZN => n7179);
   U2688 : OAI22_X1 port map( A1 => n1846, A2 => n1872, B1 => n1195, B2 => 
                           n3527, ZN => n7180);
   U2690 : OAI22_X1 port map( A1 => n1846, A2 => n1873, B1 => n1197, B2 => 
                           n3527, ZN => n7181);
   U2692 : OAI22_X1 port map( A1 => n1846, A2 => n1874, B1 => n1199, B2 => 
                           n3527, ZN => n7182);
   U2694 : OAI22_X1 port map( A1 => n1846, A2 => n1875, B1 => n1201, B2 => 
                           n3527, ZN => n7183);
   U2696 : OAI22_X1 port map( A1 => n1846, A2 => n1876, B1 => n1203, B2 => 
                           n3527, ZN => n7184);
   U2698 : OAI22_X1 port map( A1 => n1846, A2 => n1877, B1 => n1205, B2 => 
                           n3527, ZN => n7185);
   U2701 : NAND2_X1 port map( A1 => n1878, A2 => n38, ZN => n1848);
   U2702 : OAI22_X1 port map( A1 => n1879, A2 => n1880, B1 => n1147, B2 => 
                           n1256, ZN => n7186);
   U2704 : OAI22_X1 port map( A1 => n1879, A2 => n1882, B1 => n1150, B2 => 
                           n1259, ZN => n7187);
   U2706 : OAI22_X1 port map( A1 => n1879, A2 => n1883, B1 => n1152, B2 => 
                           n1259, ZN => n7188);
   U2708 : OAI22_X1 port map( A1 => n1879, A2 => n1884, B1 => n1154, B2 => 
                           n1259, ZN => n7189);
   U2710 : OAI22_X1 port map( A1 => n1879, A2 => n1885, B1 => n1156, B2 => 
                           n1259, ZN => n7190);
   U2712 : OAI22_X1 port map( A1 => n1879, A2 => n1886, B1 => n1158, B2 => 
                           n1259, ZN => n7191);
   U2714 : OAI22_X1 port map( A1 => n1879, A2 => n1887, B1 => n1160, B2 => 
                           n1259, ZN => n7192);
   U2716 : OAI22_X1 port map( A1 => n1879, A2 => n1888, B1 => n1162, B2 => 
                           n1259, ZN => n7193);
   U2718 : OAI22_X1 port map( A1 => n1879, A2 => n1889, B1 => n1164, B2 => 
                           n1259, ZN => n7194);
   U2720 : OAI22_X1 port map( A1 => n1879, A2 => n1890, B1 => n1166, B2 => 
                           n1259, ZN => n7195);
   U2722 : OAI22_X1 port map( A1 => n1879, A2 => n1891, B1 => n1168, B2 => 
                           n1259, ZN => n7196);
   U2724 : OAI22_X1 port map( A1 => n1879, A2 => n1892, B1 => n1170, B2 => 
                           n1259, ZN => n7197);
   U2726 : OAI22_X1 port map( A1 => n1879, A2 => n1893, B1 => n1172, B2 => 
                           n1259, ZN => n7198);
   U2731 : INV_X1 port map( A => n1894, ZN => n7202);
   U2732 : AOI22_X1 port map( A1 => n1256, A2 => pc_lut_10_1_port, B1 => n3521,
                           B2 => n1879, ZN => n1894);
   U2733 : INV_X1 port map( A => n1895, ZN => n7203);
   U2734 : AOI22_X1 port map( A1 => n1256, A2 => pc_lut_10_3_port, B1 => n3521,
                           B2 => n1879, ZN => n1895);
   U2735 : OAI22_X1 port map( A1 => n1879, A2 => n1896, B1 => n1179, B2 => 
                           n1259, ZN => n7204);
   U2737 : OAI22_X1 port map( A1 => n1879, A2 => n1897, B1 => n1181, B2 => 
                           n1259, ZN => n7205);
   U2739 : OAI22_X1 port map( A1 => n1879, A2 => n1898, B1 => n1183, B2 => 
                           n1259, ZN => n7206);
   U2741 : OAI22_X1 port map( A1 => n1879, A2 => n1899, B1 => n1185, B2 => 
                           n1259, ZN => n7207);
   U2743 : OAI22_X1 port map( A1 => n1879, A2 => n1900, B1 => n1187, B2 => 
                           n1259, ZN => n7208);
   U2745 : OAI22_X1 port map( A1 => n1879, A2 => n1901, B1 => n1189, B2 => 
                           n1259, ZN => n7209);
   U2747 : OAI22_X1 port map( A1 => n1879, A2 => n1902, B1 => n1191, B2 => 
                           n1259, ZN => n7210);
   U2749 : OAI22_X1 port map( A1 => n1879, A2 => n1903, B1 => n1193, B2 => 
                           n1259, ZN => n7211);
   U2751 : OAI22_X1 port map( A1 => n1879, A2 => n1904, B1 => n1195, B2 => 
                           n1259, ZN => n7212);
   U2753 : OAI22_X1 port map( A1 => n1879, A2 => n1905, B1 => n1197, B2 => 
                           n1259, ZN => n7213);
   U2755 : OAI22_X1 port map( A1 => n1879, A2 => n1906, B1 => n1199, B2 => 
                           n1259, ZN => n7214);
   U2757 : OAI22_X1 port map( A1 => n1879, A2 => n1907, B1 => n1201, B2 => 
                           n1259, ZN => n7215);
   U2759 : OAI22_X1 port map( A1 => n1879, A2 => n1908, B1 => n1203, B2 => 
                           n1259, ZN => n7216);
   U2761 : OAI22_X1 port map( A1 => n1879, A2 => n1909, B1 => n1205, B2 => 
                           n1259, ZN => n7217);
   U2765 : OAI22_X1 port map( A1 => n1910, A2 => n1911, B1 => n1147, B2 => 
                           n1912, ZN => n7218);
   U2766 : OAI22_X1 port map( A1 => n1910, A2 => n1913, B1 => n1150, B2 => 
                           n1912, ZN => n7219);
   U2767 : OAI22_X1 port map( A1 => n1910, A2 => n1914, B1 => n1152, B2 => 
                           n1912, ZN => n7220);
   U2768 : OAI22_X1 port map( A1 => n1910, A2 => n1915, B1 => n1154, B2 => 
                           n1912, ZN => n7221);
   U2769 : OAI22_X1 port map( A1 => n1910, A2 => n1916, B1 => n1156, B2 => 
                           n1912, ZN => n7222);
   U2770 : OAI22_X1 port map( A1 => n1910, A2 => n1917, B1 => n1158, B2 => 
                           n1912, ZN => n7223);
   U2771 : OAI22_X1 port map( A1 => n1910, A2 => n1918, B1 => n1160, B2 => 
                           n1912, ZN => n7224);
   U2772 : OAI22_X1 port map( A1 => n1910, A2 => n1919, B1 => n1162, B2 => 
                           n1912, ZN => n7225);
   U2773 : OAI22_X1 port map( A1 => n1910, A2 => n1920, B1 => n1164, B2 => 
                           n1912, ZN => n7226);
   U2774 : OAI22_X1 port map( A1 => n1910, A2 => n1921, B1 => n1166, B2 => 
                           n1912, ZN => n7227);
   U2775 : OAI22_X1 port map( A1 => n1910, A2 => n1922, B1 => n1168, B2 => 
                           n1912, ZN => n7228);
   U2776 : OAI22_X1 port map( A1 => n1910, A2 => n1923, B1 => n1170, B2 => 
                           n1912, ZN => n7229);
   U2777 : OAI22_X1 port map( A1 => n1910, A2 => n1924, B1 => n1172, B2 => 
                           n1912, ZN => n7230);
   U2780 : OAI22_X1 port map( A1 => n1910, A2 => n1927, B1 => n1496, B2 => 
                           n1912, ZN => n7233);
   U2782 : OAI22_X1 port map( A1 => n1910, A2 => n1929, B1 => n1496, B2 => 
                           n1912, ZN => n7235);
   U2783 : OAI22_X1 port map( A1 => n1910, A2 => n1930, B1 => n1179, B2 => 
                           n1912, ZN => n7236);
   U2784 : OAI22_X1 port map( A1 => n1910, A2 => n1931, B1 => n1181, B2 => 
                           n1912, ZN => n7237);
   U2785 : OAI22_X1 port map( A1 => n1910, A2 => n1932, B1 => n1183, B2 => 
                           n1912, ZN => n7238);
   U2786 : OAI22_X1 port map( A1 => n1910, A2 => n1933, B1 => n1185, B2 => 
                           n1912, ZN => n7239);
   U2787 : OAI22_X1 port map( A1 => n1910, A2 => n1934, B1 => n1187, B2 => 
                           n1912, ZN => n7240);
   U2788 : OAI22_X1 port map( A1 => n1910, A2 => n1935, B1 => n1189, B2 => 
                           n1912, ZN => n7241);
   U2789 : OAI22_X1 port map( A1 => n1910, A2 => n1936, B1 => n1191, B2 => 
                           n1912, ZN => n7242);
   U2790 : OAI22_X1 port map( A1 => n1910, A2 => n1937, B1 => n1193, B2 => 
                           n1912, ZN => n7243);
   U2791 : OAI22_X1 port map( A1 => n1910, A2 => n1938, B1 => n1195, B2 => 
                           n1912, ZN => n7244);
   U2792 : OAI22_X1 port map( A1 => n1910, A2 => n1939, B1 => n1197, B2 => 
                           n1912, ZN => n7245);
   U2793 : OAI22_X1 port map( A1 => n1910, A2 => n1940, B1 => n1199, B2 => 
                           n1912, ZN => n7246);
   U2794 : OAI22_X1 port map( A1 => n1910, A2 => n1941, B1 => n1201, B2 => 
                           n1912, ZN => n7247);
   U2795 : OAI22_X1 port map( A1 => n1910, A2 => n1942, B1 => n1203, B2 => 
                           n1912, ZN => n7248);
   U2796 : OAI22_X1 port map( A1 => n1910, A2 => n1943, B1 => n1205, B2 => 
                           n1912, ZN => n7249);
   U2799 : OAI22_X1 port map( A1 => n1944, A2 => n1945, B1 => n1147, B2 => 
                           n1946, ZN => n7250);
   U2800 : OAI22_X1 port map( A1 => n1944, A2 => n1947, B1 => n1150, B2 => 
                           n1946, ZN => n7251);
   U2801 : OAI22_X1 port map( A1 => n1944, A2 => n1948, B1 => n1152, B2 => 
                           n1946, ZN => n7252);
   U2802 : OAI22_X1 port map( A1 => n1944, A2 => n1949, B1 => n1154, B2 => 
                           n1946, ZN => n7253);
   U2803 : OAI22_X1 port map( A1 => n1944, A2 => n1950, B1 => n1156, B2 => 
                           n1946, ZN => n7254);
   U2804 : OAI22_X1 port map( A1 => n1944, A2 => n1951, B1 => n1158, B2 => 
                           n1946, ZN => n7255);
   U2805 : OAI22_X1 port map( A1 => n1944, A2 => n1952, B1 => n1160, B2 => 
                           n1946, ZN => n7256);
   U2806 : OAI22_X1 port map( A1 => n1944, A2 => n1953, B1 => n1162, B2 => 
                           n1946, ZN => n7257);
   U2807 : OAI22_X1 port map( A1 => n1944, A2 => n1954, B1 => n1164, B2 => 
                           n1946, ZN => n7258);
   U2808 : OAI22_X1 port map( A1 => n1944, A2 => n1955, B1 => n1166, B2 => 
                           n1946, ZN => n7259);
   U2809 : OAI22_X1 port map( A1 => n1944, A2 => n1956, B1 => n1168, B2 => 
                           n1946, ZN => n7260);
   U2810 : OAI22_X1 port map( A1 => n1944, A2 => n1957, B1 => n1170, B2 => 
                           n1946, ZN => n7261);
   U2811 : OAI22_X1 port map( A1 => n1944, A2 => n1958, B1 => n1172, B2 => 
                           n1946, ZN => n7262);
   U2816 : OAI22_X1 port map( A1 => n1944, A2 => n1963, B1 => n1496, B2 => 
                           n1946, ZN => n7267);
   U2817 : OAI22_X1 port map( A1 => n1944, A2 => n1964, B1 => n1179, B2 => 
                           n1946, ZN => n7268);
   U2818 : OAI22_X1 port map( A1 => n1944, A2 => n1965, B1 => n1181, B2 => 
                           n1946, ZN => n7269);
   U2819 : OAI22_X1 port map( A1 => n1944, A2 => n1966, B1 => n1183, B2 => 
                           n1946, ZN => n7270);
   U2820 : OAI22_X1 port map( A1 => n1944, A2 => n1967, B1 => n1185, B2 => 
                           n1946, ZN => n7271);
   U2821 : OAI22_X1 port map( A1 => n1944, A2 => n1968, B1 => n1187, B2 => 
                           n1946, ZN => n7272);
   U2822 : OAI22_X1 port map( A1 => n1944, A2 => n1969, B1 => n1189, B2 => 
                           n1946, ZN => n7273);
   U2823 : OAI22_X1 port map( A1 => n1944, A2 => n1970, B1 => n1191, B2 => 
                           n1946, ZN => n7274);
   U2824 : OAI22_X1 port map( A1 => n1944, A2 => n1971, B1 => n1193, B2 => 
                           n1946, ZN => n7275);
   U2825 : OAI22_X1 port map( A1 => n1944, A2 => n1972, B1 => n1195, B2 => 
                           n1946, ZN => n7276);
   U2826 : OAI22_X1 port map( A1 => n1944, A2 => n1973, B1 => n1197, B2 => 
                           n1946, ZN => n7277);
   U2827 : OAI22_X1 port map( A1 => n1944, A2 => n1974, B1 => n1199, B2 => 
                           n1946, ZN => n7278);
   U2828 : OAI22_X1 port map( A1 => n1944, A2 => n1975, B1 => n1201, B2 => 
                           n1946, ZN => n7279);
   U2829 : OAI22_X1 port map( A1 => n1944, A2 => n1976, B1 => n1203, B2 => 
                           n1946, ZN => n7280);
   U2830 : OAI22_X1 port map( A1 => n1944, A2 => n1977, B1 => n1205, B2 => 
                           n1946, ZN => n7281);
   U2833 : AND2_X1 port map( A1 => n3794, A2 => n316, ZN => n1878);
   U2834 : NOR2_X1 port map( A1 => n1844, A2 => PC_write(2), ZN => n316);
   U2835 : INV_X1 port map( A => PC_write(3), ZN => n1844);
   U2836 : OAI22_X1 port map( A1 => n1978, A2 => n1979, B1 => n1147, B2 => 
                           n3524, ZN => n7282);
   U2838 : OAI22_X1 port map( A1 => n1978, A2 => n1981, B1 => n1150, B2 => 
                           n3524, ZN => n7283);
   U2840 : OAI22_X1 port map( A1 => n1978, A2 => n1982, B1 => n1152, B2 => 
                           n3524, ZN => n7284);
   U2842 : OAI22_X1 port map( A1 => n1978, A2 => n1983, B1 => n1154, B2 => 
                           n3524, ZN => n7285);
   U2844 : OAI22_X1 port map( A1 => n1978, A2 => n1984, B1 => n1156, B2 => 
                           n3524, ZN => n7286);
   U2846 : OAI22_X1 port map( A1 => n1978, A2 => n1985, B1 => n1158, B2 => 
                           n3524, ZN => n7287);
   U2848 : OAI22_X1 port map( A1 => n1978, A2 => n1986, B1 => n1160, B2 => 
                           n3524, ZN => n7288);
   U2850 : OAI22_X1 port map( A1 => n1978, A2 => n1987, B1 => n1162, B2 => 
                           n3524, ZN => n7289);
   U2852 : OAI22_X1 port map( A1 => n1978, A2 => n1988, B1 => n1164, B2 => 
                           n3524, ZN => n7290);
   U2854 : OAI22_X1 port map( A1 => n1978, A2 => n1989, B1 => n1166, B2 => 
                           n3524, ZN => n7291);
   U2856 : OAI22_X1 port map( A1 => n1978, A2 => n1990, B1 => n1168, B2 => 
                           n3524, ZN => n7292);
   U2858 : OAI22_X1 port map( A1 => n1978, A2 => n1991, B1 => n1170, B2 => 
                           n3524, ZN => n7293);
   U2860 : OAI22_X1 port map( A1 => n1978, A2 => n1992, B1 => n1172, B2 => 
                           n3524, ZN => n7294);
   U2863 : INV_X1 port map( A => n1993, ZN => n7296);
   U2864 : AOI22_X1 port map( A1 => n3524, A2 => pc_lut_7_2_port, B1 => n3521, 
                           B2 => n1978, ZN => n1993);
   U2865 : INV_X1 port map( A => n1994, ZN => n7297);
   U2866 : AOI22_X1 port map( A1 => n3524, A2 => pc_lut_7_0_port, B1 => n3521, 
                           B2 => n1978, ZN => n1994);
   U2867 : INV_X1 port map( A => n1995, ZN => n7298);
   U2868 : AOI22_X1 port map( A1 => n3524, A2 => pc_lut_7_1_port, B1 => n3521, 
                           B2 => n1978, ZN => n1995);
   U2870 : OAI22_X1 port map( A1 => n1978, A2 => n1996, B1 => n1179, B2 => 
                           n3524, ZN => n7300);
   U2872 : OAI22_X1 port map( A1 => n1978, A2 => n1997, B1 => n1181, B2 => 
                           n3524, ZN => n7301);
   U2874 : OAI22_X1 port map( A1 => n1978, A2 => n1998, B1 => n1183, B2 => 
                           n3524, ZN => n7302);
   U2876 : OAI22_X1 port map( A1 => n1978, A2 => n1999, B1 => n1185, B2 => 
                           n3524, ZN => n7303);
   U2878 : OAI22_X1 port map( A1 => n1978, A2 => n2000, B1 => n1187, B2 => 
                           n3524, ZN => n7304);
   U2880 : OAI22_X1 port map( A1 => n1978, A2 => n2001, B1 => n1189, B2 => 
                           n3524, ZN => n7305);
   U2882 : OAI22_X1 port map( A1 => n1978, A2 => n2002, B1 => n1191, B2 => 
                           n3524, ZN => n7306);
   U2884 : OAI22_X1 port map( A1 => n1978, A2 => n2003, B1 => n1193, B2 => 
                           n3524, ZN => n7307);
   U2886 : OAI22_X1 port map( A1 => n1978, A2 => n2004, B1 => n1195, B2 => 
                           n3524, ZN => n7308);
   U2888 : OAI22_X1 port map( A1 => n1978, A2 => n2005, B1 => n1197, B2 => 
                           n3524, ZN => n7309);
   U2890 : OAI22_X1 port map( A1 => n1978, A2 => n2006, B1 => n1199, B2 => 
                           n3524, ZN => n7310);
   U2892 : OAI22_X1 port map( A1 => n1978, A2 => n2007, B1 => n1201, B2 => 
                           n3524, ZN => n7311);
   U2894 : OAI22_X1 port map( A1 => n1978, A2 => n2008, B1 => n1203, B2 => 
                           n3524, ZN => n7312);
   U2896 : OAI22_X1 port map( A1 => n1978, A2 => n2009, B1 => n1205, B2 => 
                           n3524, ZN => n7313);
   U2899 : NAND2_X1 port map( A1 => n2010, A2 => n38, ZN => n1980);
   U2900 : OAI22_X1 port map( A1 => n2011, A2 => n2012, B1 => n1147, B2 => 
                           n1292, ZN => n7314);
   U2902 : OAI22_X1 port map( A1 => n2011, A2 => n2014, B1 => n1150, B2 => 
                           n1293, ZN => n7315);
   U2904 : OAI22_X1 port map( A1 => n2011, A2 => n2015, B1 => n1152, B2 => 
                           n1293, ZN => n7316);
   U2906 : OAI22_X1 port map( A1 => n2011, A2 => n2016, B1 => n1154, B2 => 
                           n1293, ZN => n7317);
   U2908 : OAI22_X1 port map( A1 => n2011, A2 => n2017, B1 => n1156, B2 => 
                           n1293, ZN => n7318);
   U2910 : OAI22_X1 port map( A1 => n2011, A2 => n2018, B1 => n1158, B2 => 
                           n1293, ZN => n7319);
   U2912 : OAI22_X1 port map( A1 => n2011, A2 => n2019, B1 => n1160, B2 => 
                           n1293, ZN => n7320);
   U2914 : OAI22_X1 port map( A1 => n2011, A2 => n2020, B1 => n1162, B2 => 
                           n1293, ZN => n7321);
   U2916 : OAI22_X1 port map( A1 => n2011, A2 => n2021, B1 => n1164, B2 => 
                           n1293, ZN => n7322);
   U2918 : OAI22_X1 port map( A1 => n2011, A2 => n2022, B1 => n1166, B2 => 
                           n1293, ZN => n7323);
   U2920 : OAI22_X1 port map( A1 => n2011, A2 => n2023, B1 => n1168, B2 => 
                           n1293, ZN => n7324);
   U2922 : OAI22_X1 port map( A1 => n2011, A2 => n2024, B1 => n1170, B2 => 
                           n1293, ZN => n7325);
   U2924 : OAI22_X1 port map( A1 => n2011, A2 => n2025, B1 => n1172, B2 => 
                           n1293, ZN => n7326);
   U2927 : INV_X1 port map( A => n2026, ZN => n7328);
   U2928 : AOI22_X1 port map( A1 => n1292, A2 => pc_lut_6_2_port, B1 => n3521, 
                           B2 => n2011, ZN => n2026);
   U2930 : INV_X1 port map( A => n2027, ZN => n7330);
   U2931 : AOI22_X1 port map( A1 => n1292, A2 => pc_lut_6_1_port, B1 => n3521, 
                           B2 => n2011, ZN => n2027);
   U2933 : OAI22_X1 port map( A1 => n2011, A2 => n2028, B1 => n1179, B2 => 
                           n1293, ZN => n7332);
   U2935 : OAI22_X1 port map( A1 => n2011, A2 => n2029, B1 => n1181, B2 => 
                           n1293, ZN => n7333);
   U2937 : OAI22_X1 port map( A1 => n2011, A2 => n2030, B1 => n1183, B2 => 
                           n1293, ZN => n7334);
   U2939 : OAI22_X1 port map( A1 => n2011, A2 => n2031, B1 => n1185, B2 => 
                           n1293, ZN => n7335);
   U2941 : OAI22_X1 port map( A1 => n2011, A2 => n2032, B1 => n1187, B2 => 
                           n1293, ZN => n7336);
   U2943 : OAI22_X1 port map( A1 => n2011, A2 => n2033, B1 => n1189, B2 => 
                           n1293, ZN => n7337);
   U2945 : OAI22_X1 port map( A1 => n2011, A2 => n2034, B1 => n1191, B2 => 
                           n1293, ZN => n7338);
   U2947 : OAI22_X1 port map( A1 => n2011, A2 => n2035, B1 => n1193, B2 => 
                           n1293, ZN => n7339);
   U2949 : OAI22_X1 port map( A1 => n2011, A2 => n2036, B1 => n1195, B2 => 
                           n1293, ZN => n7340);
   U2951 : OAI22_X1 port map( A1 => n2011, A2 => n2037, B1 => n1197, B2 => 
                           n1293, ZN => n7341);
   U2953 : OAI22_X1 port map( A1 => n2011, A2 => n2038, B1 => n1199, B2 => 
                           n1293, ZN => n7342);
   U2955 : OAI22_X1 port map( A1 => n2011, A2 => n2039, B1 => n1201, B2 => 
                           n1293, ZN => n7343);
   U2957 : OAI22_X1 port map( A1 => n2011, A2 => n2040, B1 => n1203, B2 => 
                           n1293, ZN => n7344);
   U2959 : OAI22_X1 port map( A1 => n2011, A2 => n2041, B1 => n1205, B2 => 
                           n1293, ZN => n7345);
   U2963 : OAI22_X1 port map( A1 => n2042, A2 => n2043, B1 => n1147, B2 => 
                           n2044, ZN => n7346);
   U2964 : OAI22_X1 port map( A1 => n2042, A2 => n2045, B1 => n1150, B2 => 
                           n2044, ZN => n7347);
   U2965 : OAI22_X1 port map( A1 => n2042, A2 => n2046, B1 => n1152, B2 => 
                           n2044, ZN => n7348);
   U2966 : OAI22_X1 port map( A1 => n2042, A2 => n2047, B1 => n1154, B2 => 
                           n2044, ZN => n7349);
   U2967 : OAI22_X1 port map( A1 => n2042, A2 => n2048, B1 => n1156, B2 => 
                           n2044, ZN => n7350);
   U2968 : OAI22_X1 port map( A1 => n2042, A2 => n2049, B1 => n1158, B2 => 
                           n2044, ZN => n7351);
   U2969 : OAI22_X1 port map( A1 => n2042, A2 => n2050, B1 => n1160, B2 => 
                           n2044, ZN => n7352);
   U2970 : OAI22_X1 port map( A1 => n2042, A2 => n2051, B1 => n1162, B2 => 
                           n2044, ZN => n7353);
   U2971 : OAI22_X1 port map( A1 => n2042, A2 => n2052, B1 => n1164, B2 => 
                           n2044, ZN => n7354);
   U2972 : OAI22_X1 port map( A1 => n2042, A2 => n2053, B1 => n1166, B2 => 
                           n2044, ZN => n7355);
   U2973 : OAI22_X1 port map( A1 => n2042, A2 => n2054, B1 => n1168, B2 => 
                           n2044, ZN => n7356);
   U2974 : OAI22_X1 port map( A1 => n2042, A2 => n2055, B1 => n1170, B2 => 
                           n2044, ZN => n7357);
   U2975 : OAI22_X1 port map( A1 => n2042, A2 => n2056, B1 => n1172, B2 => 
                           n2044, ZN => n7358);
   U2977 : OAI22_X1 port map( A1 => n2042, A2 => n2058, B1 => n1496, B2 => 
                           n2044, ZN => n7360);
   U2978 : OAI22_X1 port map( A1 => n2042, A2 => n2059, B1 => n1496, B2 => 
                           n2044, ZN => n7361);
   U2981 : OAI22_X1 port map( A1 => n2042, A2 => n2062, B1 => n1179, B2 => 
                           n2044, ZN => n7364);
   U2982 : OAI22_X1 port map( A1 => n2042, A2 => n2063, B1 => n1181, B2 => 
                           n2044, ZN => n7365);
   U2983 : OAI22_X1 port map( A1 => n2042, A2 => n2064, B1 => n1183, B2 => 
                           n2044, ZN => n7366);
   U2984 : OAI22_X1 port map( A1 => n2042, A2 => n2065, B1 => n1185, B2 => 
                           n2044, ZN => n7367);
   U2985 : OAI22_X1 port map( A1 => n2042, A2 => n2066, B1 => n1187, B2 => 
                           n2044, ZN => n7368);
   U2986 : OAI22_X1 port map( A1 => n2042, A2 => n2067, B1 => n1189, B2 => 
                           n2044, ZN => n7369);
   U2987 : OAI22_X1 port map( A1 => n2042, A2 => n2068, B1 => n1191, B2 => 
                           n2044, ZN => n7370);
   U2988 : OAI22_X1 port map( A1 => n2042, A2 => n2069, B1 => n1193, B2 => 
                           n2044, ZN => n7371);
   U2989 : OAI22_X1 port map( A1 => n2042, A2 => n2070, B1 => n1195, B2 => 
                           n2044, ZN => n7372);
   U2990 : OAI22_X1 port map( A1 => n2042, A2 => n2071, B1 => n1197, B2 => 
                           n2044, ZN => n7373);
   U2991 : OAI22_X1 port map( A1 => n2042, A2 => n2072, B1 => n1199, B2 => 
                           n2044, ZN => n7374);
   U2992 : OAI22_X1 port map( A1 => n2042, A2 => n2073, B1 => n1201, B2 => 
                           n2044, ZN => n7375);
   U2993 : OAI22_X1 port map( A1 => n2042, A2 => n2074, B1 => n1203, B2 => 
                           n2044, ZN => n7376);
   U2994 : OAI22_X1 port map( A1 => n2042, A2 => n2075, B1 => n1205, B2 => 
                           n2044, ZN => n7377);
   U2997 : OAI22_X1 port map( A1 => n2076, A2 => n2077, B1 => n1147, B2 => 
                           n2078, ZN => n7378);
   U2998 : OAI22_X1 port map( A1 => n2076, A2 => n2079, B1 => n1150, B2 => 
                           n2078, ZN => n7379);
   U2999 : OAI22_X1 port map( A1 => n2076, A2 => n2080, B1 => n1152, B2 => 
                           n2078, ZN => n7380);
   U3000 : OAI22_X1 port map( A1 => n2076, A2 => n2081, B1 => n1154, B2 => 
                           n2078, ZN => n7381);
   U3001 : OAI22_X1 port map( A1 => n2076, A2 => n2082, B1 => n1156, B2 => 
                           n2078, ZN => n7382);
   U3002 : OAI22_X1 port map( A1 => n2076, A2 => n2083, B1 => n1158, B2 => 
                           n2078, ZN => n7383);
   U3003 : OAI22_X1 port map( A1 => n2076, A2 => n2084, B1 => n1160, B2 => 
                           n2078, ZN => n7384);
   U3004 : OAI22_X1 port map( A1 => n2076, A2 => n2085, B1 => n1162, B2 => 
                           n2078, ZN => n7385);
   U3005 : OAI22_X1 port map( A1 => n2076, A2 => n2086, B1 => n1164, B2 => 
                           n2078, ZN => n7386);
   U3006 : OAI22_X1 port map( A1 => n2076, A2 => n2087, B1 => n1166, B2 => 
                           n2078, ZN => n7387);
   U3007 : OAI22_X1 port map( A1 => n2076, A2 => n2088, B1 => n1168, B2 => 
                           n2078, ZN => n7388);
   U3008 : OAI22_X1 port map( A1 => n2076, A2 => n2089, B1 => n1170, B2 => 
                           n2078, ZN => n7389);
   U3009 : OAI22_X1 port map( A1 => n2076, A2 => n2090, B1 => n1172, B2 => 
                           n2078, ZN => n7390);
   U3011 : OAI22_X1 port map( A1 => n2076, A2 => n2092, B1 => n1496, B2 => 
                           n2078, ZN => n7392);
   U3015 : OAI22_X1 port map( A1 => n2076, A2 => n2096, B1 => n1179, B2 => 
                           n2078, ZN => n7396);
   U3016 : OAI22_X1 port map( A1 => n2076, A2 => n2097, B1 => n1181, B2 => 
                           n2078, ZN => n7397);
   U3017 : OAI22_X1 port map( A1 => n2076, A2 => n2098, B1 => n1183, B2 => 
                           n2078, ZN => n7398);
   U3018 : OAI22_X1 port map( A1 => n2076, A2 => n2099, B1 => n1185, B2 => 
                           n2078, ZN => n7399);
   U3019 : OAI22_X1 port map( A1 => n2076, A2 => n2100, B1 => n1187, B2 => 
                           n2078, ZN => n7400);
   U3020 : OAI22_X1 port map( A1 => n2076, A2 => n2101, B1 => n1189, B2 => 
                           n2078, ZN => n7401);
   U3021 : OAI22_X1 port map( A1 => n2076, A2 => n2102, B1 => n1191, B2 => 
                           n2078, ZN => n7402);
   U3022 : OAI22_X1 port map( A1 => n2076, A2 => n2103, B1 => n1193, B2 => 
                           n2078, ZN => n7403);
   U3023 : OAI22_X1 port map( A1 => n2076, A2 => n2104, B1 => n1195, B2 => 
                           n2078, ZN => n7404);
   U3024 : OAI22_X1 port map( A1 => n2076, A2 => n2105, B1 => n1197, B2 => 
                           n2078, ZN => n7405);
   U3025 : OAI22_X1 port map( A1 => n2076, A2 => n2106, B1 => n1199, B2 => 
                           n2078, ZN => n7406);
   U3026 : OAI22_X1 port map( A1 => n2076, A2 => n2107, B1 => n1201, B2 => 
                           n2078, ZN => n7407);
   U3027 : OAI22_X1 port map( A1 => n2076, A2 => n2108, B1 => n1203, B2 => 
                           n2078, ZN => n7408);
   U3028 : OAI22_X1 port map( A1 => n2076, A2 => n2109, B1 => n1205, B2 => 
                           n2078, ZN => n7409);
   U3031 : AND2_X1 port map( A1 => n1843, A2 => n454, ZN => n2010);
   U3032 : NOR2_X1 port map( A1 => n1845, A2 => PC_write(3), ZN => n454);
   U3033 : INV_X1 port map( A => PC_write(2), ZN => n1845);
   U3034 : OAI22_X1 port map( A1 => n2110, A2 => n2111, B1 => n1147, B2 => n871
                           , ZN => n7410);
   U3036 : OAI22_X1 port map( A1 => n2110, A2 => n2113, B1 => n1150, B2 => n973
                           , ZN => n7411);
   U3038 : OAI22_X1 port map( A1 => n2110, A2 => n2114, B1 => n1152, B2 => n973
                           , ZN => n7412);
   U3040 : OAI22_X1 port map( A1 => n2110, A2 => n2115, B1 => n1154, B2 => n973
                           , ZN => n7413);
   U3042 : OAI22_X1 port map( A1 => n2110, A2 => n2116, B1 => n1156, B2 => n973
                           , ZN => n7414);
   U3044 : OAI22_X1 port map( A1 => n2110, A2 => n2117, B1 => n1158, B2 => n973
                           , ZN => n7415);
   U3046 : OAI22_X1 port map( A1 => n2110, A2 => n2118, B1 => n1160, B2 => n973
                           , ZN => n7416);
   U3048 : OAI22_X1 port map( A1 => n2110, A2 => n2119, B1 => n1162, B2 => n973
                           , ZN => n7417);
   U3050 : OAI22_X1 port map( A1 => n2110, A2 => n2120, B1 => n1164, B2 => n973
                           , ZN => n7418);
   U3052 : OAI22_X1 port map( A1 => n2110, A2 => n2121, B1 => n1166, B2 => n973
                           , ZN => n7419);
   U3054 : OAI22_X1 port map( A1 => n2110, A2 => n2122, B1 => n1168, B2 => n973
                           , ZN => n7420);
   U3056 : OAI22_X1 port map( A1 => n2110, A2 => n2123, B1 => n1170, B2 => n973
                           , ZN => n7421);
   U3058 : OAI22_X1 port map( A1 => n2110, A2 => n2124, B1 => n1172, B2 => n973
                           , ZN => n7422);
   U3062 : INV_X1 port map( A => n2125, ZN => n7425);
   U3063 : AOI22_X1 port map( A1 => n871, A2 => pc_lut_3_0_port, B1 => n3521, 
                           B2 => n2110, ZN => n2125);
   U3064 : INV_X1 port map( A => n2126, ZN => n7426);
   U3065 : AOI22_X1 port map( A1 => n871, A2 => pc_lut_3_1_port, B1 => n3521, 
                           B2 => n2110, ZN => n2126);
   U3067 : OAI22_X1 port map( A1 => n2110, A2 => n2127, B1 => n1179, B2 => n973
                           , ZN => n7428);
   U3069 : OAI22_X1 port map( A1 => n2110, A2 => n2128, B1 => n1181, B2 => n973
                           , ZN => n7429);
   U3071 : OAI22_X1 port map( A1 => n2110, A2 => n2129, B1 => n1183, B2 => n973
                           , ZN => n7430);
   U3073 : OAI22_X1 port map( A1 => n2110, A2 => n2130, B1 => n1185, B2 => n973
                           , ZN => n7431);
   U3075 : OAI22_X1 port map( A1 => n2110, A2 => n2131, B1 => n1187, B2 => n973
                           , ZN => n7432);
   U3077 : OAI22_X1 port map( A1 => n2110, A2 => n2132, B1 => n1189, B2 => n973
                           , ZN => n7433);
   U3079 : OAI22_X1 port map( A1 => n2110, A2 => n2133, B1 => n1191, B2 => n973
                           , ZN => n7434);
   U3081 : OAI22_X1 port map( A1 => n2110, A2 => n2134, B1 => n1193, B2 => n973
                           , ZN => n7435);
   U3083 : OAI22_X1 port map( A1 => n2110, A2 => n2135, B1 => n1195, B2 => n973
                           , ZN => n7436);
   U3085 : OAI22_X1 port map( A1 => n2110, A2 => n2136, B1 => n1197, B2 => n973
                           , ZN => n7437);
   U3087 : OAI22_X1 port map( A1 => n2110, A2 => n2137, B1 => n1199, B2 => n973
                           , ZN => n7438);
   U3089 : OAI22_X1 port map( A1 => n2110, A2 => n2138, B1 => n1201, B2 => n973
                           , ZN => n7439);
   U3091 : OAI22_X1 port map( A1 => n2110, A2 => n2139, B1 => n1203, B2 => n973
                           , ZN => n7440);
   U3093 : OAI22_X1 port map( A1 => n2110, A2 => n2140, B1 => n1205, B2 => n973
                           , ZN => n7441);
   U3098 : OAI22_X1 port map( A1 => n2144, A2 => n2145, B1 => n1147, B2 => n3, 
                           ZN => n7442);
   U3100 : OAI22_X1 port map( A1 => n2144, A2 => n2147, B1 => n1150, B2 => n283
                           , ZN => n7443);
   U3102 : OAI22_X1 port map( A1 => n2144, A2 => n2148, B1 => n1152, B2 => n283
                           , ZN => n7444);
   U3104 : OAI22_X1 port map( A1 => n2144, A2 => n2149, B1 => n1154, B2 => n283
                           , ZN => n7445);
   U3106 : OAI22_X1 port map( A1 => n2144, A2 => n2150, B1 => n1156, B2 => n283
                           , ZN => n7446);
   U3108 : OAI22_X1 port map( A1 => n2144, A2 => n2151, B1 => n1158, B2 => n283
                           , ZN => n7447);
   U3110 : OAI22_X1 port map( A1 => n2144, A2 => n2152, B1 => n1160, B2 => n283
                           , ZN => n7448);
   U3112 : OAI22_X1 port map( A1 => n2144, A2 => n2153, B1 => n1162, B2 => n283
                           , ZN => n7449);
   U3114 : OAI22_X1 port map( A1 => n2144, A2 => n2154, B1 => n1164, B2 => n283
                           , ZN => n7450);
   U3116 : OAI22_X1 port map( A1 => n2144, A2 => n2155, B1 => n1166, B2 => n283
                           , ZN => n7451);
   U3118 : OAI22_X1 port map( A1 => n2144, A2 => n2156, B1 => n1168, B2 => n283
                           , ZN => n7452);
   U3120 : OAI22_X1 port map( A1 => n2144, A2 => n2157, B1 => n1170, B2 => n283
                           , ZN => n7453);
   U3122 : OAI22_X1 port map( A1 => n2144, A2 => n2158, B1 => n1172, B2 => n283
                           , ZN => n7454);
   U3127 : INV_X1 port map( A => n2159, ZN => n7458);
   U3128 : AOI22_X1 port map( A1 => n3, A2 => pc_lut_2_1_port, B1 => n3521, B2 
                           => n2144, ZN => n2159);
   U3130 : OAI22_X1 port map( A1 => n2144, A2 => n2160, B1 => n1179, B2 => n283
                           , ZN => n7460);
   U3132 : OAI22_X1 port map( A1 => n2144, A2 => n2161, B1 => n1181, B2 => n283
                           , ZN => n7461);
   U3134 : OAI22_X1 port map( A1 => n2144, A2 => n2162, B1 => n1183, B2 => n283
                           , ZN => n7462);
   U3136 : OAI22_X1 port map( A1 => n2144, A2 => n2163, B1 => n1185, B2 => n283
                           , ZN => n7463);
   U3138 : OAI22_X1 port map( A1 => n2144, A2 => n2164, B1 => n1187, B2 => n283
                           , ZN => n7464);
   U3140 : OAI22_X1 port map( A1 => n2144, A2 => n2165, B1 => n1189, B2 => n283
                           , ZN => n7465);
   U3142 : OAI22_X1 port map( A1 => n2144, A2 => n2166, B1 => n1191, B2 => n283
                           , ZN => n7466);
   U3144 : OAI22_X1 port map( A1 => n2144, A2 => n2167, B1 => n1193, B2 => n283
                           , ZN => n7467);
   U3146 : OAI22_X1 port map( A1 => n2144, A2 => n2168, B1 => n1195, B2 => n283
                           , ZN => n7468);
   U3148 : OAI22_X1 port map( A1 => n2144, A2 => n2169, B1 => n1197, B2 => n283
                           , ZN => n7469);
   U3150 : OAI22_X1 port map( A1 => n2144, A2 => n2170, B1 => n1199, B2 => n283
                           , ZN => n7470);
   U3152 : OAI22_X1 port map( A1 => n2144, A2 => n2171, B1 => n1201, B2 => n283
                           , ZN => n7471);
   U3154 : OAI22_X1 port map( A1 => n2144, A2 => n2172, B1 => n1203, B2 => n283
                           , ZN => n7472);
   U3156 : OAI22_X1 port map( A1 => n2144, A2 => n2173, B1 => n1205, B2 => n283
                           , ZN => n7473);
   U3161 : INV_X1 port map( A => PC_write(1), ZN => n2142);
   U3162 : OAI22_X1 port map( A1 => n2174, A2 => n2175, B1 => n1147, B2 => 
                           n2176, ZN => n7474);
   U3163 : OAI22_X1 port map( A1 => n2174, A2 => n2177, B1 => n1150, B2 => 
                           n2176, ZN => n7475);
   U3164 : OAI22_X1 port map( A1 => n2174, A2 => n2178, B1 => n1152, B2 => 
                           n2176, ZN => n7476);
   U3165 : OAI22_X1 port map( A1 => n2174, A2 => n2179, B1 => n1154, B2 => 
                           n2176, ZN => n7477);
   U3166 : OAI22_X1 port map( A1 => n2174, A2 => n2180, B1 => n1156, B2 => 
                           n2176, ZN => n7478);
   U3167 : OAI22_X1 port map( A1 => n2174, A2 => n2181, B1 => n1158, B2 => 
                           n2176, ZN => n7479);
   U3168 : OAI22_X1 port map( A1 => n2174, A2 => n2182, B1 => n1160, B2 => 
                           n2176, ZN => n7480);
   U3169 : OAI22_X1 port map( A1 => n2174, A2 => n2183, B1 => n1162, B2 => 
                           n2176, ZN => n7481);
   U3170 : OAI22_X1 port map( A1 => n2174, A2 => n2184, B1 => n1164, B2 => 
                           n2176, ZN => n7482);
   U3171 : OAI22_X1 port map( A1 => n2174, A2 => n2185, B1 => n1166, B2 => 
                           n2176, ZN => n7483);
   U3172 : OAI22_X1 port map( A1 => n2174, A2 => n2186, B1 => n1168, B2 => 
                           n2176, ZN => n7484);
   U3173 : OAI22_X1 port map( A1 => n2174, A2 => n2187, B1 => n1170, B2 => 
                           n2176, ZN => n7485);
   U3174 : OAI22_X1 port map( A1 => n2174, A2 => n2188, B1 => n1172, B2 => 
                           n2176, ZN => n7486);
   U3177 : OAI22_X1 port map( A1 => n2174, A2 => n2191, B1 => n1496, B2 => 
                           n2176, ZN => n7489);
   U3180 : OAI22_X1 port map( A1 => n2174, A2 => n2194, B1 => n1179, B2 => 
                           n2176, ZN => n7492);
   U3181 : OAI22_X1 port map( A1 => n2174, A2 => n2195, B1 => n1181, B2 => 
                           n2176, ZN => n7493);
   U3182 : OAI22_X1 port map( A1 => n2174, A2 => n2196, B1 => n1183, B2 => 
                           n2176, ZN => n7494);
   U3183 : OAI22_X1 port map( A1 => n2174, A2 => n2197, B1 => n1185, B2 => 
                           n2176, ZN => n7495);
   U3184 : OAI22_X1 port map( A1 => n2174, A2 => n2198, B1 => n1187, B2 => 
                           n2176, ZN => n7496);
   U3185 : OAI22_X1 port map( A1 => n2174, A2 => n2199, B1 => n1189, B2 => 
                           n2176, ZN => n7497);
   U3186 : OAI22_X1 port map( A1 => n2174, A2 => n2200, B1 => n1191, B2 => 
                           n2176, ZN => n7498);
   U3187 : OAI22_X1 port map( A1 => n2174, A2 => n2201, B1 => n1193, B2 => 
                           n2176, ZN => n7499);
   U3188 : OAI22_X1 port map( A1 => n2174, A2 => n2202, B1 => n1195, B2 => 
                           n2176, ZN => n7500);
   U3189 : OAI22_X1 port map( A1 => n2174, A2 => n2203, B1 => n1197, B2 => 
                           n2176, ZN => n7501);
   U3190 : OAI22_X1 port map( A1 => n2174, A2 => n2204, B1 => n1199, B2 => 
                           n2176, ZN => n7502);
   U3191 : OAI22_X1 port map( A1 => n2174, A2 => n2205, B1 => n1201, B2 => 
                           n2176, ZN => n7503);
   U3192 : OAI22_X1 port map( A1 => n2174, A2 => n2206, B1 => n1203, B2 => 
                           n2176, ZN => n7504);
   U3193 : OAI22_X1 port map( A1 => n2174, A2 => n2207, B1 => n1205, B2 => 
                           n2176, ZN => n7505);
   U3197 : INV_X1 port map( A => PC_write(0), ZN => n2143);
   U3198 : OAI22_X1 port map( A1 => n2208, A2 => n2209, B1 => n1147, B2 => 
                           n2210, ZN => n7506);
   U3200 : OAI22_X1 port map( A1 => n2208, A2 => n2211, B1 => n1150, B2 => 
                           n2210, ZN => n7507);
   U3202 : OAI22_X1 port map( A1 => n2208, A2 => n2212, B1 => n1152, B2 => 
                           n2210, ZN => n7508);
   U3204 : OAI22_X1 port map( A1 => n2208, A2 => n2213, B1 => n1154, B2 => 
                           n2210, ZN => n7509);
   U3206 : OAI22_X1 port map( A1 => n2208, A2 => n2214, B1 => n1156, B2 => 
                           n2210, ZN => n7510);
   U3208 : OAI22_X1 port map( A1 => n2208, A2 => n2215, B1 => n1158, B2 => 
                           n2210, ZN => n7511);
   U3210 : OAI22_X1 port map( A1 => n2208, A2 => n2216, B1 => n1160, B2 => 
                           n2210, ZN => n7512);
   U3212 : OAI22_X1 port map( A1 => n2208, A2 => n2217, B1 => n1162, B2 => 
                           n2210, ZN => n7513);
   U3214 : OAI22_X1 port map( A1 => n2208, A2 => n2218, B1 => n1164, B2 => 
                           n2210, ZN => n7514);
   U3216 : OAI22_X1 port map( A1 => n2208, A2 => n2219, B1 => n1166, B2 => 
                           n2210, ZN => n7515);
   U3218 : OAI22_X1 port map( A1 => n2208, A2 => n2220, B1 => n1168, B2 => 
                           n2210, ZN => n7516);
   U3220 : OAI22_X1 port map( A1 => n2208, A2 => n2221, B1 => n1170, B2 => 
                           n2210, ZN => n7517);
   U3222 : OAI22_X1 port map( A1 => n2208, A2 => n2222, B1 => n1172, B2 => 
                           n2210, ZN => n7518);
   U3229 : OAI22_X1 port map( A1 => n2208, A2 => n2228, B1 => n1179, B2 => 
                           n2210, ZN => n7524);
   U3231 : OAI22_X1 port map( A1 => n2208, A2 => n2229, B1 => n1181, B2 => 
                           n2210, ZN => n7525);
   U3233 : OAI22_X1 port map( A1 => n2208, A2 => n2230, B1 => n1183, B2 => 
                           n2210, ZN => n7526);
   U3235 : OAI22_X1 port map( A1 => n2208, A2 => n2231, B1 => n1185, B2 => 
                           n2210, ZN => n7527);
   U3237 : OAI22_X1 port map( A1 => n2208, A2 => n2232, B1 => n1187, B2 => 
                           n2210, ZN => n7528);
   U3239 : OAI22_X1 port map( A1 => n2208, A2 => n2233, B1 => n1189, B2 => 
                           n2210, ZN => n7529);
   U3241 : OAI22_X1 port map( A1 => n2208, A2 => n2234, B1 => n1191, B2 => 
                           n2210, ZN => n7530);
   U3243 : OAI22_X1 port map( A1 => n2208, A2 => n2235, B1 => n1193, B2 => 
                           n2210, ZN => n7531);
   U3245 : OAI22_X1 port map( A1 => n2208, A2 => n2236, B1 => n1195, B2 => 
                           n2210, ZN => n7532);
   U3247 : OAI22_X1 port map( A1 => n2208, A2 => n2237, B1 => n1197, B2 => 
                           n2210, ZN => n7533);
   U3249 : OAI22_X1 port map( A1 => n2208, A2 => n2238, B1 => n1199, B2 => 
                           n2210, ZN => n7534);
   U3251 : OAI22_X1 port map( A1 => n2208, A2 => n2239, B1 => n1201, B2 => 
                           n2210, ZN => n7535);
   U3253 : OAI22_X1 port map( A1 => n2208, A2 => n2240, B1 => n1203, B2 => 
                           n2210, ZN => n7536);
   U3255 : OAI22_X1 port map( A1 => n2208, A2 => n2241, B1 => n1205, B2 => 
                           n2210, ZN => n7537);
   U3260 : AND2_X1 port map( A1 => n3794, A2 => n592, ZN => n2141);
   U3261 : NOR2_X1 port map( A1 => PC_write(2), A2 => PC_write(3), ZN => n592);
   U3262 : NOR2_X1 port map( A1 => n1708, A2 => PC_write(4), ZN => n1843);
   U3263 : OAI211_X1 port map( C1 => n3528, C2 => n1144, A => Enable, B => WR, 
                           ZN => n1708);
   U3264 : INV_X1 port map( A => prevT_NT_port, ZN => n1144);
   U3266 : NAND2_X1 port map( A1 => n2242, A2 => n2243, ZN => N99);
   U3267 : NOR4_X1 port map( A1 => n2244, A2 => n2245, A3 => n2246, A4 => n2247
                           , ZN => n2243);
   U3268 : OAI221_X1 port map( B1 => n285, B2 => n2248, C1 => n251, C2 => n2249
                           , A => n2250, ZN => n2247);
   U3269 : AOI22_X1 port map( A1 => n2251, A2 => pc_target_26_28_port, B1 => 
                           n2252, B2 => pc_target_27_28_port, ZN => n2250);
   U3272 : OAI221_X1 port map( B1 => n145, B2 => n2253, C1 => n80, C2 => n2254,
                           A => n2255, ZN => n2246);
   U3273 : AOI22_X1 port map( A1 => n2256, A2 => pc_target_30_28_port, B1 => 
                           n2257, B2 => pc_target_31_28_port, ZN => n2255);
   U3276 : OAI221_X1 port map( B1 => n561, B2 => n2258, C1 => n527, C2 => n2259
                           , A => n2260, ZN => n2245);
   U3277 : AOI22_X1 port map( A1 => n2261, A2 => pc_target_18_28_port, B1 => 
                           n2262, B2 => pc_target_19_28_port, ZN => n2260);
   U3280 : OAI221_X1 port map( B1 => n355, B2 => n2263, C1 => n320, C2 => n2264
                           , A => n2265, ZN => n2244);
   U3281 : AOI22_X1 port map( A1 => n2266, A2 => pc_target_20_28_port, B1 => 
                           n2267, B2 => pc_target_21_28_port, ZN => n2265);
   U3284 : NOR4_X1 port map( A1 => n2268, A2 => n2269, A3 => n2270, A4 => n2271
                           , ZN => n2242);
   U3285 : OAI221_X1 port map( B1 => n838, B2 => n2272, C1 => n804, C2 => n2273
                           , A => n2274, ZN => n2271);
   U3286 : AOI22_X1 port map( A1 => n2275, A2 => pc_target_10_28_port, B1 => 
                           n2276, B2 => pc_target_11_28_port, ZN => n2274);
   U3289 : OAI221_X1 port map( B1 => n700, B2 => n2277, C1 => n666, C2 => n2278
                           , A => n2279, ZN => n2270);
   U3290 : AOI22_X1 port map( A1 => n2280, A2 => pc_target_14_28_port, B1 => 
                           n2281, B2 => pc_target_15_28_port, ZN => n2279);
   U3293 : OAI221_X1 port map( B1 => n1112, B2 => n2282, C1 => n1078, C2 => 
                           n2283, A => n2284, ZN => n2269);
   U3294 : AOI22_X1 port map( A1 => n2285, A2 => pc_target_2_28_port, B1 => 
                           n2286, B2 => pc_target_3_28_port, ZN => n2284);
   U3297 : OAI221_X1 port map( B1 => n975, B2 => n2287, C1 => n941, C2 => n2288
                           , A => n2289, ZN => n2268);
   U3298 : AOI22_X1 port map( A1 => n2290, A2 => pc_target_6_28_port, B1 => 
                           n2291, B2 => pc_target_7_28_port, ZN => n2289);
   U3301 : NAND2_X1 port map( A1 => n2292, A2 => n2293, ZN => N98);
   U3302 : NOR4_X1 port map( A1 => n2294, A2 => n2295, A3 => n2296, A4 => n2297
                           , ZN => n2293);
   U3303 : OAI221_X1 port map( B1 => n314, B2 => n2248, C1 => n280, C2 => n2249
                           , A => n2298, ZN => n2297);
   U3304 : AOI22_X1 port map( A1 => n2251, A2 => pc_target_26_29_port, B1 => 
                           n2252, B2 => pc_target_27_29_port, ZN => n2298);
   U3307 : OAI221_X1 port map( B1 => n174, B2 => n2253, C1 => n138, C2 => n2254
                           , A => n2299, ZN => n2296);
   U3308 : AOI22_X1 port map( A1 => n2256, A2 => pc_target_30_29_port, B1 => 
                           n2257, B2 => pc_target_31_29_port, ZN => n2299);
   U3311 : OAI221_X1 port map( B1 => n590, B2 => n2258, C1 => n556, C2 => n2259
                           , A => n2300, ZN => n2295);
   U3312 : AOI22_X1 port map( A1 => n2261, A2 => pc_target_18_29_port, B1 => 
                           n2262, B2 => pc_target_19_29_port, ZN => n2300);
   U3315 : OAI221_X1 port map( B1 => n384, B2 => n2263, C1 => n349, C2 => n2264
                           , A => n2301, ZN => n2294);
   U3316 : AOI22_X1 port map( A1 => n2266, A2 => pc_target_20_29_port, B1 => 
                           n2267, B2 => pc_target_21_29_port, ZN => n2301);
   U3319 : NOR4_X1 port map( A1 => n2302, A2 => n2303, A3 => n2304, A4 => n2305
                           , ZN => n2292);
   U3320 : OAI221_X1 port map( B1 => n867, B2 => n2272, C1 => n833, C2 => n2273
                           , A => n2306, ZN => n2305);
   U3321 : AOI22_X1 port map( A1 => n2275, A2 => pc_target_10_29_port, B1 => 
                           n2276, B2 => pc_target_11_29_port, ZN => n2306);
   U3324 : OAI221_X1 port map( B1 => n729, B2 => n2277, C1 => n695, C2 => n2278
                           , A => n2307, ZN => n2304);
   U3325 : AOI22_X1 port map( A1 => n2280, A2 => pc_target_14_29_port, B1 => 
                           n2281, B2 => pc_target_15_29_port, ZN => n2307);
   U3328 : OAI221_X1 port map( B1 => n1141, B2 => n2282, C1 => n1107, C2 => 
                           n2283, A => n2308, ZN => n2303);
   U3329 : AOI22_X1 port map( A1 => n2285, A2 => pc_target_2_29_port, B1 => 
                           n2286, B2 => pc_target_3_29_port, ZN => n2308);
   U3332 : OAI221_X1 port map( B1 => n1004, B2 => n2287, C1 => n970, C2 => 
                           n2288, A => n2309, ZN => n2302);
   U3333 : AOI22_X1 port map( A1 => n2290, A2 => pc_target_6_29_port, B1 => 
                           n2291, B2 => pc_target_7_29_port, ZN => n2309);
   U3336 : NAND2_X1 port map( A1 => n2310, A2 => n2311, ZN => N97);
   U3337 : NOR4_X1 port map( A1 => n2312, A2 => n2313, A3 => n2314, A4 => n2315
                           , ZN => n2311);
   U3338 : OAI221_X1 port map( B1 => n284, B2 => n2248, C1 => n250, C2 => n2249
                           , A => n2316, ZN => n2315);
   U3339 : AOI22_X1 port map( A1 => n2251, A2 => pc_target_26_30_port, B1 => 
                           n2252, B2 => pc_target_27_30_port, ZN => n2316);
   U3342 : OAI221_X1 port map( B1 => n144, B2 => n2253, C1 => n78, C2 => n2254,
                           A => n2317, ZN => n2314);
   U3343 : AOI22_X1 port map( A1 => n2256, A2 => pc_target_30_30_port, B1 => 
                           n2257, B2 => pc_target_31_30_port, ZN => n2317);
   U3346 : OAI221_X1 port map( B1 => n560, B2 => n2258, C1 => n526, C2 => n2259
                           , A => n2318, ZN => n2313);
   U3347 : AOI22_X1 port map( A1 => n2261, A2 => pc_target_18_30_port, B1 => 
                           n2262, B2 => pc_target_19_30_port, ZN => n2318);
   U3350 : OAI221_X1 port map( B1 => n354, B2 => n2263, C1 => n319, C2 => n2264
                           , A => n2319, ZN => n2312);
   U3351 : AOI22_X1 port map( A1 => n2266, A2 => pc_target_20_30_port, B1 => 
                           n2267, B2 => pc_target_21_30_port, ZN => n2319);
   U3354 : NOR4_X1 port map( A1 => n2320, A2 => n2321, A3 => n2322, A4 => n2323
                           , ZN => n2310);
   U3355 : OAI221_X1 port map( B1 => n837, B2 => n2272, C1 => n803, C2 => n2273
                           , A => n2324, ZN => n2323);
   U3356 : AOI22_X1 port map( A1 => n2275, A2 => pc_target_10_30_port, B1 => 
                           n2276, B2 => pc_target_11_30_port, ZN => n2324);
   U3359 : OAI221_X1 port map( B1 => n699, B2 => n2277, C1 => n665, C2 => n2278
                           , A => n2325, ZN => n2322);
   U3360 : AOI22_X1 port map( A1 => n2280, A2 => pc_target_14_30_port, B1 => 
                           n2281, B2 => pc_target_15_30_port, ZN => n2325);
   U3363 : OAI221_X1 port map( B1 => n1111, B2 => n2282, C1 => n1077, C2 => 
                           n2283, A => n2326, ZN => n2321);
   U3364 : AOI22_X1 port map( A1 => n2285, A2 => pc_target_2_30_port, B1 => 
                           n2286, B2 => pc_target_3_30_port, ZN => n2326);
   U3367 : OAI221_X1 port map( B1 => n974, B2 => n2287, C1 => n940, C2 => n2288
                           , A => n2327, ZN => n2320);
   U3368 : AOI22_X1 port map( A1 => n2290, A2 => pc_target_6_30_port, B1 => 
                           n2291, B2 => pc_target_7_30_port, ZN => n2327);
   U3371 : NAND2_X1 port map( A1 => n2328, A2 => n2329, ZN => N96);
   U3372 : NOR4_X1 port map( A1 => n2330, A2 => n2331, A3 => n2332, A4 => n2333
                           , ZN => n2329);
   U3373 : OAI221_X1 port map( B1 => n315, B2 => n2248, C1 => n281, C2 => n2249
                           , A => n2334, ZN => n2333);
   U3374 : AOI22_X1 port map( A1 => n2251, A2 => pc_target_26_31_port, B1 => 
                           n2252, B2 => pc_target_27_31_port, ZN => n2334);
   U3377 : OAI221_X1 port map( B1 => n175, B2 => n2253, C1 => n140, C2 => n2254
                           , A => n2335, ZN => n2332);
   U3378 : AOI22_X1 port map( A1 => n2256, A2 => pc_target_30_31_port, B1 => 
                           n2257, B2 => pc_target_31_31_port, ZN => n2335);
   U3381 : OAI221_X1 port map( B1 => n591, B2 => n2258, C1 => n557, C2 => n2259
                           , A => n2336, ZN => n2331);
   U3382 : AOI22_X1 port map( A1 => n2261, A2 => pc_target_18_31_port, B1 => 
                           n2262, B2 => pc_target_19_31_port, ZN => n2336);
   U3385 : OAI221_X1 port map( B1 => n385, B2 => n2263, C1 => n350, C2 => n2264
                           , A => n2337, ZN => n2330);
   U3386 : AOI22_X1 port map( A1 => n2266, A2 => pc_target_20_31_port, B1 => 
                           n2267, B2 => pc_target_21_31_port, ZN => n2337);
   U3389 : NOR4_X1 port map( A1 => n2338, A2 => n2339, A3 => n2340, A4 => n2341
                           , ZN => n2328);
   U3390 : OAI221_X1 port map( B1 => n868, B2 => n2272, C1 => n834, C2 => n2273
                           , A => n2342, ZN => n2341);
   U3391 : AOI22_X1 port map( A1 => n2275, A2 => pc_target_10_31_port, B1 => 
                           n2276, B2 => pc_target_11_31_port, ZN => n2342);
   U3394 : OAI221_X1 port map( B1 => n730, B2 => n2277, C1 => n696, C2 => n2278
                           , A => n2343, ZN => n2340);
   U3395 : AOI22_X1 port map( A1 => n2280, A2 => pc_target_14_31_port, B1 => 
                           n2281, B2 => pc_target_15_31_port, ZN => n2343);
   U3398 : OAI221_X1 port map( B1 => n1142, B2 => n2282, C1 => n1108, C2 => 
                           n2283, A => n2344, ZN => n2339);
   U3399 : AOI22_X1 port map( A1 => n2285, A2 => pc_target_2_31_port, B1 => 
                           n2286, B2 => pc_target_3_31_port, ZN => n2344);
   U3402 : OAI221_X1 port map( B1 => n1005, B2 => n2287, C1 => n971, C2 => 
                           n2288, A => n2345, ZN => n2338);
   U3403 : AOI22_X1 port map( A1 => n2290, A2 => pc_target_6_31_port, B1 => 
                           n2291, B2 => pc_target_7_31_port, ZN => n2345);
   U3406 : NAND2_X1 port map( A1 => n2346, A2 => n2347, ZN => N219);
   U3407 : NOR4_X1 port map( A1 => n2348, A2 => n2349, A3 => n2350, A4 => n2351
                           , ZN => n2347);
   U3424 : NOR4_X1 port map( A1 => n2356, A2 => n2357, A3 => n2358, A4 => n2359
                           , ZN => n2346);
   U3441 : NAND2_X1 port map( A1 => n2364, A2 => n2365, ZN => N218);
   U3442 : NOR4_X1 port map( A1 => n2366, A2 => n2367, A3 => n2368, A4 => n2369
                           , ZN => n2365);
   U3444 : AOI22_X1 port map( A1 => n2251, A2 => pc_lut_26_1_port, B1 => n2252,
                           B2 => pc_lut_27_1_port, ZN => n2370);
   U3448 : AOI22_X1 port map( A1 => n2256, A2 => pc_lut_30_1_port, B1 => n2257,
                           B2 => pc_lut_31_1_port, ZN => n2371);
   U3452 : AOI22_X1 port map( A1 => n2261, A2 => pc_lut_18_1_port, B1 => n2262,
                           B2 => pc_lut_19_1_port, ZN => n2372);
   U3459 : NOR4_X1 port map( A1 => n2374, A2 => n2375, A3 => n2376, A4 => n2377
                           , ZN => n2364);
   U3461 : AOI22_X1 port map( A1 => n2275, A2 => pc_lut_10_1_port, B1 => n2276,
                           B2 => pc_lut_11_1_port, ZN => n2378);
   U3465 : AOI22_X1 port map( A1 => n2280, A2 => pc_lut_14_1_port, B1 => n2281,
                           B2 => pc_lut_15_1_port, ZN => n2379);
   U3469 : AOI22_X1 port map( A1 => n2285, A2 => pc_lut_2_1_port, B1 => n2286, 
                           B2 => pc_lut_3_1_port, ZN => n2380);
   U3473 : AOI22_X1 port map( A1 => n2290, A2 => pc_lut_6_1_port, B1 => n2291, 
                           B2 => pc_lut_7_1_port, ZN => n2381);
   U3476 : NAND2_X1 port map( A1 => n2382, A2 => n2383, ZN => N217);
   U3482 : OAI221_X1 port map( B1 => n1291, B2 => n2253, C1 => n1257, C2 => 
                           n2254, A => n2389, ZN => n2386);
   U3483 : AOI22_X1 port map( A1 => n2256, A2 => pc_lut_30_2_port, B1 => n2257,
                           B2 => pc_lut_31_2_port, ZN => n2389);
   U3490 : OAI221_X1 port map( B1 => n1495, B2 => n2263, C1 => n1460, C2 => 
                           n2264, A => n2391, ZN => n2384);
   U3491 : AOI22_X1 port map( A1 => n2266, A2 => pc_lut_20_2_port, B1 => n2267,
                           B2 => pc_lut_21_2_port, ZN => n2391);
   U3499 : OAI221_X1 port map( B1 => n1825, B2 => n2277, C1 => n1791, C2 => 
                           n2278, A => n2397, ZN => n2394);
   U3500 : AOI22_X1 port map( A1 => n2280, A2 => pc_lut_14_2_port, B1 => n2281,
                           B2 => pc_lut_15_2_port, ZN => n2397);
   U3507 : OAI221_X1 port map( B1 => n2092, B2 => n2287, C1 => n2058, C2 => 
                           n2288, A => n2399, ZN => n2392);
   U3508 : AOI22_X1 port map( A1 => n2290, A2 => pc_lut_6_2_port, B1 => n2291, 
                           B2 => pc_lut_7_2_port, ZN => n2399);
   U3511 : NAND2_X1 port map( A1 => n2400, A2 => n2401, ZN => N216);
   U3513 : OAI221_X1 port map( B1 => n1429, B2 => n2248, C1 => n1395, C2 => 
                           n2249, A => n2406, ZN => n2405);
   U3514 : AOI22_X1 port map( A1 => n2251, A2 => pc_lut_26_3_port, B1 => n2252,
                           B2 => pc_lut_27_3_port, ZN => n2406);
   U3517 : OAI221_X1 port map( B1 => n1294, B2 => n2253, C1 => n1260, C2 => 
                           n2254, A => n2407, ZN => n2404);
   U3518 : AOI22_X1 port map( A1 => n2256, A2 => pc_lut_30_3_port, B1 => n2257,
                           B2 => pc_lut_31_3_port, ZN => n2407);
   U3530 : OAI221_X1 port map( B1 => n1963, B2 => n2272, C1 => n1929, C2 => 
                           n2273, A => n2414, ZN => n2413);
   U3531 : AOI22_X1 port map( A1 => n2275, A2 => pc_lut_10_3_port, B1 => n2276,
                           B2 => pc_lut_11_3_port, ZN => n2414);
   U3534 : OAI221_X1 port map( B1 => n1828, B2 => n2277, C1 => n1794, C2 => 
                           n2278, A => n2415, ZN => n2412);
   U3535 : AOI22_X1 port map( A1 => n2280, A2 => pc_lut_14_3_port, B1 => n2281,
                           B2 => pc_lut_15_3_port, ZN => n2415);
   U3547 : NOR4_X1 port map( A1 => n2420, A2 => n2421, A3 => n2422, A4 => n2423
                           , ZN => n2419);
   U3548 : OAI221_X1 port map( B1 => n1425, B2 => n2248, C1 => n1391, C2 => 
                           n2249, A => n2424, ZN => n2423);
   U3549 : AOI22_X1 port map( A1 => n2251, A2 => pc_lut_26_4_port, B1 => n2252,
                           B2 => pc_lut_27_4_port, ZN => n2424);
   U3552 : OAI221_X1 port map( B1 => n1290, B2 => n2253, C1 => n1255, C2 => 
                           n2254, A => n2425, ZN => n2422);
   U3553 : AOI22_X1 port map( A1 => n2256, A2 => pc_lut_30_4_port, B1 => n2257,
                           B2 => pc_lut_31_4_port, ZN => n2425);
   U3556 : OAI221_X1 port map( B1 => n1689, B2 => n2258, C1 => n1655, C2 => 
                           n2259, A => n2426, ZN => n2421);
   U3557 : AOI22_X1 port map( A1 => n2261, A2 => pc_lut_18_4_port, B1 => n2262,
                           B2 => pc_lut_19_4_port, ZN => n2426);
   U3560 : OAI221_X1 port map( B1 => n1494, B2 => n2263, C1 => n1459, C2 => 
                           n2264, A => n2427, ZN => n2420);
   U3561 : AOI22_X1 port map( A1 => n2266, A2 => pc_lut_20_4_port, B1 => n2267,
                           B2 => pc_lut_21_4_port, ZN => n2427);
   U3581 : NAND2_X1 port map( A1 => n2436, A2 => n2437, ZN => N214);
   U3582 : NOR4_X1 port map( A1 => n2438, A2 => n2439, A3 => n2440, A4 => n2441
                           , ZN => n2437);
   U3583 : OAI221_X1 port map( B1 => n1430, B2 => n2248, C1 => n1396, C2 => 
                           n2249, A => n2442, ZN => n2441);
   U3584 : AOI22_X1 port map( A1 => n2251, A2 => pc_lut_26_5_port, B1 => n2252,
                           B2 => pc_lut_27_5_port, ZN => n2442);
   U3587 : OAI221_X1 port map( B1 => n1295, B2 => n2253, C1 => n1261, C2 => 
                           n2254, A => n2443, ZN => n2440);
   U3588 : AOI22_X1 port map( A1 => n2256, A2 => pc_lut_30_5_port, B1 => n2257,
                           B2 => pc_lut_31_5_port, ZN => n2443);
   U3591 : OAI221_X1 port map( B1 => n1694, B2 => n2258, C1 => n1660, C2 => 
                           n2259, A => n2444, ZN => n2439);
   U3592 : AOI22_X1 port map( A1 => n2261, A2 => pc_lut_18_5_port, B1 => n2262,
                           B2 => pc_lut_19_5_port, ZN => n2444);
   U3595 : OAI221_X1 port map( B1 => n1499, B2 => n2263, C1 => n1464, C2 => 
                           n2264, A => n2445, ZN => n2438);
   U3596 : AOI22_X1 port map( A1 => n2266, A2 => pc_lut_20_5_port, B1 => n2267,
                           B2 => pc_lut_21_5_port, ZN => n2445);
   U3599 : NOR4_X1 port map( A1 => n2446, A2 => n2447, A3 => n2448, A4 => n2449
                           , ZN => n2436);
   U3600 : OAI221_X1 port map( B1 => n1964, B2 => n2272, C1 => n1930, C2 => 
                           n2273, A => n2450, ZN => n2449);
   U3601 : AOI22_X1 port map( A1 => n2275, A2 => pc_lut_10_5_port, B1 => n2276,
                           B2 => pc_lut_11_5_port, ZN => n2450);
   U3604 : OAI221_X1 port map( B1 => n1829, B2 => n2277, C1 => n1795, C2 => 
                           n2278, A => n2451, ZN => n2448);
   U3605 : AOI22_X1 port map( A1 => n2280, A2 => pc_lut_14_5_port, B1 => n2281,
                           B2 => pc_lut_15_5_port, ZN => n2451);
   U3608 : OAI221_X1 port map( B1 => n2228, B2 => n2282, C1 => n2194, C2 => 
                           n2283, A => n2452, ZN => n2447);
   U3609 : AOI22_X1 port map( A1 => n2285, A2 => pc_lut_2_5_port, B1 => n2286, 
                           B2 => pc_lut_3_5_port, ZN => n2452);
   U3612 : OAI221_X1 port map( B1 => n2096, B2 => n2287, C1 => n2062, C2 => 
                           n2288, A => n2453, ZN => n2446);
   U3613 : AOI22_X1 port map( A1 => n2290, A2 => pc_lut_6_5_port, B1 => n2291, 
                           B2 => pc_lut_7_5_port, ZN => n2453);
   U3616 : NAND2_X1 port map( A1 => n2454, A2 => n2455, ZN => N213);
   U3617 : NOR4_X1 port map( A1 => n2456, A2 => n2457, A3 => n2458, A4 => n2459
                           , ZN => n2455);
   U3618 : OAI221_X1 port map( B1 => n1424, B2 => n2248, C1 => n1390, C2 => 
                           n2249, A => n2460, ZN => n2459);
   U3619 : AOI22_X1 port map( A1 => n2251, A2 => pc_lut_26_6_port, B1 => n2252,
                           B2 => pc_lut_27_6_port, ZN => n2460);
   U3622 : OAI221_X1 port map( B1 => n1289, B2 => n2253, C1 => n1254, C2 => 
                           n2254, A => n2461, ZN => n2458);
   U3623 : AOI22_X1 port map( A1 => n2256, A2 => pc_lut_30_6_port, B1 => n2257,
                           B2 => pc_lut_31_6_port, ZN => n2461);
   U3626 : OAI221_X1 port map( B1 => n1688, B2 => n2258, C1 => n1654, C2 => 
                           n2259, A => n2462, ZN => n2457);
   U3627 : AOI22_X1 port map( A1 => n2261, A2 => pc_lut_18_6_port, B1 => n2262,
                           B2 => pc_lut_19_6_port, ZN => n2462);
   U3630 : OAI221_X1 port map( B1 => n1493, B2 => n2263, C1 => n1458, C2 => 
                           n2264, A => n2463, ZN => n2456);
   U3631 : AOI22_X1 port map( A1 => n2266, A2 => pc_lut_20_6_port, B1 => n2267,
                           B2 => pc_lut_21_6_port, ZN => n2463);
   U3634 : NOR4_X1 port map( A1 => n2464, A2 => n2465, A3 => n2466, A4 => n2467
                           , ZN => n2454);
   U3635 : OAI221_X1 port map( B1 => n1958, B2 => n2272, C1 => n1924, C2 => 
                           n2273, A => n2468, ZN => n2467);
   U3636 : AOI22_X1 port map( A1 => n2275, A2 => pc_lut_10_6_port, B1 => n2276,
                           B2 => pc_lut_11_6_port, ZN => n2468);
   U3639 : OAI221_X1 port map( B1 => n1823, B2 => n2277, C1 => n1789, C2 => 
                           n2278, A => n2469, ZN => n2466);
   U3640 : AOI22_X1 port map( A1 => n2280, A2 => pc_lut_14_6_port, B1 => n2281,
                           B2 => pc_lut_15_6_port, ZN => n2469);
   U3643 : OAI221_X1 port map( B1 => n2222, B2 => n2282, C1 => n2188, C2 => 
                           n2283, A => n2470, ZN => n2465);
   U3644 : AOI22_X1 port map( A1 => n2285, A2 => pc_lut_2_6_port, B1 => n2286, 
                           B2 => pc_lut_3_6_port, ZN => n2470);
   U3647 : OAI221_X1 port map( B1 => n2090, B2 => n2287, C1 => n2056, C2 => 
                           n2288, A => n2471, ZN => n2464);
   U3648 : AOI22_X1 port map( A1 => n2290, A2 => pc_lut_6_6_port, B1 => n2291, 
                           B2 => pc_lut_7_6_port, ZN => n2471);
   U3651 : NAND2_X1 port map( A1 => n2472, A2 => n2473, ZN => N212);
   U3652 : NOR4_X1 port map( A1 => n2474, A2 => n2475, A3 => n2476, A4 => n2477
                           , ZN => n2473);
   U3653 : OAI221_X1 port map( B1 => n1431, B2 => n2248, C1 => n1397, C2 => 
                           n2249, A => n2478, ZN => n2477);
   U3654 : AOI22_X1 port map( A1 => n2251, A2 => pc_lut_26_7_port, B1 => n2252,
                           B2 => pc_lut_27_7_port, ZN => n2478);
   U3657 : OAI221_X1 port map( B1 => n1296, B2 => n2253, C1 => n1262, C2 => 
                           n2254, A => n2479, ZN => n2476);
   U3658 : AOI22_X1 port map( A1 => n2256, A2 => pc_lut_30_7_port, B1 => n2257,
                           B2 => pc_lut_31_7_port, ZN => n2479);
   U3661 : OAI221_X1 port map( B1 => n1695, B2 => n2258, C1 => n1661, C2 => 
                           n2259, A => n2480, ZN => n2475);
   U3662 : AOI22_X1 port map( A1 => n2261, A2 => pc_lut_18_7_port, B1 => n2262,
                           B2 => pc_lut_19_7_port, ZN => n2480);
   U3665 : OAI221_X1 port map( B1 => n1500, B2 => n2263, C1 => n1465, C2 => 
                           n2264, A => n2481, ZN => n2474);
   U3666 : AOI22_X1 port map( A1 => n2266, A2 => pc_lut_20_7_port, B1 => n2267,
                           B2 => pc_lut_21_7_port, ZN => n2481);
   U3669 : NOR4_X1 port map( A1 => n2482, A2 => n2483, A3 => n2484, A4 => n2485
                           , ZN => n2472);
   U3670 : OAI221_X1 port map( B1 => n1965, B2 => n2272, C1 => n1931, C2 => 
                           n2273, A => n2486, ZN => n2485);
   U3671 : AOI22_X1 port map( A1 => n2275, A2 => pc_lut_10_7_port, B1 => n2276,
                           B2 => pc_lut_11_7_port, ZN => n2486);
   U3674 : OAI221_X1 port map( B1 => n1830, B2 => n2277, C1 => n1796, C2 => 
                           n2278, A => n2487, ZN => n2484);
   U3675 : AOI22_X1 port map( A1 => n2280, A2 => pc_lut_14_7_port, B1 => n2281,
                           B2 => pc_lut_15_7_port, ZN => n2487);
   U3678 : OAI221_X1 port map( B1 => n2229, B2 => n2282, C1 => n2195, C2 => 
                           n2283, A => n2488, ZN => n2483);
   U3679 : AOI22_X1 port map( A1 => n2285, A2 => pc_lut_2_7_port, B1 => n2286, 
                           B2 => pc_lut_3_7_port, ZN => n2488);
   U3682 : OAI221_X1 port map( B1 => n2097, B2 => n2287, C1 => n2063, C2 => 
                           n2288, A => n2489, ZN => n2482);
   U3683 : AOI22_X1 port map( A1 => n2290, A2 => pc_lut_6_7_port, B1 => n2291, 
                           B2 => pc_lut_7_7_port, ZN => n2489);
   U3686 : NAND2_X1 port map( A1 => n2490, A2 => n2491, ZN => N211);
   U3687 : NOR4_X1 port map( A1 => n2492, A2 => n2493, A3 => n2494, A4 => n2495
                           , ZN => n2491);
   U3688 : OAI221_X1 port map( B1 => n1423, B2 => n2248, C1 => n1389, C2 => 
                           n2249, A => n2496, ZN => n2495);
   U3689 : AOI22_X1 port map( A1 => n2251, A2 => pc_lut_26_8_port, B1 => n2252,
                           B2 => pc_lut_27_8_port, ZN => n2496);
   U3692 : OAI221_X1 port map( B1 => n1288, B2 => n2253, C1 => n1253, C2 => 
                           n2254, A => n2497, ZN => n2494);
   U3693 : AOI22_X1 port map( A1 => n2256, A2 => pc_lut_30_8_port, B1 => n2257,
                           B2 => pc_lut_31_8_port, ZN => n2497);
   U3696 : OAI221_X1 port map( B1 => n1687, B2 => n2258, C1 => n1653, C2 => 
                           n2259, A => n2498, ZN => n2493);
   U3697 : AOI22_X1 port map( A1 => n2261, A2 => pc_lut_18_8_port, B1 => n2262,
                           B2 => pc_lut_19_8_port, ZN => n2498);
   U3700 : OAI221_X1 port map( B1 => n1492, B2 => n2263, C1 => n1457, C2 => 
                           n2264, A => n2499, ZN => n2492);
   U3701 : AOI22_X1 port map( A1 => n2266, A2 => pc_lut_20_8_port, B1 => n2267,
                           B2 => pc_lut_21_8_port, ZN => n2499);
   U3704 : NOR4_X1 port map( A1 => n2500, A2 => n2501, A3 => n2502, A4 => n2503
                           , ZN => n2490);
   U3705 : OAI221_X1 port map( B1 => n1957, B2 => n2272, C1 => n1923, C2 => 
                           n2273, A => n2504, ZN => n2503);
   U3706 : AOI22_X1 port map( A1 => n2275, A2 => pc_lut_10_8_port, B1 => n2276,
                           B2 => pc_lut_11_8_port, ZN => n2504);
   U3709 : OAI221_X1 port map( B1 => n1822, B2 => n2277, C1 => n1788, C2 => 
                           n2278, A => n2505, ZN => n2502);
   U3710 : AOI22_X1 port map( A1 => n2280, A2 => pc_lut_14_8_port, B1 => n2281,
                           B2 => pc_lut_15_8_port, ZN => n2505);
   U3713 : OAI221_X1 port map( B1 => n2221, B2 => n2282, C1 => n2187, C2 => 
                           n2283, A => n2506, ZN => n2501);
   U3714 : AOI22_X1 port map( A1 => n2285, A2 => pc_lut_2_8_port, B1 => n2286, 
                           B2 => pc_lut_3_8_port, ZN => n2506);
   U3717 : OAI221_X1 port map( B1 => n2089, B2 => n2287, C1 => n2055, C2 => 
                           n2288, A => n2507, ZN => n2500);
   U3718 : AOI22_X1 port map( A1 => n2290, A2 => pc_lut_6_8_port, B1 => n2291, 
                           B2 => pc_lut_7_8_port, ZN => n2507);
   U3721 : NAND2_X1 port map( A1 => n2508, A2 => n2509, ZN => N210);
   U3722 : NOR4_X1 port map( A1 => n2510, A2 => n2511, A3 => n2512, A4 => n2513
                           , ZN => n2509);
   U3723 : OAI221_X1 port map( B1 => n1432, B2 => n2248, C1 => n1398, C2 => 
                           n2249, A => n2514, ZN => n2513);
   U3724 : AOI22_X1 port map( A1 => n2251, A2 => pc_lut_26_9_port, B1 => n2252,
                           B2 => pc_lut_27_9_port, ZN => n2514);
   U3727 : OAI221_X1 port map( B1 => n1297, B2 => n2253, C1 => n1263, C2 => 
                           n2254, A => n2515, ZN => n2512);
   U3728 : AOI22_X1 port map( A1 => n2256, A2 => pc_lut_30_9_port, B1 => n2257,
                           B2 => pc_lut_31_9_port, ZN => n2515);
   U3731 : OAI221_X1 port map( B1 => n1696, B2 => n2258, C1 => n1662, C2 => 
                           n2259, A => n2516, ZN => n2511);
   U3732 : AOI22_X1 port map( A1 => n2261, A2 => pc_lut_18_9_port, B1 => n2262,
                           B2 => pc_lut_19_9_port, ZN => n2516);
   U3735 : OAI221_X1 port map( B1 => n1501, B2 => n2263, C1 => n1466, C2 => 
                           n2264, A => n2517, ZN => n2510);
   U3736 : AOI22_X1 port map( A1 => n2266, A2 => pc_lut_20_9_port, B1 => n2267,
                           B2 => pc_lut_21_9_port, ZN => n2517);
   U3739 : NOR4_X1 port map( A1 => n2518, A2 => n2519, A3 => n2520, A4 => n2521
                           , ZN => n2508);
   U3740 : OAI221_X1 port map( B1 => n1966, B2 => n2272, C1 => n1932, C2 => 
                           n2273, A => n2522, ZN => n2521);
   U3741 : AOI22_X1 port map( A1 => n2275, A2 => pc_lut_10_9_port, B1 => n2276,
                           B2 => pc_lut_11_9_port, ZN => n2522);
   U3744 : OAI221_X1 port map( B1 => n1831, B2 => n2277, C1 => n1797, C2 => 
                           n2278, A => n2523, ZN => n2520);
   U3745 : AOI22_X1 port map( A1 => n2280, A2 => pc_lut_14_9_port, B1 => n2281,
                           B2 => pc_lut_15_9_port, ZN => n2523);
   U3748 : OAI221_X1 port map( B1 => n2230, B2 => n2282, C1 => n2196, C2 => 
                           n2283, A => n2524, ZN => n2519);
   U3749 : AOI22_X1 port map( A1 => n2285, A2 => pc_lut_2_9_port, B1 => n2286, 
                           B2 => pc_lut_3_9_port, ZN => n2524);
   U3752 : OAI221_X1 port map( B1 => n2098, B2 => n2287, C1 => n2064, C2 => 
                           n2288, A => n2525, ZN => n2518);
   U3753 : AOI22_X1 port map( A1 => n2290, A2 => pc_lut_6_9_port, B1 => n2291, 
                           B2 => pc_lut_7_9_port, ZN => n2525);
   U3756 : NAND2_X1 port map( A1 => n2526, A2 => n2527, ZN => N209);
   U3757 : NOR4_X1 port map( A1 => n2528, A2 => n2529, A3 => n2530, A4 => n2531
                           , ZN => n2527);
   U3758 : OAI221_X1 port map( B1 => n1422, B2 => n2248, C1 => n1388, C2 => 
                           n2249, A => n2532, ZN => n2531);
   U3759 : AOI22_X1 port map( A1 => n2251, A2 => pc_lut_26_10_port, B1 => n2252
                           , B2 => pc_lut_27_10_port, ZN => n2532);
   U3762 : OAI221_X1 port map( B1 => n1287, B2 => n2253, C1 => n1252, C2 => 
                           n2254, A => n2533, ZN => n2530);
   U3763 : AOI22_X1 port map( A1 => n2256, A2 => pc_lut_30_10_port, B1 => n2257
                           , B2 => pc_lut_31_10_port, ZN => n2533);
   U3766 : OAI221_X1 port map( B1 => n1686, B2 => n2258, C1 => n1652, C2 => 
                           n2259, A => n2534, ZN => n2529);
   U3767 : AOI22_X1 port map( A1 => n2261, A2 => pc_lut_18_10_port, B1 => n2262
                           , B2 => pc_lut_19_10_port, ZN => n2534);
   U3770 : OAI221_X1 port map( B1 => n1491, B2 => n2263, C1 => n1456, C2 => 
                           n2264, A => n2535, ZN => n2528);
   U3771 : AOI22_X1 port map( A1 => n2266, A2 => pc_lut_20_10_port, B1 => n2267
                           , B2 => pc_lut_21_10_port, ZN => n2535);
   U3774 : NOR4_X1 port map( A1 => n2536, A2 => n2537, A3 => n2538, A4 => n2539
                           , ZN => n2526);
   U3775 : OAI221_X1 port map( B1 => n1956, B2 => n2272, C1 => n1922, C2 => 
                           n2273, A => n2540, ZN => n2539);
   U3776 : AOI22_X1 port map( A1 => n2275, A2 => pc_lut_10_10_port, B1 => n2276
                           , B2 => pc_lut_11_10_port, ZN => n2540);
   U3779 : OAI221_X1 port map( B1 => n1821, B2 => n2277, C1 => n1787, C2 => 
                           n2278, A => n2541, ZN => n2538);
   U3780 : AOI22_X1 port map( A1 => n2280, A2 => pc_lut_14_10_port, B1 => n2281
                           , B2 => pc_lut_15_10_port, ZN => n2541);
   U3783 : OAI221_X1 port map( B1 => n2220, B2 => n2282, C1 => n2186, C2 => 
                           n2283, A => n2542, ZN => n2537);
   U3784 : AOI22_X1 port map( A1 => n2285, A2 => pc_lut_2_10_port, B1 => n2286,
                           B2 => pc_lut_3_10_port, ZN => n2542);
   U3787 : OAI221_X1 port map( B1 => n2088, B2 => n2287, C1 => n2054, C2 => 
                           n2288, A => n2543, ZN => n2536);
   U3788 : AOI22_X1 port map( A1 => n2290, A2 => pc_lut_6_10_port, B1 => n2291,
                           B2 => pc_lut_7_10_port, ZN => n2543);
   U3791 : NAND2_X1 port map( A1 => n2544, A2 => n2545, ZN => N208);
   U3792 : NOR4_X1 port map( A1 => n2546, A2 => n2547, A3 => n2548, A4 => n2549
                           , ZN => n2545);
   U3793 : OAI221_X1 port map( B1 => n1433, B2 => n2248, C1 => n1399, C2 => 
                           n2249, A => n2550, ZN => n2549);
   U3794 : AOI22_X1 port map( A1 => n2251, A2 => pc_lut_26_11_port, B1 => n2252
                           , B2 => pc_lut_27_11_port, ZN => n2550);
   U3797 : OAI221_X1 port map( B1 => n1298, B2 => n2253, C1 => n1264, C2 => 
                           n2254, A => n2551, ZN => n2548);
   U3798 : AOI22_X1 port map( A1 => n2256, A2 => pc_lut_30_11_port, B1 => n2257
                           , B2 => pc_lut_31_11_port, ZN => n2551);
   U3801 : OAI221_X1 port map( B1 => n1697, B2 => n2258, C1 => n1663, C2 => 
                           n2259, A => n2552, ZN => n2547);
   U3802 : AOI22_X1 port map( A1 => n2261, A2 => pc_lut_18_11_port, B1 => n2262
                           , B2 => pc_lut_19_11_port, ZN => n2552);
   U3805 : OAI221_X1 port map( B1 => n1502, B2 => n2263, C1 => n1467, C2 => 
                           n2264, A => n2553, ZN => n2546);
   U3806 : AOI22_X1 port map( A1 => n2266, A2 => pc_lut_20_11_port, B1 => n2267
                           , B2 => pc_lut_21_11_port, ZN => n2553);
   U3809 : NOR4_X1 port map( A1 => n2554, A2 => n2555, A3 => n2556, A4 => n2557
                           , ZN => n2544);
   U3810 : OAI221_X1 port map( B1 => n1967, B2 => n2272, C1 => n1933, C2 => 
                           n2273, A => n2558, ZN => n2557);
   U3811 : AOI22_X1 port map( A1 => n2275, A2 => pc_lut_10_11_port, B1 => n2276
                           , B2 => pc_lut_11_11_port, ZN => n2558);
   U3814 : OAI221_X1 port map( B1 => n1832, B2 => n2277, C1 => n1798, C2 => 
                           n2278, A => n2559, ZN => n2556);
   U3815 : AOI22_X1 port map( A1 => n2280, A2 => pc_lut_14_11_port, B1 => n2281
                           , B2 => pc_lut_15_11_port, ZN => n2559);
   U3818 : OAI221_X1 port map( B1 => n2231, B2 => n2282, C1 => n2197, C2 => 
                           n2283, A => n2560, ZN => n2555);
   U3819 : AOI22_X1 port map( A1 => n2285, A2 => pc_lut_2_11_port, B1 => n2286,
                           B2 => pc_lut_3_11_port, ZN => n2560);
   U3822 : OAI221_X1 port map( B1 => n2099, B2 => n2287, C1 => n2065, C2 => 
                           n2288, A => n2561, ZN => n2554);
   U3823 : AOI22_X1 port map( A1 => n2290, A2 => pc_lut_6_11_port, B1 => n2291,
                           B2 => pc_lut_7_11_port, ZN => n2561);
   U3826 : NAND2_X1 port map( A1 => n2562, A2 => n2563, ZN => N207);
   U3827 : NOR4_X1 port map( A1 => n2564, A2 => n2565, A3 => n2566, A4 => n2567
                           , ZN => n2563);
   U3828 : OAI221_X1 port map( B1 => n1421, B2 => n2248, C1 => n1387, C2 => 
                           n2249, A => n2568, ZN => n2567);
   U3829 : AOI22_X1 port map( A1 => n2251, A2 => pc_lut_26_12_port, B1 => n2252
                           , B2 => pc_lut_27_12_port, ZN => n2568);
   U3832 : OAI221_X1 port map( B1 => n1286, B2 => n2253, C1 => n1251, C2 => 
                           n2254, A => n2569, ZN => n2566);
   U3833 : AOI22_X1 port map( A1 => n2256, A2 => pc_lut_30_12_port, B1 => n2257
                           , B2 => pc_lut_31_12_port, ZN => n2569);
   U3836 : OAI221_X1 port map( B1 => n1685, B2 => n2258, C1 => n1651, C2 => 
                           n2259, A => n2570, ZN => n2565);
   U3837 : AOI22_X1 port map( A1 => n2261, A2 => pc_lut_18_12_port, B1 => n2262
                           , B2 => pc_lut_19_12_port, ZN => n2570);
   U3840 : OAI221_X1 port map( B1 => n1490, B2 => n2263, C1 => n1455, C2 => 
                           n2264, A => n2571, ZN => n2564);
   U3841 : AOI22_X1 port map( A1 => n2266, A2 => pc_lut_20_12_port, B1 => n2267
                           , B2 => pc_lut_21_12_port, ZN => n2571);
   U3844 : NOR4_X1 port map( A1 => n2572, A2 => n2573, A3 => n2574, A4 => n2575
                           , ZN => n2562);
   U3845 : OAI221_X1 port map( B1 => n1955, B2 => n2272, C1 => n1921, C2 => 
                           n2273, A => n2576, ZN => n2575);
   U3846 : AOI22_X1 port map( A1 => n2275, A2 => pc_lut_10_12_port, B1 => n2276
                           , B2 => pc_lut_11_12_port, ZN => n2576);
   U3849 : OAI221_X1 port map( B1 => n1820, B2 => n2277, C1 => n1786, C2 => 
                           n2278, A => n2577, ZN => n2574);
   U3850 : AOI22_X1 port map( A1 => n2280, A2 => pc_lut_14_12_port, B1 => n2281
                           , B2 => pc_lut_15_12_port, ZN => n2577);
   U3853 : OAI221_X1 port map( B1 => n2219, B2 => n2282, C1 => n2185, C2 => 
                           n2283, A => n2578, ZN => n2573);
   U3854 : AOI22_X1 port map( A1 => n2285, A2 => pc_lut_2_12_port, B1 => n2286,
                           B2 => pc_lut_3_12_port, ZN => n2578);
   U3857 : OAI221_X1 port map( B1 => n2087, B2 => n2287, C1 => n2053, C2 => 
                           n2288, A => n2579, ZN => n2572);
   U3858 : AOI22_X1 port map( A1 => n2290, A2 => pc_lut_6_12_port, B1 => n2291,
                           B2 => pc_lut_7_12_port, ZN => n2579);
   U3861 : NAND2_X1 port map( A1 => n2580, A2 => n2581, ZN => N206);
   U3862 : NOR4_X1 port map( A1 => n2582, A2 => n2583, A3 => n2584, A4 => n2585
                           , ZN => n2581);
   U3863 : OAI221_X1 port map( B1 => n1434, B2 => n2248, C1 => n1400, C2 => 
                           n2249, A => n2586, ZN => n2585);
   U3864 : AOI22_X1 port map( A1 => n2251, A2 => pc_lut_26_13_port, B1 => n2252
                           , B2 => pc_lut_27_13_port, ZN => n2586);
   U3867 : OAI221_X1 port map( B1 => n1299, B2 => n2253, C1 => n1265, C2 => 
                           n2254, A => n2587, ZN => n2584);
   U3868 : AOI22_X1 port map( A1 => n2256, A2 => pc_lut_30_13_port, B1 => n2257
                           , B2 => pc_lut_31_13_port, ZN => n2587);
   U3871 : OAI221_X1 port map( B1 => n1698, B2 => n2258, C1 => n1664, C2 => 
                           n2259, A => n2588, ZN => n2583);
   U3872 : AOI22_X1 port map( A1 => n2261, A2 => pc_lut_18_13_port, B1 => n2262
                           , B2 => pc_lut_19_13_port, ZN => n2588);
   U3875 : OAI221_X1 port map( B1 => n1503, B2 => n2263, C1 => n1468, C2 => 
                           n2264, A => n2589, ZN => n2582);
   U3876 : AOI22_X1 port map( A1 => n2266, A2 => pc_lut_20_13_port, B1 => n2267
                           , B2 => pc_lut_21_13_port, ZN => n2589);
   U3879 : NOR4_X1 port map( A1 => n2590, A2 => n2591, A3 => n2592, A4 => n2593
                           , ZN => n2580);
   U3880 : OAI221_X1 port map( B1 => n1968, B2 => n2272, C1 => n1934, C2 => 
                           n2273, A => n2594, ZN => n2593);
   U3881 : AOI22_X1 port map( A1 => n2275, A2 => pc_lut_10_13_port, B1 => n2276
                           , B2 => pc_lut_11_13_port, ZN => n2594);
   U3884 : OAI221_X1 port map( B1 => n1833, B2 => n2277, C1 => n1799, C2 => 
                           n2278, A => n2595, ZN => n2592);
   U3885 : AOI22_X1 port map( A1 => n2280, A2 => pc_lut_14_13_port, B1 => n2281
                           , B2 => pc_lut_15_13_port, ZN => n2595);
   U3888 : OAI221_X1 port map( B1 => n2232, B2 => n2282, C1 => n2198, C2 => 
                           n2283, A => n2596, ZN => n2591);
   U3889 : AOI22_X1 port map( A1 => n2285, A2 => pc_lut_2_13_port, B1 => n2286,
                           B2 => pc_lut_3_13_port, ZN => n2596);
   U3892 : OAI221_X1 port map( B1 => n2100, B2 => n2287, C1 => n2066, C2 => 
                           n2288, A => n2597, ZN => n2590);
   U3893 : AOI22_X1 port map( A1 => n2290, A2 => pc_lut_6_13_port, B1 => n2291,
                           B2 => pc_lut_7_13_port, ZN => n2597);
   U3896 : NAND2_X1 port map( A1 => n2598, A2 => n2599, ZN => N205);
   U3897 : NOR4_X1 port map( A1 => n2600, A2 => n2601, A3 => n2602, A4 => n2603
                           , ZN => n2599);
   U3898 : OAI221_X1 port map( B1 => n1420, B2 => n2248, C1 => n1386, C2 => 
                           n2249, A => n2604, ZN => n2603);
   U3899 : AOI22_X1 port map( A1 => n2251, A2 => pc_lut_26_14_port, B1 => n2252
                           , B2 => pc_lut_27_14_port, ZN => n2604);
   U3902 : OAI221_X1 port map( B1 => n1285, B2 => n2253, C1 => n1250, C2 => 
                           n2254, A => n2605, ZN => n2602);
   U3903 : AOI22_X1 port map( A1 => n2256, A2 => pc_lut_30_14_port, B1 => n2257
                           , B2 => pc_lut_31_14_port, ZN => n2605);
   U3906 : OAI221_X1 port map( B1 => n1684, B2 => n2258, C1 => n1650, C2 => 
                           n2259, A => n2606, ZN => n2601);
   U3907 : AOI22_X1 port map( A1 => n2261, A2 => pc_lut_18_14_port, B1 => n2262
                           , B2 => pc_lut_19_14_port, ZN => n2606);
   U3910 : OAI221_X1 port map( B1 => n1489, B2 => n2263, C1 => n1454, C2 => 
                           n2264, A => n2607, ZN => n2600);
   U3911 : AOI22_X1 port map( A1 => n2266, A2 => pc_lut_20_14_port, B1 => n2267
                           , B2 => pc_lut_21_14_port, ZN => n2607);
   U3914 : NOR4_X1 port map( A1 => n2608, A2 => n2609, A3 => n2610, A4 => n2611
                           , ZN => n2598);
   U3915 : OAI221_X1 port map( B1 => n1954, B2 => n2272, C1 => n1920, C2 => 
                           n2273, A => n2612, ZN => n2611);
   U3916 : AOI22_X1 port map( A1 => n2275, A2 => pc_lut_10_14_port, B1 => n2276
                           , B2 => pc_lut_11_14_port, ZN => n2612);
   U3919 : OAI221_X1 port map( B1 => n1819, B2 => n2277, C1 => n1785, C2 => 
                           n2278, A => n2613, ZN => n2610);
   U3920 : AOI22_X1 port map( A1 => n2280, A2 => pc_lut_14_14_port, B1 => n2281
                           , B2 => pc_lut_15_14_port, ZN => n2613);
   U3923 : OAI221_X1 port map( B1 => n2218, B2 => n2282, C1 => n2184, C2 => 
                           n2283, A => n2614, ZN => n2609);
   U3924 : AOI22_X1 port map( A1 => n2285, A2 => pc_lut_2_14_port, B1 => n2286,
                           B2 => pc_lut_3_14_port, ZN => n2614);
   U3927 : OAI221_X1 port map( B1 => n2086, B2 => n2287, C1 => n2052, C2 => 
                           n2288, A => n2615, ZN => n2608);
   U3928 : AOI22_X1 port map( A1 => n2290, A2 => pc_lut_6_14_port, B1 => n2291,
                           B2 => pc_lut_7_14_port, ZN => n2615);
   U3931 : NAND2_X1 port map( A1 => n2616, A2 => n2617, ZN => N204);
   U3932 : NOR4_X1 port map( A1 => n2618, A2 => n2619, A3 => n2620, A4 => n2621
                           , ZN => n2617);
   U3933 : OAI221_X1 port map( B1 => n1435, B2 => n2248, C1 => n1401, C2 => 
                           n2249, A => n2622, ZN => n2621);
   U3934 : AOI22_X1 port map( A1 => n2251, A2 => pc_lut_26_15_port, B1 => n2252
                           , B2 => pc_lut_27_15_port, ZN => n2622);
   U3937 : OAI221_X1 port map( B1 => n1300, B2 => n2253, C1 => n1266, C2 => 
                           n2254, A => n2623, ZN => n2620);
   U3938 : AOI22_X1 port map( A1 => n2256, A2 => pc_lut_30_15_port, B1 => n2257
                           , B2 => pc_lut_31_15_port, ZN => n2623);
   U3941 : OAI221_X1 port map( B1 => n1699, B2 => n2258, C1 => n1665, C2 => 
                           n2259, A => n2624, ZN => n2619);
   U3942 : AOI22_X1 port map( A1 => n2261, A2 => pc_lut_18_15_port, B1 => n2262
                           , B2 => pc_lut_19_15_port, ZN => n2624);
   U3945 : OAI221_X1 port map( B1 => n1504, B2 => n2263, C1 => n1469, C2 => 
                           n2264, A => n2625, ZN => n2618);
   U3946 : AOI22_X1 port map( A1 => n2266, A2 => pc_lut_20_15_port, B1 => n2267
                           , B2 => pc_lut_21_15_port, ZN => n2625);
   U3949 : NOR4_X1 port map( A1 => n2626, A2 => n2627, A3 => n2628, A4 => n2629
                           , ZN => n2616);
   U3950 : OAI221_X1 port map( B1 => n1969, B2 => n2272, C1 => n1935, C2 => 
                           n2273, A => n2630, ZN => n2629);
   U3951 : AOI22_X1 port map( A1 => n2275, A2 => pc_lut_10_15_port, B1 => n2276
                           , B2 => pc_lut_11_15_port, ZN => n2630);
   U3954 : OAI221_X1 port map( B1 => n1834, B2 => n2277, C1 => n1800, C2 => 
                           n2278, A => n2631, ZN => n2628);
   U3955 : AOI22_X1 port map( A1 => n2280, A2 => pc_lut_14_15_port, B1 => n2281
                           , B2 => pc_lut_15_15_port, ZN => n2631);
   U3958 : OAI221_X1 port map( B1 => n2233, B2 => n2282, C1 => n2199, C2 => 
                           n2283, A => n2632, ZN => n2627);
   U3959 : AOI22_X1 port map( A1 => n2285, A2 => pc_lut_2_15_port, B1 => n2286,
                           B2 => pc_lut_3_15_port, ZN => n2632);
   U3962 : OAI221_X1 port map( B1 => n2101, B2 => n2287, C1 => n2067, C2 => 
                           n2288, A => n2633, ZN => n2626);
   U3963 : AOI22_X1 port map( A1 => n2290, A2 => pc_lut_6_15_port, B1 => n2291,
                           B2 => pc_lut_7_15_port, ZN => n2633);
   U3966 : NAND2_X1 port map( A1 => n2634, A2 => n2635, ZN => N203);
   U3967 : NOR4_X1 port map( A1 => n2636, A2 => n2637, A3 => n2638, A4 => n2639
                           , ZN => n2635);
   U3968 : OAI221_X1 port map( B1 => n1419, B2 => n2248, C1 => n1385, C2 => 
                           n2249, A => n2640, ZN => n2639);
   U3969 : AOI22_X1 port map( A1 => n2251, A2 => pc_lut_26_16_port, B1 => n2252
                           , B2 => pc_lut_27_16_port, ZN => n2640);
   U3972 : OAI221_X1 port map( B1 => n1284, B2 => n2253, C1 => n1249, C2 => 
                           n2254, A => n2641, ZN => n2638);
   U3973 : AOI22_X1 port map( A1 => n2256, A2 => pc_lut_30_16_port, B1 => n2257
                           , B2 => pc_lut_31_16_port, ZN => n2641);
   U3976 : OAI221_X1 port map( B1 => n1683, B2 => n2258, C1 => n1649, C2 => 
                           n2259, A => n2642, ZN => n2637);
   U3977 : AOI22_X1 port map( A1 => n2261, A2 => pc_lut_18_16_port, B1 => n2262
                           , B2 => pc_lut_19_16_port, ZN => n2642);
   U3980 : OAI221_X1 port map( B1 => n1488, B2 => n2263, C1 => n1453, C2 => 
                           n2264, A => n2643, ZN => n2636);
   U3981 : AOI22_X1 port map( A1 => n2266, A2 => pc_lut_20_16_port, B1 => n2267
                           , B2 => pc_lut_21_16_port, ZN => n2643);
   U3984 : NOR4_X1 port map( A1 => n2644, A2 => n2645, A3 => n2646, A4 => n2647
                           , ZN => n2634);
   U3985 : OAI221_X1 port map( B1 => n1953, B2 => n2272, C1 => n1919, C2 => 
                           n2273, A => n2648, ZN => n2647);
   U3986 : AOI22_X1 port map( A1 => n2275, A2 => pc_lut_10_16_port, B1 => n2276
                           , B2 => pc_lut_11_16_port, ZN => n2648);
   U3989 : OAI221_X1 port map( B1 => n1818, B2 => n2277, C1 => n1784, C2 => 
                           n2278, A => n2649, ZN => n2646);
   U3990 : AOI22_X1 port map( A1 => n2280, A2 => pc_lut_14_16_port, B1 => n2281
                           , B2 => pc_lut_15_16_port, ZN => n2649);
   U3993 : OAI221_X1 port map( B1 => n2217, B2 => n2282, C1 => n2183, C2 => 
                           n2283, A => n2650, ZN => n2645);
   U3994 : AOI22_X1 port map( A1 => n2285, A2 => pc_lut_2_16_port, B1 => n2286,
                           B2 => pc_lut_3_16_port, ZN => n2650);
   U3997 : OAI221_X1 port map( B1 => n2085, B2 => n2287, C1 => n2051, C2 => 
                           n2288, A => n2651, ZN => n2644);
   U3998 : AOI22_X1 port map( A1 => n2290, A2 => pc_lut_6_16_port, B1 => n2291,
                           B2 => pc_lut_7_16_port, ZN => n2651);
   U4001 : NAND2_X1 port map( A1 => n2652, A2 => n2653, ZN => N202);
   U4002 : NOR4_X1 port map( A1 => n2654, A2 => n2655, A3 => n2656, A4 => n2657
                           , ZN => n2653);
   U4003 : OAI221_X1 port map( B1 => n1436, B2 => n2248, C1 => n1402, C2 => 
                           n2249, A => n2658, ZN => n2657);
   U4004 : AOI22_X1 port map( A1 => n2251, A2 => pc_lut_26_17_port, B1 => n2252
                           , B2 => pc_lut_27_17_port, ZN => n2658);
   U4007 : OAI221_X1 port map( B1 => n1301, B2 => n2253, C1 => n1267, C2 => 
                           n2254, A => n2659, ZN => n2656);
   U4008 : AOI22_X1 port map( A1 => n2256, A2 => pc_lut_30_17_port, B1 => n2257
                           , B2 => pc_lut_31_17_port, ZN => n2659);
   U4011 : OAI221_X1 port map( B1 => n1700, B2 => n2258, C1 => n1666, C2 => 
                           n2259, A => n2660, ZN => n2655);
   U4012 : AOI22_X1 port map( A1 => n2261, A2 => pc_lut_18_17_port, B1 => n2262
                           , B2 => pc_lut_19_17_port, ZN => n2660);
   U4015 : OAI221_X1 port map( B1 => n1505, B2 => n2263, C1 => n1470, C2 => 
                           n2264, A => n2661, ZN => n2654);
   U4016 : AOI22_X1 port map( A1 => n2266, A2 => pc_lut_20_17_port, B1 => n2267
                           , B2 => pc_lut_21_17_port, ZN => n2661);
   U4019 : NOR4_X1 port map( A1 => n2662, A2 => n2663, A3 => n2664, A4 => n2665
                           , ZN => n2652);
   U4020 : OAI221_X1 port map( B1 => n1970, B2 => n2272, C1 => n1936, C2 => 
                           n2273, A => n2666, ZN => n2665);
   U4021 : AOI22_X1 port map( A1 => n2275, A2 => pc_lut_10_17_port, B1 => n2276
                           , B2 => pc_lut_11_17_port, ZN => n2666);
   U4024 : OAI221_X1 port map( B1 => n1835, B2 => n2277, C1 => n1801, C2 => 
                           n2278, A => n2667, ZN => n2664);
   U4025 : AOI22_X1 port map( A1 => n2280, A2 => pc_lut_14_17_port, B1 => n2281
                           , B2 => pc_lut_15_17_port, ZN => n2667);
   U4028 : OAI221_X1 port map( B1 => n2234, B2 => n2282, C1 => n2200, C2 => 
                           n2283, A => n2668, ZN => n2663);
   U4029 : AOI22_X1 port map( A1 => n2285, A2 => pc_lut_2_17_port, B1 => n2286,
                           B2 => pc_lut_3_17_port, ZN => n2668);
   U4032 : OAI221_X1 port map( B1 => n2102, B2 => n2287, C1 => n2068, C2 => 
                           n2288, A => n2669, ZN => n2662);
   U4033 : AOI22_X1 port map( A1 => n2290, A2 => pc_lut_6_17_port, B1 => n2291,
                           B2 => pc_lut_7_17_port, ZN => n2669);
   U4036 : NAND2_X1 port map( A1 => n2670, A2 => n2671, ZN => N201);
   U4037 : NOR4_X1 port map( A1 => n2672, A2 => n2673, A3 => n2674, A4 => n2675
                           , ZN => n2671);
   U4038 : OAI221_X1 port map( B1 => n1418, B2 => n2248, C1 => n1384, C2 => 
                           n2249, A => n2676, ZN => n2675);
   U4039 : AOI22_X1 port map( A1 => n2251, A2 => pc_lut_26_18_port, B1 => n2252
                           , B2 => pc_lut_27_18_port, ZN => n2676);
   U4042 : OAI221_X1 port map( B1 => n1283, B2 => n2253, C1 => n1248, C2 => 
                           n2254, A => n2677, ZN => n2674);
   U4043 : AOI22_X1 port map( A1 => n2256, A2 => pc_lut_30_18_port, B1 => n2257
                           , B2 => pc_lut_31_18_port, ZN => n2677);
   U4046 : OAI221_X1 port map( B1 => n1682, B2 => n2258, C1 => n1648, C2 => 
                           n2259, A => n2678, ZN => n2673);
   U4047 : AOI22_X1 port map( A1 => n2261, A2 => pc_lut_18_18_port, B1 => n2262
                           , B2 => pc_lut_19_18_port, ZN => n2678);
   U4050 : OAI221_X1 port map( B1 => n1487, B2 => n2263, C1 => n1452, C2 => 
                           n2264, A => n2679, ZN => n2672);
   U4051 : AOI22_X1 port map( A1 => n2266, A2 => pc_lut_20_18_port, B1 => n2267
                           , B2 => pc_lut_21_18_port, ZN => n2679);
   U4054 : NOR4_X1 port map( A1 => n2680, A2 => n2681, A3 => n2682, A4 => n2683
                           , ZN => n2670);
   U4055 : OAI221_X1 port map( B1 => n1952, B2 => n2272, C1 => n1918, C2 => 
                           n2273, A => n2684, ZN => n2683);
   U4056 : AOI22_X1 port map( A1 => n2275, A2 => pc_lut_10_18_port, B1 => n2276
                           , B2 => pc_lut_11_18_port, ZN => n2684);
   U4059 : OAI221_X1 port map( B1 => n1817, B2 => n2277, C1 => n1783, C2 => 
                           n2278, A => n2685, ZN => n2682);
   U4060 : AOI22_X1 port map( A1 => n2280, A2 => pc_lut_14_18_port, B1 => n2281
                           , B2 => pc_lut_15_18_port, ZN => n2685);
   U4063 : OAI221_X1 port map( B1 => n2216, B2 => n2282, C1 => n2182, C2 => 
                           n2283, A => n2686, ZN => n2681);
   U4064 : AOI22_X1 port map( A1 => n2285, A2 => pc_lut_2_18_port, B1 => n2286,
                           B2 => pc_lut_3_18_port, ZN => n2686);
   U4067 : OAI221_X1 port map( B1 => n2084, B2 => n2287, C1 => n2050, C2 => 
                           n2288, A => n2687, ZN => n2680);
   U4068 : AOI22_X1 port map( A1 => n2290, A2 => pc_lut_6_18_port, B1 => n2291,
                           B2 => pc_lut_7_18_port, ZN => n2687);
   U4071 : NAND2_X1 port map( A1 => n2688, A2 => n2689, ZN => N200);
   U4072 : NOR4_X1 port map( A1 => n2690, A2 => n2691, A3 => n2692, A4 => n2693
                           , ZN => n2689);
   U4073 : OAI221_X1 port map( B1 => n1437, B2 => n2248, C1 => n1403, C2 => 
                           n2249, A => n2694, ZN => n2693);
   U4074 : AOI22_X1 port map( A1 => n2251, A2 => pc_lut_26_19_port, B1 => n2252
                           , B2 => pc_lut_27_19_port, ZN => n2694);
   U4077 : OAI221_X1 port map( B1 => n1302, B2 => n2253, C1 => n1268, C2 => 
                           n2254, A => n2695, ZN => n2692);
   U4078 : AOI22_X1 port map( A1 => n2256, A2 => pc_lut_30_19_port, B1 => n2257
                           , B2 => pc_lut_31_19_port, ZN => n2695);
   U4081 : OAI221_X1 port map( B1 => n1701, B2 => n2258, C1 => n1667, C2 => 
                           n2259, A => n2696, ZN => n2691);
   U4082 : AOI22_X1 port map( A1 => n2261, A2 => pc_lut_18_19_port, B1 => n2262
                           , B2 => pc_lut_19_19_port, ZN => n2696);
   U4085 : OAI221_X1 port map( B1 => n1506, B2 => n2263, C1 => n1471, C2 => 
                           n2264, A => n2697, ZN => n2690);
   U4086 : AOI22_X1 port map( A1 => n2266, A2 => pc_lut_20_19_port, B1 => n2267
                           , B2 => pc_lut_21_19_port, ZN => n2697);
   U4089 : NOR4_X1 port map( A1 => n2698, A2 => n2699, A3 => n2700, A4 => n2701
                           , ZN => n2688);
   U4090 : OAI221_X1 port map( B1 => n1971, B2 => n2272, C1 => n1937, C2 => 
                           n2273, A => n2702, ZN => n2701);
   U4091 : AOI22_X1 port map( A1 => n2275, A2 => pc_lut_10_19_port, B1 => n2276
                           , B2 => pc_lut_11_19_port, ZN => n2702);
   U4094 : OAI221_X1 port map( B1 => n1836, B2 => n2277, C1 => n1802, C2 => 
                           n2278, A => n2703, ZN => n2700);
   U4095 : AOI22_X1 port map( A1 => n2280, A2 => pc_lut_14_19_port, B1 => n2281
                           , B2 => pc_lut_15_19_port, ZN => n2703);
   U4098 : OAI221_X1 port map( B1 => n2235, B2 => n2282, C1 => n2201, C2 => 
                           n2283, A => n2704, ZN => n2699);
   U4099 : AOI22_X1 port map( A1 => n2285, A2 => pc_lut_2_19_port, B1 => n2286,
                           B2 => pc_lut_3_19_port, ZN => n2704);
   U4102 : OAI221_X1 port map( B1 => n2103, B2 => n2287, C1 => n2069, C2 => 
                           n2288, A => n2705, ZN => n2698);
   U4103 : AOI22_X1 port map( A1 => n2290, A2 => pc_lut_6_19_port, B1 => n2291,
                           B2 => pc_lut_7_19_port, ZN => n2705);
   U4106 : NAND2_X1 port map( A1 => n2706, A2 => n2707, ZN => N199);
   U4107 : NOR4_X1 port map( A1 => n2708, A2 => n2709, A3 => n2710, A4 => n2711
                           , ZN => n2707);
   U4108 : OAI221_X1 port map( B1 => n1417, B2 => n2248, C1 => n1383, C2 => 
                           n2249, A => n2712, ZN => n2711);
   U4109 : AOI22_X1 port map( A1 => n2251, A2 => pc_lut_26_20_port, B1 => n2252
                           , B2 => pc_lut_27_20_port, ZN => n2712);
   U4112 : OAI221_X1 port map( B1 => n1282, B2 => n2253, C1 => n1247, C2 => 
                           n2254, A => n2713, ZN => n2710);
   U4113 : AOI22_X1 port map( A1 => n2256, A2 => pc_lut_30_20_port, B1 => n2257
                           , B2 => pc_lut_31_20_port, ZN => n2713);
   U4116 : OAI221_X1 port map( B1 => n1681, B2 => n2258, C1 => n1647, C2 => 
                           n2259, A => n2714, ZN => n2709);
   U4117 : AOI22_X1 port map( A1 => n2261, A2 => pc_lut_18_20_port, B1 => n2262
                           , B2 => pc_lut_19_20_port, ZN => n2714);
   U4120 : OAI221_X1 port map( B1 => n1486, B2 => n2263, C1 => n1451, C2 => 
                           n2264, A => n2715, ZN => n2708);
   U4121 : AOI22_X1 port map( A1 => n2266, A2 => pc_lut_20_20_port, B1 => n2267
                           , B2 => pc_lut_21_20_port, ZN => n2715);
   U4124 : NOR4_X1 port map( A1 => n2716, A2 => n2717, A3 => n2718, A4 => n2719
                           , ZN => n2706);
   U4125 : OAI221_X1 port map( B1 => n1951, B2 => n2272, C1 => n1917, C2 => 
                           n2273, A => n2720, ZN => n2719);
   U4126 : AOI22_X1 port map( A1 => n2275, A2 => pc_lut_10_20_port, B1 => n2276
                           , B2 => pc_lut_11_20_port, ZN => n2720);
   U4129 : OAI221_X1 port map( B1 => n1816, B2 => n2277, C1 => n1782, C2 => 
                           n2278, A => n2721, ZN => n2718);
   U4130 : AOI22_X1 port map( A1 => n2280, A2 => pc_lut_14_20_port, B1 => n2281
                           , B2 => pc_lut_15_20_port, ZN => n2721);
   U4133 : OAI221_X1 port map( B1 => n2215, B2 => n2282, C1 => n2181, C2 => 
                           n2283, A => n2722, ZN => n2717);
   U4134 : AOI22_X1 port map( A1 => n2285, A2 => pc_lut_2_20_port, B1 => n2286,
                           B2 => pc_lut_3_20_port, ZN => n2722);
   U4137 : OAI221_X1 port map( B1 => n2083, B2 => n2287, C1 => n2049, C2 => 
                           n2288, A => n2723, ZN => n2716);
   U4138 : AOI22_X1 port map( A1 => n2290, A2 => pc_lut_6_20_port, B1 => n2291,
                           B2 => pc_lut_7_20_port, ZN => n2723);
   U4141 : NAND2_X1 port map( A1 => n2724, A2 => n2725, ZN => N198);
   U4142 : NOR4_X1 port map( A1 => n2726, A2 => n2727, A3 => n2728, A4 => n2729
                           , ZN => n2725);
   U4143 : OAI221_X1 port map( B1 => n1438, B2 => n2248, C1 => n1404, C2 => 
                           n2249, A => n2730, ZN => n2729);
   U4144 : AOI22_X1 port map( A1 => n2251, A2 => pc_lut_26_21_port, B1 => n2252
                           , B2 => pc_lut_27_21_port, ZN => n2730);
   U4147 : OAI221_X1 port map( B1 => n1303, B2 => n2253, C1 => n1269, C2 => 
                           n2254, A => n2731, ZN => n2728);
   U4148 : AOI22_X1 port map( A1 => n2256, A2 => pc_lut_30_21_port, B1 => n2257
                           , B2 => pc_lut_31_21_port, ZN => n2731);
   U4151 : OAI221_X1 port map( B1 => n1702, B2 => n2258, C1 => n1668, C2 => 
                           n2259, A => n2732, ZN => n2727);
   U4152 : AOI22_X1 port map( A1 => n2261, A2 => pc_lut_18_21_port, B1 => n2262
                           , B2 => pc_lut_19_21_port, ZN => n2732);
   U4155 : OAI221_X1 port map( B1 => n1507, B2 => n2263, C1 => n1472, C2 => 
                           n2264, A => n2733, ZN => n2726);
   U4156 : AOI22_X1 port map( A1 => n2266, A2 => pc_lut_20_21_port, B1 => n2267
                           , B2 => pc_lut_21_21_port, ZN => n2733);
   U4159 : NOR4_X1 port map( A1 => n2734, A2 => n2735, A3 => n2736, A4 => n2737
                           , ZN => n2724);
   U4160 : OAI221_X1 port map( B1 => n1972, B2 => n2272, C1 => n1938, C2 => 
                           n2273, A => n2738, ZN => n2737);
   U4161 : AOI22_X1 port map( A1 => n2275, A2 => pc_lut_10_21_port, B1 => n2276
                           , B2 => pc_lut_11_21_port, ZN => n2738);
   U4164 : OAI221_X1 port map( B1 => n1837, B2 => n2277, C1 => n1803, C2 => 
                           n2278, A => n2739, ZN => n2736);
   U4165 : AOI22_X1 port map( A1 => n2280, A2 => pc_lut_14_21_port, B1 => n2281
                           , B2 => pc_lut_15_21_port, ZN => n2739);
   U4168 : OAI221_X1 port map( B1 => n2236, B2 => n2282, C1 => n2202, C2 => 
                           n2283, A => n2740, ZN => n2735);
   U4169 : AOI22_X1 port map( A1 => n2285, A2 => pc_lut_2_21_port, B1 => n2286,
                           B2 => pc_lut_3_21_port, ZN => n2740);
   U4172 : OAI221_X1 port map( B1 => n2104, B2 => n2287, C1 => n2070, C2 => 
                           n2288, A => n2741, ZN => n2734);
   U4173 : AOI22_X1 port map( A1 => n2290, A2 => pc_lut_6_21_port, B1 => n2291,
                           B2 => pc_lut_7_21_port, ZN => n2741);
   U4176 : NAND2_X1 port map( A1 => n2742, A2 => n2743, ZN => N197);
   U4177 : NOR4_X1 port map( A1 => n2744, A2 => n2745, A3 => n2746, A4 => n2747
                           , ZN => n2743);
   U4178 : OAI221_X1 port map( B1 => n1416, B2 => n2248, C1 => n1382, C2 => 
                           n2249, A => n2748, ZN => n2747);
   U4179 : AOI22_X1 port map( A1 => n2251, A2 => pc_lut_26_22_port, B1 => n2252
                           , B2 => pc_lut_27_22_port, ZN => n2748);
   U4182 : OAI221_X1 port map( B1 => n1281, B2 => n2253, C1 => n1246, C2 => 
                           n2254, A => n2749, ZN => n2746);
   U4183 : AOI22_X1 port map( A1 => n2256, A2 => pc_lut_30_22_port, B1 => n2257
                           , B2 => pc_lut_31_22_port, ZN => n2749);
   U4186 : OAI221_X1 port map( B1 => n1680, B2 => n2258, C1 => n1646, C2 => 
                           n2259, A => n2750, ZN => n2745);
   U4187 : AOI22_X1 port map( A1 => n2261, A2 => pc_lut_18_22_port, B1 => n2262
                           , B2 => pc_lut_19_22_port, ZN => n2750);
   U4190 : OAI221_X1 port map( B1 => n1485, B2 => n2263, C1 => n1450, C2 => 
                           n2264, A => n2751, ZN => n2744);
   U4191 : AOI22_X1 port map( A1 => n2266, A2 => pc_lut_20_22_port, B1 => n2267
                           , B2 => pc_lut_21_22_port, ZN => n2751);
   U4194 : NOR4_X1 port map( A1 => n2752, A2 => n2753, A3 => n2754, A4 => n2755
                           , ZN => n2742);
   U4195 : OAI221_X1 port map( B1 => n1950, B2 => n2272, C1 => n1916, C2 => 
                           n2273, A => n2756, ZN => n2755);
   U4196 : AOI22_X1 port map( A1 => n2275, A2 => pc_lut_10_22_port, B1 => n2276
                           , B2 => pc_lut_11_22_port, ZN => n2756);
   U4199 : OAI221_X1 port map( B1 => n1815, B2 => n2277, C1 => n1781, C2 => 
                           n2278, A => n2757, ZN => n2754);
   U4200 : AOI22_X1 port map( A1 => n2280, A2 => pc_lut_14_22_port, B1 => n2281
                           , B2 => pc_lut_15_22_port, ZN => n2757);
   U4203 : OAI221_X1 port map( B1 => n2214, B2 => n2282, C1 => n2180, C2 => 
                           n2283, A => n2758, ZN => n2753);
   U4204 : AOI22_X1 port map( A1 => n2285, A2 => pc_lut_2_22_port, B1 => n2286,
                           B2 => pc_lut_3_22_port, ZN => n2758);
   U4207 : OAI221_X1 port map( B1 => n2082, B2 => n2287, C1 => n2048, C2 => 
                           n2288, A => n2759, ZN => n2752);
   U4208 : AOI22_X1 port map( A1 => n2290, A2 => pc_lut_6_22_port, B1 => n2291,
                           B2 => pc_lut_7_22_port, ZN => n2759);
   U4211 : NAND2_X1 port map( A1 => n2760, A2 => n2761, ZN => N196);
   U4212 : NOR4_X1 port map( A1 => n2762, A2 => n2763, A3 => n2764, A4 => n2765
                           , ZN => n2761);
   U4213 : OAI221_X1 port map( B1 => n1439, B2 => n2248, C1 => n1405, C2 => 
                           n2249, A => n2766, ZN => n2765);
   U4214 : AOI22_X1 port map( A1 => n2251, A2 => pc_lut_26_23_port, B1 => n2252
                           , B2 => pc_lut_27_23_port, ZN => n2766);
   U4217 : OAI221_X1 port map( B1 => n1304, B2 => n2253, C1 => n1270, C2 => 
                           n2254, A => n2767, ZN => n2764);
   U4218 : AOI22_X1 port map( A1 => n2256, A2 => pc_lut_30_23_port, B1 => n2257
                           , B2 => pc_lut_31_23_port, ZN => n2767);
   U4221 : OAI221_X1 port map( B1 => n1703, B2 => n2258, C1 => n1669, C2 => 
                           n2259, A => n2768, ZN => n2763);
   U4222 : AOI22_X1 port map( A1 => n2261, A2 => pc_lut_18_23_port, B1 => n2262
                           , B2 => pc_lut_19_23_port, ZN => n2768);
   U4225 : OAI221_X1 port map( B1 => n1508, B2 => n2263, C1 => n1473, C2 => 
                           n2264, A => n2769, ZN => n2762);
   U4226 : AOI22_X1 port map( A1 => n2266, A2 => pc_lut_20_23_port, B1 => n2267
                           , B2 => pc_lut_21_23_port, ZN => n2769);
   U4229 : NOR4_X1 port map( A1 => n2770, A2 => n2771, A3 => n2772, A4 => n2773
                           , ZN => n2760);
   U4230 : OAI221_X1 port map( B1 => n1973, B2 => n2272, C1 => n1939, C2 => 
                           n2273, A => n2774, ZN => n2773);
   U4231 : AOI22_X1 port map( A1 => n2275, A2 => pc_lut_10_23_port, B1 => n2276
                           , B2 => pc_lut_11_23_port, ZN => n2774);
   U4234 : OAI221_X1 port map( B1 => n1838, B2 => n2277, C1 => n1804, C2 => 
                           n2278, A => n2775, ZN => n2772);
   U4235 : AOI22_X1 port map( A1 => n2280, A2 => pc_lut_14_23_port, B1 => n2281
                           , B2 => pc_lut_15_23_port, ZN => n2775);
   U4238 : OAI221_X1 port map( B1 => n2237, B2 => n2282, C1 => n2203, C2 => 
                           n2283, A => n2776, ZN => n2771);
   U4239 : AOI22_X1 port map( A1 => n2285, A2 => pc_lut_2_23_port, B1 => n2286,
                           B2 => pc_lut_3_23_port, ZN => n2776);
   U4242 : OAI221_X1 port map( B1 => n2105, B2 => n2287, C1 => n2071, C2 => 
                           n2288, A => n2777, ZN => n2770);
   U4243 : AOI22_X1 port map( A1 => n2290, A2 => pc_lut_6_23_port, B1 => n2291,
                           B2 => pc_lut_7_23_port, ZN => n2777);
   U4246 : NAND2_X1 port map( A1 => n2778, A2 => n2779, ZN => N195);
   U4247 : NOR4_X1 port map( A1 => n2780, A2 => n2781, A3 => n2782, A4 => n2783
                           , ZN => n2779);
   U4248 : OAI221_X1 port map( B1 => n1415, B2 => n2248, C1 => n1381, C2 => 
                           n2249, A => n2784, ZN => n2783);
   U4249 : AOI22_X1 port map( A1 => n2251, A2 => pc_lut_26_24_port, B1 => n2252
                           , B2 => pc_lut_27_24_port, ZN => n2784);
   U4252 : OAI221_X1 port map( B1 => n1280, B2 => n2253, C1 => n1245, C2 => 
                           n2254, A => n2785, ZN => n2782);
   U4253 : AOI22_X1 port map( A1 => n2256, A2 => pc_lut_30_24_port, B1 => n2257
                           , B2 => pc_lut_31_24_port, ZN => n2785);
   U4256 : OAI221_X1 port map( B1 => n1679, B2 => n2258, C1 => n1645, C2 => 
                           n2259, A => n2786, ZN => n2781);
   U4257 : AOI22_X1 port map( A1 => n2261, A2 => pc_lut_18_24_port, B1 => n2262
                           , B2 => pc_lut_19_24_port, ZN => n2786);
   U4260 : OAI221_X1 port map( B1 => n1484, B2 => n2263, C1 => n1449, C2 => 
                           n2264, A => n2787, ZN => n2780);
   U4261 : AOI22_X1 port map( A1 => n2266, A2 => pc_lut_20_24_port, B1 => n2267
                           , B2 => pc_lut_21_24_port, ZN => n2787);
   U4264 : NOR4_X1 port map( A1 => n2788, A2 => n2789, A3 => n2790, A4 => n2791
                           , ZN => n2778);
   U4265 : OAI221_X1 port map( B1 => n1949, B2 => n2272, C1 => n1915, C2 => 
                           n2273, A => n2792, ZN => n2791);
   U4266 : AOI22_X1 port map( A1 => n2275, A2 => pc_lut_10_24_port, B1 => n2276
                           , B2 => pc_lut_11_24_port, ZN => n2792);
   U4269 : OAI221_X1 port map( B1 => n1814, B2 => n2277, C1 => n1780, C2 => 
                           n2278, A => n2793, ZN => n2790);
   U4270 : AOI22_X1 port map( A1 => n2280, A2 => pc_lut_14_24_port, B1 => n2281
                           , B2 => pc_lut_15_24_port, ZN => n2793);
   U4273 : OAI221_X1 port map( B1 => n2213, B2 => n2282, C1 => n2179, C2 => 
                           n2283, A => n2794, ZN => n2789);
   U4274 : AOI22_X1 port map( A1 => n2285, A2 => pc_lut_2_24_port, B1 => n2286,
                           B2 => pc_lut_3_24_port, ZN => n2794);
   U4277 : OAI221_X1 port map( B1 => n2081, B2 => n2287, C1 => n2047, C2 => 
                           n2288, A => n2795, ZN => n2788);
   U4278 : AOI22_X1 port map( A1 => n2290, A2 => pc_lut_6_24_port, B1 => n2291,
                           B2 => pc_lut_7_24_port, ZN => n2795);
   U4281 : NAND2_X1 port map( A1 => n2796, A2 => n2797, ZN => N194);
   U4282 : NOR4_X1 port map( A1 => n2798, A2 => n2799, A3 => n2800, A4 => n2801
                           , ZN => n2797);
   U4283 : OAI221_X1 port map( B1 => n1440, B2 => n2248, C1 => n1406, C2 => 
                           n2249, A => n2802, ZN => n2801);
   U4284 : AOI22_X1 port map( A1 => n2251, A2 => pc_lut_26_25_port, B1 => n2252
                           , B2 => pc_lut_27_25_port, ZN => n2802);
   U4287 : OAI221_X1 port map( B1 => n1305, B2 => n2253, C1 => n1271, C2 => 
                           n2254, A => n2803, ZN => n2800);
   U4288 : AOI22_X1 port map( A1 => n2256, A2 => pc_lut_30_25_port, B1 => n2257
                           , B2 => pc_lut_31_25_port, ZN => n2803);
   U4291 : OAI221_X1 port map( B1 => n1704, B2 => n2258, C1 => n1670, C2 => 
                           n2259, A => n2804, ZN => n2799);
   U4292 : AOI22_X1 port map( A1 => n2261, A2 => pc_lut_18_25_port, B1 => n2262
                           , B2 => pc_lut_19_25_port, ZN => n2804);
   U4295 : OAI221_X1 port map( B1 => n1509, B2 => n2263, C1 => n1474, C2 => 
                           n2264, A => n2805, ZN => n2798);
   U4296 : AOI22_X1 port map( A1 => n2266, A2 => pc_lut_20_25_port, B1 => n2267
                           , B2 => pc_lut_21_25_port, ZN => n2805);
   U4299 : NOR4_X1 port map( A1 => n2806, A2 => n2807, A3 => n2808, A4 => n2809
                           , ZN => n2796);
   U4300 : OAI221_X1 port map( B1 => n1974, B2 => n2272, C1 => n1940, C2 => 
                           n2273, A => n2810, ZN => n2809);
   U4301 : AOI22_X1 port map( A1 => n2275, A2 => pc_lut_10_25_port, B1 => n2276
                           , B2 => pc_lut_11_25_port, ZN => n2810);
   U4304 : OAI221_X1 port map( B1 => n1839, B2 => n2277, C1 => n1805, C2 => 
                           n2278, A => n2811, ZN => n2808);
   U4305 : AOI22_X1 port map( A1 => n2280, A2 => pc_lut_14_25_port, B1 => n2281
                           , B2 => pc_lut_15_25_port, ZN => n2811);
   U4308 : OAI221_X1 port map( B1 => n2238, B2 => n2282, C1 => n2204, C2 => 
                           n2283, A => n2812, ZN => n2807);
   U4309 : AOI22_X1 port map( A1 => n2285, A2 => pc_lut_2_25_port, B1 => n2286,
                           B2 => pc_lut_3_25_port, ZN => n2812);
   U4312 : OAI221_X1 port map( B1 => n2106, B2 => n2287, C1 => n2072, C2 => 
                           n2288, A => n2813, ZN => n2806);
   U4313 : AOI22_X1 port map( A1 => n2290, A2 => pc_lut_6_25_port, B1 => n2291,
                           B2 => pc_lut_7_25_port, ZN => n2813);
   U4316 : NAND2_X1 port map( A1 => n2814, A2 => n2815, ZN => N193);
   U4317 : NOR4_X1 port map( A1 => n2816, A2 => n2817, A3 => n2818, A4 => n2819
                           , ZN => n2815);
   U4318 : OAI221_X1 port map( B1 => n1414, B2 => n2248, C1 => n1380, C2 => 
                           n2249, A => n2820, ZN => n2819);
   U4319 : AOI22_X1 port map( A1 => n2251, A2 => pc_lut_26_26_port, B1 => n2252
                           , B2 => pc_lut_27_26_port, ZN => n2820);
   U4322 : OAI221_X1 port map( B1 => n1279, B2 => n2253, C1 => n1244, C2 => 
                           n2254, A => n2821, ZN => n2818);
   U4323 : AOI22_X1 port map( A1 => n2256, A2 => pc_lut_30_26_port, B1 => n2257
                           , B2 => pc_lut_31_26_port, ZN => n2821);
   U4326 : OAI221_X1 port map( B1 => n1678, B2 => n2258, C1 => n1644, C2 => 
                           n2259, A => n2822, ZN => n2817);
   U4327 : AOI22_X1 port map( A1 => n2261, A2 => pc_lut_18_26_port, B1 => n2262
                           , B2 => pc_lut_19_26_port, ZN => n2822);
   U4330 : OAI221_X1 port map( B1 => n1483, B2 => n2263, C1 => n1448, C2 => 
                           n2264, A => n2823, ZN => n2816);
   U4331 : AOI22_X1 port map( A1 => n2266, A2 => pc_lut_20_26_port, B1 => n2267
                           , B2 => pc_lut_21_26_port, ZN => n2823);
   U4334 : NOR4_X1 port map( A1 => n2824, A2 => n2825, A3 => n2826, A4 => n2827
                           , ZN => n2814);
   U4335 : OAI221_X1 port map( B1 => n1948, B2 => n2272, C1 => n1914, C2 => 
                           n2273, A => n2828, ZN => n2827);
   U4336 : AOI22_X1 port map( A1 => n2275, A2 => pc_lut_10_26_port, B1 => n2276
                           , B2 => pc_lut_11_26_port, ZN => n2828);
   U4339 : OAI221_X1 port map( B1 => n1813, B2 => n2277, C1 => n1779, C2 => 
                           n2278, A => n2829, ZN => n2826);
   U4340 : AOI22_X1 port map( A1 => n2280, A2 => pc_lut_14_26_port, B1 => n2281
                           , B2 => pc_lut_15_26_port, ZN => n2829);
   U4343 : OAI221_X1 port map( B1 => n2212, B2 => n2282, C1 => n2178, C2 => 
                           n2283, A => n2830, ZN => n2825);
   U4344 : AOI22_X1 port map( A1 => n2285, A2 => pc_lut_2_26_port, B1 => n2286,
                           B2 => pc_lut_3_26_port, ZN => n2830);
   U4347 : OAI221_X1 port map( B1 => n2080, B2 => n2287, C1 => n2046, C2 => 
                           n2288, A => n2831, ZN => n2824);
   U4348 : AOI22_X1 port map( A1 => n2290, A2 => pc_lut_6_26_port, B1 => n2291,
                           B2 => pc_lut_7_26_port, ZN => n2831);
   U4351 : NAND2_X1 port map( A1 => n2832, A2 => n2833, ZN => N192);
   U4352 : NOR4_X1 port map( A1 => n2834, A2 => n2835, A3 => n2836, A4 => n2837
                           , ZN => n2833);
   U4353 : OAI221_X1 port map( B1 => n1441, B2 => n2248, C1 => n1407, C2 => 
                           n2249, A => n2838, ZN => n2837);
   U4354 : AOI22_X1 port map( A1 => n2251, A2 => pc_lut_26_27_port, B1 => n2252
                           , B2 => pc_lut_27_27_port, ZN => n2838);
   U4357 : OAI221_X1 port map( B1 => n1306, B2 => n2253, C1 => n1272, C2 => 
                           n2254, A => n2839, ZN => n2836);
   U4358 : AOI22_X1 port map( A1 => n2256, A2 => pc_lut_30_27_port, B1 => n2257
                           , B2 => pc_lut_31_27_port, ZN => n2839);
   U4361 : OAI221_X1 port map( B1 => n1705, B2 => n2258, C1 => n1671, C2 => 
                           n2259, A => n2840, ZN => n2835);
   U4362 : AOI22_X1 port map( A1 => n2261, A2 => pc_lut_18_27_port, B1 => n2262
                           , B2 => pc_lut_19_27_port, ZN => n2840);
   U4365 : OAI221_X1 port map( B1 => n1510, B2 => n2263, C1 => n1475, C2 => 
                           n2264, A => n2841, ZN => n2834);
   U4366 : AOI22_X1 port map( A1 => n2266, A2 => pc_lut_20_27_port, B1 => n2267
                           , B2 => pc_lut_21_27_port, ZN => n2841);
   U4369 : NOR4_X1 port map( A1 => n2842, A2 => n2843, A3 => n2844, A4 => n2845
                           , ZN => n2832);
   U4370 : OAI221_X1 port map( B1 => n1975, B2 => n2272, C1 => n1941, C2 => 
                           n2273, A => n2846, ZN => n2845);
   U4371 : AOI22_X1 port map( A1 => n2275, A2 => pc_lut_10_27_port, B1 => n2276
                           , B2 => pc_lut_11_27_port, ZN => n2846);
   U4374 : OAI221_X1 port map( B1 => n1840, B2 => n2277, C1 => n1806, C2 => 
                           n2278, A => n2847, ZN => n2844);
   U4375 : AOI22_X1 port map( A1 => n2280, A2 => pc_lut_14_27_port, B1 => n2281
                           , B2 => pc_lut_15_27_port, ZN => n2847);
   U4378 : OAI221_X1 port map( B1 => n2239, B2 => n2282, C1 => n2205, C2 => 
                           n2283, A => n2848, ZN => n2843);
   U4379 : AOI22_X1 port map( A1 => n2285, A2 => pc_lut_2_27_port, B1 => n2286,
                           B2 => pc_lut_3_27_port, ZN => n2848);
   U4382 : OAI221_X1 port map( B1 => n2107, B2 => n2287, C1 => n2073, C2 => 
                           n2288, A => n2849, ZN => n2842);
   U4383 : AOI22_X1 port map( A1 => n2290, A2 => pc_lut_6_27_port, B1 => n2291,
                           B2 => pc_lut_7_27_port, ZN => n2849);
   U4386 : NAND2_X1 port map( A1 => n2850, A2 => n2851, ZN => N191);
   U4387 : NOR4_X1 port map( A1 => n2852, A2 => n2853, A3 => n2854, A4 => n2855
                           , ZN => n2851);
   U4388 : OAI221_X1 port map( B1 => n1413, B2 => n2248, C1 => n1379, C2 => 
                           n2249, A => n2856, ZN => n2855);
   U4389 : AOI22_X1 port map( A1 => n2251, A2 => pc_lut_26_28_port, B1 => n2252
                           , B2 => pc_lut_27_28_port, ZN => n2856);
   U4392 : OAI221_X1 port map( B1 => n1278, B2 => n2253, C1 => n1243, C2 => 
                           n2254, A => n2857, ZN => n2854);
   U4393 : AOI22_X1 port map( A1 => n2256, A2 => pc_lut_30_28_port, B1 => n2257
                           , B2 => pc_lut_31_28_port, ZN => n2857);
   U4396 : OAI221_X1 port map( B1 => n1677, B2 => n2258, C1 => n1643, C2 => 
                           n2259, A => n2858, ZN => n2853);
   U4397 : AOI22_X1 port map( A1 => n2261, A2 => pc_lut_18_28_port, B1 => n2262
                           , B2 => pc_lut_19_28_port, ZN => n2858);
   U4400 : OAI221_X1 port map( B1 => n1482, B2 => n2263, C1 => n1447, C2 => 
                           n2264, A => n2859, ZN => n2852);
   U4401 : AOI22_X1 port map( A1 => n2266, A2 => pc_lut_20_28_port, B1 => n2267
                           , B2 => pc_lut_21_28_port, ZN => n2859);
   U4404 : NOR4_X1 port map( A1 => n2860, A2 => n2861, A3 => n2862, A4 => n2863
                           , ZN => n2850);
   U4405 : OAI221_X1 port map( B1 => n1947, B2 => n2272, C1 => n1913, C2 => 
                           n2273, A => n2864, ZN => n2863);
   U4406 : AOI22_X1 port map( A1 => n2275, A2 => pc_lut_10_28_port, B1 => n2276
                           , B2 => pc_lut_11_28_port, ZN => n2864);
   U4409 : OAI221_X1 port map( B1 => n1812, B2 => n2277, C1 => n1778, C2 => 
                           n2278, A => n2865, ZN => n2862);
   U4410 : AOI22_X1 port map( A1 => n2280, A2 => pc_lut_14_28_port, B1 => n2281
                           , B2 => pc_lut_15_28_port, ZN => n2865);
   U4413 : OAI221_X1 port map( B1 => n2211, B2 => n2282, C1 => n2177, C2 => 
                           n2283, A => n2866, ZN => n2861);
   U4414 : AOI22_X1 port map( A1 => n2285, A2 => pc_lut_2_28_port, B1 => n2286,
                           B2 => pc_lut_3_28_port, ZN => n2866);
   U4417 : OAI221_X1 port map( B1 => n2079, B2 => n2287, C1 => n2045, C2 => 
                           n2288, A => n2867, ZN => n2860);
   U4418 : AOI22_X1 port map( A1 => n2290, A2 => pc_lut_6_28_port, B1 => n2291,
                           B2 => pc_lut_7_28_port, ZN => n2867);
   U4421 : NAND2_X1 port map( A1 => n2868, A2 => n2869, ZN => N190);
   U4422 : NOR4_X1 port map( A1 => n2870, A2 => n2871, A3 => n2872, A4 => n2873
                           , ZN => n2869);
   U4423 : OAI221_X1 port map( B1 => n1442, B2 => n2248, C1 => n1408, C2 => 
                           n2249, A => n2874, ZN => n2873);
   U4424 : AOI22_X1 port map( A1 => n2251, A2 => pc_lut_26_29_port, B1 => n2252
                           , B2 => pc_lut_27_29_port, ZN => n2874);
   U4427 : OAI221_X1 port map( B1 => n1307, B2 => n2253, C1 => n1273, C2 => 
                           n2254, A => n2875, ZN => n2872);
   U4428 : AOI22_X1 port map( A1 => n2256, A2 => pc_lut_30_29_port, B1 => n2257
                           , B2 => pc_lut_31_29_port, ZN => n2875);
   U4431 : OAI221_X1 port map( B1 => n1706, B2 => n2258, C1 => n1672, C2 => 
                           n2259, A => n2876, ZN => n2871);
   U4432 : AOI22_X1 port map( A1 => n2261, A2 => pc_lut_18_29_port, B1 => n2262
                           , B2 => pc_lut_19_29_port, ZN => n2876);
   U4435 : OAI221_X1 port map( B1 => n1511, B2 => n2263, C1 => n1476, C2 => 
                           n2264, A => n2877, ZN => n2870);
   U4436 : AOI22_X1 port map( A1 => n2266, A2 => pc_lut_20_29_port, B1 => n2267
                           , B2 => pc_lut_21_29_port, ZN => n2877);
   U4439 : NOR4_X1 port map( A1 => n2878, A2 => n2879, A3 => n2880, A4 => n2881
                           , ZN => n2868);
   U4440 : OAI221_X1 port map( B1 => n1976, B2 => n2272, C1 => n1942, C2 => 
                           n2273, A => n2882, ZN => n2881);
   U4441 : AOI22_X1 port map( A1 => n2275, A2 => pc_lut_10_29_port, B1 => n2276
                           , B2 => pc_lut_11_29_port, ZN => n2882);
   U4444 : OAI221_X1 port map( B1 => n1841, B2 => n2277, C1 => n1807, C2 => 
                           n2278, A => n2883, ZN => n2880);
   U4445 : AOI22_X1 port map( A1 => n2280, A2 => pc_lut_14_29_port, B1 => n2281
                           , B2 => pc_lut_15_29_port, ZN => n2883);
   U4448 : OAI221_X1 port map( B1 => n2240, B2 => n2282, C1 => n2206, C2 => 
                           n2283, A => n2884, ZN => n2879);
   U4449 : AOI22_X1 port map( A1 => n2285, A2 => pc_lut_2_29_port, B1 => n2286,
                           B2 => pc_lut_3_29_port, ZN => n2884);
   U4452 : OAI221_X1 port map( B1 => n2108, B2 => n2287, C1 => n2074, C2 => 
                           n2288, A => n2885, ZN => n2878);
   U4453 : AOI22_X1 port map( A1 => n2290, A2 => pc_lut_6_29_port, B1 => n2291,
                           B2 => pc_lut_7_29_port, ZN => n2885);
   U4456 : NAND2_X1 port map( A1 => n2886, A2 => n2887, ZN => N189);
   U4457 : NOR4_X1 port map( A1 => n2888, A2 => n2889, A3 => n2890, A4 => n2891
                           , ZN => n2887);
   U4458 : OAI221_X1 port map( B1 => n1411, B2 => n2248, C1 => n1377, C2 => 
                           n2249, A => n2892, ZN => n2891);
   U4459 : AOI22_X1 port map( A1 => n2251, A2 => pc_lut_26_30_port, B1 => n2252
                           , B2 => pc_lut_27_30_port, ZN => n2892);
   U4462 : OAI221_X1 port map( B1 => n1276, B2 => n2253, C1 => n1241, C2 => 
                           n2254, A => n2893, ZN => n2890);
   U4463 : AOI22_X1 port map( A1 => n2256, A2 => pc_lut_30_30_port, B1 => n2257
                           , B2 => pc_lut_31_30_port, ZN => n2893);
   U4466 : OAI221_X1 port map( B1 => n1675, B2 => n2258, C1 => n1641, C2 => 
                           n2259, A => n2894, ZN => n2889);
   U4467 : AOI22_X1 port map( A1 => n2261, A2 => pc_lut_18_30_port, B1 => n2262
                           , B2 => pc_lut_19_30_port, ZN => n2894);
   U4470 : OAI221_X1 port map( B1 => n1480, B2 => n2263, C1 => n1445, C2 => 
                           n2264, A => n2895, ZN => n2888);
   U4471 : AOI22_X1 port map( A1 => n2266, A2 => pc_lut_20_30_port, B1 => n2267
                           , B2 => pc_lut_21_30_port, ZN => n2895);
   U4474 : NOR4_X1 port map( A1 => n2896, A2 => n2897, A3 => n2898, A4 => n2899
                           , ZN => n2886);
   U4475 : OAI221_X1 port map( B1 => n1945, B2 => n2272, C1 => n1911, C2 => 
                           n2273, A => n2900, ZN => n2899);
   U4476 : AOI22_X1 port map( A1 => n2275, A2 => pc_lut_10_30_port, B1 => n2276
                           , B2 => pc_lut_11_30_port, ZN => n2900);
   U4479 : OAI221_X1 port map( B1 => n1810, B2 => n2277, C1 => n1776, C2 => 
                           n2278, A => n2901, ZN => n2898);
   U4480 : AOI22_X1 port map( A1 => n2280, A2 => pc_lut_14_30_port, B1 => n2281
                           , B2 => pc_lut_15_30_port, ZN => n2901);
   U4483 : OAI221_X1 port map( B1 => n2209, B2 => n2282, C1 => n2175, C2 => 
                           n2283, A => n2902, ZN => n2897);
   U4484 : AOI22_X1 port map( A1 => n2285, A2 => pc_lut_2_30_port, B1 => n2286,
                           B2 => pc_lut_3_30_port, ZN => n2902);
   U4487 : OAI221_X1 port map( B1 => n2077, B2 => n2287, C1 => n2043, C2 => 
                           n2288, A => n2903, ZN => n2896);
   U4488 : AOI22_X1 port map( A1 => n2290, A2 => pc_lut_6_30_port, B1 => n2291,
                           B2 => pc_lut_7_30_port, ZN => n2903);
   U4491 : NAND2_X1 port map( A1 => n2904, A2 => n2905, ZN => N188);
   U4492 : NOR4_X1 port map( A1 => n2906, A2 => n2907, A3 => n2908, A4 => n2909
                           , ZN => n2905);
   U4493 : OAI221_X1 port map( B1 => n1443, B2 => n2248, C1 => n1409, C2 => 
                           n2249, A => n2910, ZN => n2909);
   U4494 : AOI22_X1 port map( A1 => n2251, A2 => pc_lut_26_31_port, B1 => n2252
                           , B2 => pc_lut_27_31_port, ZN => n2910);
   U4497 : OAI221_X1 port map( B1 => n1308, B2 => n2253, C1 => n1274, C2 => 
                           n2254, A => n2911, ZN => n2908);
   U4498 : AOI22_X1 port map( A1 => n2256, A2 => pc_lut_30_31_port, B1 => n2257
                           , B2 => pc_lut_31_31_port, ZN => n2911);
   U4501 : OAI221_X1 port map( B1 => n1707, B2 => n2258, C1 => n1673, C2 => 
                           n2259, A => n2912, ZN => n2907);
   U4502 : AOI22_X1 port map( A1 => n2261, A2 => pc_lut_18_31_port, B1 => n2262
                           , B2 => pc_lut_19_31_port, ZN => n2912);
   U4505 : OAI221_X1 port map( B1 => n1512, B2 => n2263, C1 => n1477, C2 => 
                           n2264, A => n2913, ZN => n2906);
   U4506 : AOI22_X1 port map( A1 => n2266, A2 => pc_lut_20_31_port, B1 => n2267
                           , B2 => pc_lut_21_31_port, ZN => n2913);
   U4509 : NOR4_X1 port map( A1 => n2914, A2 => n2915, A3 => n2916, A4 => n2917
                           , ZN => n2904);
   U4510 : OAI221_X1 port map( B1 => n1977, B2 => n2272, C1 => n1943, C2 => 
                           n2273, A => n2918, ZN => n2917);
   U4511 : AOI22_X1 port map( A1 => n2275, A2 => pc_lut_10_31_port, B1 => n2276
                           , B2 => pc_lut_11_31_port, ZN => n2918);
   U4514 : OAI221_X1 port map( B1 => n1842, B2 => n2277, C1 => n1808, C2 => 
                           n2278, A => n2919, ZN => n2916);
   U4515 : AOI22_X1 port map( A1 => n2280, A2 => pc_lut_14_31_port, B1 => n2281
                           , B2 => pc_lut_15_31_port, ZN => n2919);
   U4518 : OAI221_X1 port map( B1 => n2241, B2 => n2282, C1 => n2207, C2 => 
                           n2283, A => n2920, ZN => n2915);
   U4519 : AOI22_X1 port map( A1 => n2285, A2 => pc_lut_2_31_port, B1 => n2286,
                           B2 => pc_lut_3_31_port, ZN => n2920);
   U4522 : OAI221_X1 port map( B1 => n2109, B2 => n2287, C1 => n2075, C2 => 
                           n2288, A => n2921, ZN => n2914);
   U4523 : AOI22_X1 port map( A1 => n2290, A2 => pc_lut_6_31_port, B1 => n2291,
                           B2 => pc_lut_7_31_port, ZN => n2921);
   U4526 : NAND2_X1 port map( A1 => n2922, A2 => n2923, ZN => N127);
   U4527 : NOR4_X1 port map( A1 => n2924, A2 => n2925, A3 => n2926, A4 => n2927
                           , ZN => n2923);
   U4528 : OAI221_X1 port map( B1 => n299, B2 => n2248, C1 => n265, C2 => n2249
                           , A => n2928, ZN => n2927);
   U4529 : AOI22_X1 port map( A1 => n2251, A2 => pc_target_26_0_port, B1 => 
                           n2252, B2 => pc_target_27_0_port, ZN => n2928);
   U4532 : OAI221_X1 port map( B1 => n159, B2 => n2253, C1 => n108_port, C2 => 
                           n2254, A => n2929, ZN => n2926);
   U4533 : AOI22_X1 port map( A1 => n2256, A2 => pc_target_30_0_port, B1 => 
                           n2257, B2 => pc_target_31_0_port, ZN => n2929);
   U4536 : OAI221_X1 port map( B1 => n575, B2 => n2258, C1 => n541, C2 => n2259
                           , A => n2930, ZN => n2925);
   U4537 : AOI22_X1 port map( A1 => n2261, A2 => pc_target_18_0_port, B1 => 
                           n2262, B2 => pc_target_19_0_port, ZN => n2930);
   U4540 : OAI221_X1 port map( B1 => n369, B2 => n2263, C1 => n334, C2 => n2264
                           , A => n2931, ZN => n2924);
   U4541 : AOI22_X1 port map( A1 => n2266, A2 => pc_target_20_0_port, B1 => 
                           n2267, B2 => pc_target_21_0_port, ZN => n2931);
   U4544 : NOR4_X1 port map( A1 => n2932, A2 => n2933, A3 => n2934, A4 => n2935
                           , ZN => n2922);
   U4545 : OAI221_X1 port map( B1 => n852, B2 => n2272, C1 => n818, C2 => n2273
                           , A => n2936, ZN => n2935);
   U4546 : AOI22_X1 port map( A1 => n2275, A2 => pc_target_10_0_port, B1 => 
                           n2276, B2 => pc_target_11_0_port, ZN => n2936);
   U4549 : OAI221_X1 port map( B1 => n714, B2 => n2277, C1 => n680, C2 => n2278
                           , A => n2937, ZN => n2934);
   U4550 : AOI22_X1 port map( A1 => n2280, A2 => pc_target_14_0_port, B1 => 
                           n2281, B2 => pc_target_15_0_port, ZN => n2937);
   U4553 : OAI221_X1 port map( B1 => n1126, B2 => n2282, C1 => n1092, C2 => 
                           n2283, A => n2938, ZN => n2933);
   U4554 : AOI22_X1 port map( A1 => n2285, A2 => pc_target_2_0_port, B1 => 
                           n2286, B2 => pc_target_3_0_port, ZN => n2938);
   U4557 : OAI221_X1 port map( B1 => n989, B2 => n2287, C1 => n955, C2 => n2288
                           , A => n2939, ZN => n2932);
   U4558 : AOI22_X1 port map( A1 => n2290, A2 => pc_target_6_0_port, B1 => 
                           n2291, B2 => pc_target_7_0_port, ZN => n2939);
   U4561 : NAND2_X1 port map( A1 => n2940, A2 => n2941, ZN => N126);
   U4562 : NOR4_X1 port map( A1 => n2942, A2 => n2943, A3 => n2944, A4 => n2945
                           , ZN => n2941);
   U4563 : OAI221_X1 port map( B1 => n300, B2 => n2248, C1 => n266, C2 => n2249
                           , A => n2946, ZN => n2945);
   U4564 : AOI22_X1 port map( A1 => n2251, A2 => pc_target_26_1_port, B1 => 
                           n2252, B2 => pc_target_27_1_port, ZN => n2946);
   U4567 : OAI221_X1 port map( B1 => n160, B2 => n2253, C1 => n110_port, C2 => 
                           n2254, A => n2947, ZN => n2944);
   U4568 : AOI22_X1 port map( A1 => n2256, A2 => pc_target_30_1_port, B1 => 
                           n2257, B2 => pc_target_31_1_port, ZN => n2947);
   U4571 : OAI221_X1 port map( B1 => n576, B2 => n2258, C1 => n542, C2 => n2259
                           , A => n2948, ZN => n2943);
   U4572 : AOI22_X1 port map( A1 => n2261, A2 => pc_target_18_1_port, B1 => 
                           n2262, B2 => pc_target_19_1_port, ZN => n2948);
   U4575 : OAI221_X1 port map( B1 => n370, B2 => n2263, C1 => n335, C2 => n2264
                           , A => n2949, ZN => n2942);
   U4576 : AOI22_X1 port map( A1 => n2266, A2 => pc_target_20_1_port, B1 => 
                           n2267, B2 => pc_target_21_1_port, ZN => n2949);
   U4579 : NOR4_X1 port map( A1 => n2950, A2 => n2951, A3 => n2952, A4 => n2953
                           , ZN => n2940);
   U4580 : OAI221_X1 port map( B1 => n853, B2 => n2272, C1 => n819, C2 => n2273
                           , A => n2954, ZN => n2953);
   U4581 : AOI22_X1 port map( A1 => n2275, A2 => pc_target_10_1_port, B1 => 
                           n2276, B2 => pc_target_11_1_port, ZN => n2954);
   U4584 : OAI221_X1 port map( B1 => n715, B2 => n2277, C1 => n681, C2 => n2278
                           , A => n2955, ZN => n2952);
   U4585 : AOI22_X1 port map( A1 => n2280, A2 => pc_target_14_1_port, B1 => 
                           n2281, B2 => pc_target_15_1_port, ZN => n2955);
   U4588 : OAI221_X1 port map( B1 => n1127, B2 => n2282, C1 => n1093, C2 => 
                           n2283, A => n2956, ZN => n2951);
   U4589 : AOI22_X1 port map( A1 => n2285, A2 => pc_target_2_1_port, B1 => 
                           n2286, B2 => pc_target_3_1_port, ZN => n2956);
   U4592 : OAI221_X1 port map( B1 => n990, B2 => n2287, C1 => n956, C2 => n2288
                           , A => n2957, ZN => n2950);
   U4593 : AOI22_X1 port map( A1 => n2290, A2 => pc_target_6_1_port, B1 => 
                           n2291, B2 => pc_target_7_1_port, ZN => n2957);
   U4596 : NAND2_X1 port map( A1 => n2958, A2 => n2959, ZN => N125);
   U4597 : NOR4_X1 port map( A1 => n2960, A2 => n2961, A3 => n2962, A4 => n2963
                           , ZN => n2959);
   U4598 : OAI221_X1 port map( B1 => n298, B2 => n2248, C1 => n264, C2 => n2249
                           , A => n2964, ZN => n2963);
   U4599 : AOI22_X1 port map( A1 => n2251, A2 => pc_target_26_2_port, B1 => 
                           n2252, B2 => pc_target_27_2_port, ZN => n2964);
   U4602 : OAI221_X1 port map( B1 => n158, B2 => n2253, C1 => n106_port, C2 => 
                           n2254, A => n2965, ZN => n2962);
   U4603 : AOI22_X1 port map( A1 => n2256, A2 => pc_target_30_2_port, B1 => 
                           n2257, B2 => pc_target_31_2_port, ZN => n2965);
   U4606 : OAI221_X1 port map( B1 => n574, B2 => n2258, C1 => n540, C2 => n2259
                           , A => n2966, ZN => n2961);
   U4607 : AOI22_X1 port map( A1 => n2261, A2 => pc_target_18_2_port, B1 => 
                           n2262, B2 => pc_target_19_2_port, ZN => n2966);
   U4610 : OAI221_X1 port map( B1 => n368, B2 => n2263, C1 => n333, C2 => n2264
                           , A => n2967, ZN => n2960);
   U4611 : AOI22_X1 port map( A1 => n2266, A2 => pc_target_20_2_port, B1 => 
                           n2267, B2 => pc_target_21_2_port, ZN => n2967);
   U4614 : NOR4_X1 port map( A1 => n2968, A2 => n2969, A3 => n2970, A4 => n2971
                           , ZN => n2958);
   U4615 : OAI221_X1 port map( B1 => n851, B2 => n2272, C1 => n817, C2 => n2273
                           , A => n2972, ZN => n2971);
   U4616 : AOI22_X1 port map( A1 => n2275, A2 => pc_target_10_2_port, B1 => 
                           n2276, B2 => pc_target_11_2_port, ZN => n2972);
   U4619 : OAI221_X1 port map( B1 => n713, B2 => n2277, C1 => n679, C2 => n2278
                           , A => n2973, ZN => n2970);
   U4620 : AOI22_X1 port map( A1 => n2280, A2 => pc_target_14_2_port, B1 => 
                           n2281, B2 => pc_target_15_2_port, ZN => n2973);
   U4623 : OAI221_X1 port map( B1 => n1125, B2 => n2282, C1 => n1091, C2 => 
                           n2283, A => n2974, ZN => n2969);
   U4624 : AOI22_X1 port map( A1 => n2285, A2 => pc_target_2_2_port, B1 => 
                           n2286, B2 => pc_target_3_2_port, ZN => n2974);
   U4627 : OAI221_X1 port map( B1 => n988, B2 => n2287, C1 => n954, C2 => n2288
                           , A => n2975, ZN => n2968);
   U4628 : AOI22_X1 port map( A1 => n2290, A2 => pc_target_6_2_port, B1 => 
                           n2291, B2 => pc_target_7_2_port, ZN => n2975);
   U4631 : NAND2_X1 port map( A1 => n2976, A2 => n2977, ZN => N124);
   U4632 : NOR4_X1 port map( A1 => n2978, A2 => n2979, A3 => n2980, A4 => n2981
                           , ZN => n2977);
   U4633 : OAI221_X1 port map( B1 => n301, B2 => n2248, C1 => n267, C2 => n2249
                           , A => n2982, ZN => n2981);
   U4634 : AOI22_X1 port map( A1 => n2251, A2 => pc_target_26_3_port, B1 => 
                           n2252, B2 => pc_target_27_3_port, ZN => n2982);
   U4637 : OAI221_X1 port map( B1 => n161, B2 => n2253, C1 => n112_port, C2 => 
                           n2254, A => n2983, ZN => n2980);
   U4638 : AOI22_X1 port map( A1 => n2256, A2 => pc_target_30_3_port, B1 => 
                           n2257, B2 => pc_target_31_3_port, ZN => n2983);
   U4641 : OAI221_X1 port map( B1 => n577, B2 => n2258, C1 => n543, C2 => n2259
                           , A => n2984, ZN => n2979);
   U4642 : AOI22_X1 port map( A1 => n2261, A2 => pc_target_18_3_port, B1 => 
                           n2262, B2 => pc_target_19_3_port, ZN => n2984);
   U4645 : OAI221_X1 port map( B1 => n371, B2 => n2263, C1 => n336, C2 => n2264
                           , A => n2985, ZN => n2978);
   U4646 : AOI22_X1 port map( A1 => n2266, A2 => pc_target_20_3_port, B1 => 
                           n2267, B2 => pc_target_21_3_port, ZN => n2985);
   U4649 : NOR4_X1 port map( A1 => n2986, A2 => n2987, A3 => n2988, A4 => n2989
                           , ZN => n2976);
   U4650 : OAI221_X1 port map( B1 => n854, B2 => n2272, C1 => n820, C2 => n2273
                           , A => n2990, ZN => n2989);
   U4651 : AOI22_X1 port map( A1 => n2275, A2 => pc_target_10_3_port, B1 => 
                           n2276, B2 => pc_target_11_3_port, ZN => n2990);
   U4654 : OAI221_X1 port map( B1 => n716, B2 => n2277, C1 => n682, C2 => n2278
                           , A => n2991, ZN => n2988);
   U4655 : AOI22_X1 port map( A1 => n2280, A2 => pc_target_14_3_port, B1 => 
                           n2281, B2 => pc_target_15_3_port, ZN => n2991);
   U4658 : OAI221_X1 port map( B1 => n1128, B2 => n2282, C1 => n1094, C2 => 
                           n2283, A => n2992, ZN => n2987);
   U4659 : AOI22_X1 port map( A1 => n2285, A2 => pc_target_2_3_port, B1 => 
                           n2286, B2 => pc_target_3_3_port, ZN => n2992);
   U4662 : OAI221_X1 port map( B1 => n991, B2 => n2287, C1 => n957, C2 => n2288
                           , A => n2993, ZN => n2986);
   U4663 : AOI22_X1 port map( A1 => n2290, A2 => pc_target_6_3_port, B1 => 
                           n2291, B2 => pc_target_7_3_port, ZN => n2993);
   U4666 : NAND2_X1 port map( A1 => n2994, A2 => n2995, ZN => N123);
   U4667 : NOR4_X1 port map( A1 => n2996, A2 => n2997, A3 => n2998, A4 => n2999
                           , ZN => n2995);
   U4668 : OAI221_X1 port map( B1 => n297, B2 => n2248, C1 => n263, C2 => n2249
                           , A => n3000, ZN => n2999);
   U4669 : AOI22_X1 port map( A1 => n2251, A2 => pc_target_26_4_port, B1 => 
                           n2252, B2 => pc_target_27_4_port, ZN => n3000);
   U4672 : OAI221_X1 port map( B1 => n157, B2 => n2253, C1 => n104_port, C2 => 
                           n2254, A => n3001, ZN => n2998);
   U4673 : AOI22_X1 port map( A1 => n2256, A2 => pc_target_30_4_port, B1 => 
                           n2257, B2 => pc_target_31_4_port, ZN => n3001);
   U4676 : OAI221_X1 port map( B1 => n573, B2 => n2258, C1 => n539, C2 => n2259
                           , A => n3002, ZN => n2997);
   U4677 : AOI22_X1 port map( A1 => n2261, A2 => pc_target_18_4_port, B1 => 
                           n2262, B2 => pc_target_19_4_port, ZN => n3002);
   U4680 : OAI221_X1 port map( B1 => n367, B2 => n2263, C1 => n332, C2 => n2264
                           , A => n3003, ZN => n2996);
   U4681 : AOI22_X1 port map( A1 => n2266, A2 => pc_target_20_4_port, B1 => 
                           n2267, B2 => pc_target_21_4_port, ZN => n3003);
   U4684 : NOR4_X1 port map( A1 => n3004, A2 => n3005, A3 => n3006, A4 => n3007
                           , ZN => n2994);
   U4685 : OAI221_X1 port map( B1 => n850, B2 => n2272, C1 => n816, C2 => n2273
                           , A => n3008, ZN => n3007);
   U4686 : AOI22_X1 port map( A1 => n2275, A2 => pc_target_10_4_port, B1 => 
                           n2276, B2 => pc_target_11_4_port, ZN => n3008);
   U4689 : OAI221_X1 port map( B1 => n712, B2 => n2277, C1 => n678, C2 => n2278
                           , A => n3009, ZN => n3006);
   U4690 : AOI22_X1 port map( A1 => n2280, A2 => pc_target_14_4_port, B1 => 
                           n2281, B2 => pc_target_15_4_port, ZN => n3009);
   U4693 : OAI221_X1 port map( B1 => n1124, B2 => n2282, C1 => n1090, C2 => 
                           n2283, A => n3010, ZN => n3005);
   U4694 : AOI22_X1 port map( A1 => n2285, A2 => pc_target_2_4_port, B1 => 
                           n2286, B2 => pc_target_3_4_port, ZN => n3010);
   U4697 : OAI221_X1 port map( B1 => n987, B2 => n2287, C1 => n953, C2 => n2288
                           , A => n3011, ZN => n3004);
   U4698 : AOI22_X1 port map( A1 => n2290, A2 => pc_target_6_4_port, B1 => 
                           n2291, B2 => pc_target_7_4_port, ZN => n3011);
   U4701 : NAND2_X1 port map( A1 => n3012, A2 => n3013, ZN => N122);
   U4702 : NOR4_X1 port map( A1 => n3014, A2 => n3015, A3 => n3016, A4 => n3017
                           , ZN => n3013);
   U4703 : OAI221_X1 port map( B1 => n302, B2 => n2248, C1 => n268, C2 => n2249
                           , A => n3018, ZN => n3017);
   U4704 : AOI22_X1 port map( A1 => n2251, A2 => pc_target_26_5_port, B1 => 
                           n2252, B2 => pc_target_27_5_port, ZN => n3018);
   U4707 : OAI221_X1 port map( B1 => n162, B2 => n2253, C1 => n114_port, C2 => 
                           n2254, A => n3019, ZN => n3016);
   U4708 : AOI22_X1 port map( A1 => n2256, A2 => pc_target_30_5_port, B1 => 
                           n2257, B2 => pc_target_31_5_port, ZN => n3019);
   U4711 : OAI221_X1 port map( B1 => n578, B2 => n2258, C1 => n544, C2 => n2259
                           , A => n3020, ZN => n3015);
   U4712 : AOI22_X1 port map( A1 => n2261, A2 => pc_target_18_5_port, B1 => 
                           n2262, B2 => pc_target_19_5_port, ZN => n3020);
   U4715 : OAI221_X1 port map( B1 => n372, B2 => n2263, C1 => n337, C2 => n2264
                           , A => n3021, ZN => n3014);
   U4716 : AOI22_X1 port map( A1 => n2266, A2 => pc_target_20_5_port, B1 => 
                           n2267, B2 => pc_target_21_5_port, ZN => n3021);
   U4719 : NOR4_X1 port map( A1 => n3022, A2 => n3023, A3 => n3024, A4 => n3025
                           , ZN => n3012);
   U4720 : OAI221_X1 port map( B1 => n855, B2 => n2272, C1 => n821, C2 => n2273
                           , A => n3026, ZN => n3025);
   U4721 : AOI22_X1 port map( A1 => n2275, A2 => pc_target_10_5_port, B1 => 
                           n2276, B2 => pc_target_11_5_port, ZN => n3026);
   U4724 : OAI221_X1 port map( B1 => n717, B2 => n2277, C1 => n683, C2 => n2278
                           , A => n3027, ZN => n3024);
   U4725 : AOI22_X1 port map( A1 => n2280, A2 => pc_target_14_5_port, B1 => 
                           n2281, B2 => pc_target_15_5_port, ZN => n3027);
   U4728 : OAI221_X1 port map( B1 => n1129, B2 => n2282, C1 => n1095, C2 => 
                           n2283, A => n3028, ZN => n3023);
   U4729 : AOI22_X1 port map( A1 => n2285, A2 => pc_target_2_5_port, B1 => 
                           n2286, B2 => pc_target_3_5_port, ZN => n3028);
   U4732 : OAI221_X1 port map( B1 => n992, B2 => n2287, C1 => n958, C2 => n2288
                           , A => n3029, ZN => n3022);
   U4733 : AOI22_X1 port map( A1 => n2290, A2 => pc_target_6_5_port, B1 => 
                           n2291, B2 => pc_target_7_5_port, ZN => n3029);
   U4736 : NAND2_X1 port map( A1 => n3030, A2 => n3031, ZN => N121);
   U4737 : NOR4_X1 port map( A1 => n3032, A2 => n3033, A3 => n3034, A4 => n3035
                           , ZN => n3031);
   U4738 : OAI221_X1 port map( B1 => n296, B2 => n2248, C1 => n262, C2 => n2249
                           , A => n3036, ZN => n3035);
   U4739 : AOI22_X1 port map( A1 => n2251, A2 => pc_target_26_6_port, B1 => 
                           n2252, B2 => pc_target_27_6_port, ZN => n3036);
   U4742 : OAI221_X1 port map( B1 => n156, B2 => n2253, C1 => n102_port, C2 => 
                           n2254, A => n3037, ZN => n3034);
   U4743 : AOI22_X1 port map( A1 => n2256, A2 => pc_target_30_6_port, B1 => 
                           n2257, B2 => pc_target_31_6_port, ZN => n3037);
   U4746 : OAI221_X1 port map( B1 => n572, B2 => n2258, C1 => n538, C2 => n2259
                           , A => n3038, ZN => n3033);
   U4747 : AOI22_X1 port map( A1 => n2261, A2 => pc_target_18_6_port, B1 => 
                           n2262, B2 => pc_target_19_6_port, ZN => n3038);
   U4750 : OAI221_X1 port map( B1 => n366, B2 => n2263, C1 => n331, C2 => n2264
                           , A => n3039, ZN => n3032);
   U4751 : AOI22_X1 port map( A1 => n2266, A2 => pc_target_20_6_port, B1 => 
                           n2267, B2 => pc_target_21_6_port, ZN => n3039);
   U4754 : NOR4_X1 port map( A1 => n3040, A2 => n3041, A3 => n3042, A4 => n3043
                           , ZN => n3030);
   U4755 : OAI221_X1 port map( B1 => n849, B2 => n2272, C1 => n815, C2 => n2273
                           , A => n3044, ZN => n3043);
   U4756 : AOI22_X1 port map( A1 => n2275, A2 => pc_target_10_6_port, B1 => 
                           n2276, B2 => pc_target_11_6_port, ZN => n3044);
   U4759 : OAI221_X1 port map( B1 => n711, B2 => n2277, C1 => n677, C2 => n2278
                           , A => n3045, ZN => n3042);
   U4760 : AOI22_X1 port map( A1 => n2280, A2 => pc_target_14_6_port, B1 => 
                           n2281, B2 => pc_target_15_6_port, ZN => n3045);
   U4763 : OAI221_X1 port map( B1 => n1123, B2 => n2282, C1 => n1089, C2 => 
                           n2283, A => n3046, ZN => n3041);
   U4764 : AOI22_X1 port map( A1 => n2285, A2 => pc_target_2_6_port, B1 => 
                           n2286, B2 => pc_target_3_6_port, ZN => n3046);
   U4767 : OAI221_X1 port map( B1 => n986, B2 => n2287, C1 => n952, C2 => n2288
                           , A => n3047, ZN => n3040);
   U4768 : AOI22_X1 port map( A1 => n2290, A2 => pc_target_6_6_port, B1 => 
                           n2291, B2 => pc_target_7_6_port, ZN => n3047);
   U4771 : NAND2_X1 port map( A1 => n3048, A2 => n3049, ZN => N120);
   U4772 : NOR4_X1 port map( A1 => n3050, A2 => n3051, A3 => n3052, A4 => n3053
                           , ZN => n3049);
   U4773 : OAI221_X1 port map( B1 => n303, B2 => n2248, C1 => n269, C2 => n2249
                           , A => n3054, ZN => n3053);
   U4774 : AOI22_X1 port map( A1 => n2251, A2 => pc_target_26_7_port, B1 => 
                           n2252, B2 => pc_target_27_7_port, ZN => n3054);
   U4777 : OAI221_X1 port map( B1 => n163, B2 => n2253, C1 => n116_port, C2 => 
                           n2254, A => n3055, ZN => n3052);
   U4778 : AOI22_X1 port map( A1 => n2256, A2 => pc_target_30_7_port, B1 => 
                           n2257, B2 => pc_target_31_7_port, ZN => n3055);
   U4781 : OAI221_X1 port map( B1 => n579, B2 => n2258, C1 => n545, C2 => n2259
                           , A => n3056, ZN => n3051);
   U4782 : AOI22_X1 port map( A1 => n2261, A2 => pc_target_18_7_port, B1 => 
                           n2262, B2 => pc_target_19_7_port, ZN => n3056);
   U4785 : OAI221_X1 port map( B1 => n373, B2 => n2263, C1 => n338, C2 => n2264
                           , A => n3057, ZN => n3050);
   U4786 : AOI22_X1 port map( A1 => n2266, A2 => pc_target_20_7_port, B1 => 
                           n2267, B2 => pc_target_21_7_port, ZN => n3057);
   U4789 : NOR4_X1 port map( A1 => n3058, A2 => n3059, A3 => n3060, A4 => n3061
                           , ZN => n3048);
   U4790 : OAI221_X1 port map( B1 => n856, B2 => n2272, C1 => n822, C2 => n2273
                           , A => n3062, ZN => n3061);
   U4791 : AOI22_X1 port map( A1 => n2275, A2 => pc_target_10_7_port, B1 => 
                           n2276, B2 => pc_target_11_7_port, ZN => n3062);
   U4794 : OAI221_X1 port map( B1 => n718, B2 => n2277, C1 => n684, C2 => n2278
                           , A => n3063, ZN => n3060);
   U4795 : AOI22_X1 port map( A1 => n2280, A2 => pc_target_14_7_port, B1 => 
                           n2281, B2 => pc_target_15_7_port, ZN => n3063);
   U4798 : OAI221_X1 port map( B1 => n1130, B2 => n2282, C1 => n1096, C2 => 
                           n2283, A => n3064, ZN => n3059);
   U4799 : AOI22_X1 port map( A1 => n2285, A2 => pc_target_2_7_port, B1 => 
                           n2286, B2 => pc_target_3_7_port, ZN => n3064);
   U4802 : OAI221_X1 port map( B1 => n993, B2 => n2287, C1 => n959, C2 => n2288
                           , A => n3065, ZN => n3058);
   U4803 : AOI22_X1 port map( A1 => n2290, A2 => pc_target_6_7_port, B1 => 
                           n2291, B2 => pc_target_7_7_port, ZN => n3065);
   U4806 : NAND2_X1 port map( A1 => n3066, A2 => n3067, ZN => N119);
   U4807 : NOR4_X1 port map( A1 => n3068, A2 => n3069, A3 => n3070, A4 => n3071
                           , ZN => n3067);
   U4808 : OAI221_X1 port map( B1 => n295, B2 => n2248, C1 => n261, C2 => n2249
                           , A => n3072, ZN => n3071);
   U4809 : AOI22_X1 port map( A1 => n2251, A2 => pc_target_26_8_port, B1 => 
                           n2252, B2 => pc_target_27_8_port, ZN => n3072);
   U4812 : OAI221_X1 port map( B1 => n155, B2 => n2253, C1 => n100_port, C2 => 
                           n2254, A => n3073, ZN => n3070);
   U4813 : AOI22_X1 port map( A1 => n2256, A2 => pc_target_30_8_port, B1 => 
                           n2257, B2 => pc_target_31_8_port, ZN => n3073);
   U4816 : OAI221_X1 port map( B1 => n571, B2 => n2258, C1 => n537, C2 => n2259
                           , A => n3074, ZN => n3069);
   U4817 : AOI22_X1 port map( A1 => n2261, A2 => pc_target_18_8_port, B1 => 
                           n2262, B2 => pc_target_19_8_port, ZN => n3074);
   U4820 : OAI221_X1 port map( B1 => n365, B2 => n2263, C1 => n330, C2 => n2264
                           , A => n3075, ZN => n3068);
   U4821 : AOI22_X1 port map( A1 => n2266, A2 => pc_target_20_8_port, B1 => 
                           n2267, B2 => pc_target_21_8_port, ZN => n3075);
   U4824 : NOR4_X1 port map( A1 => n3076, A2 => n3077, A3 => n3078, A4 => n3079
                           , ZN => n3066);
   U4825 : OAI221_X1 port map( B1 => n848, B2 => n2272, C1 => n814, C2 => n2273
                           , A => n3080, ZN => n3079);
   U4826 : AOI22_X1 port map( A1 => n2275, A2 => pc_target_10_8_port, B1 => 
                           n2276, B2 => pc_target_11_8_port, ZN => n3080);
   U4829 : OAI221_X1 port map( B1 => n710, B2 => n2277, C1 => n676, C2 => n2278
                           , A => n3081, ZN => n3078);
   U4830 : AOI22_X1 port map( A1 => n2280, A2 => pc_target_14_8_port, B1 => 
                           n2281, B2 => pc_target_15_8_port, ZN => n3081);
   U4833 : OAI221_X1 port map( B1 => n1122, B2 => n2282, C1 => n1088, C2 => 
                           n2283, A => n3082, ZN => n3077);
   U4834 : AOI22_X1 port map( A1 => n2285, A2 => pc_target_2_8_port, B1 => 
                           n2286, B2 => pc_target_3_8_port, ZN => n3082);
   U4837 : OAI221_X1 port map( B1 => n985, B2 => n2287, C1 => n951, C2 => n2288
                           , A => n3083, ZN => n3076);
   U4838 : AOI22_X1 port map( A1 => n2290, A2 => pc_target_6_8_port, B1 => 
                           n2291, B2 => pc_target_7_8_port, ZN => n3083);
   U4841 : NAND2_X1 port map( A1 => n3084, A2 => n3085, ZN => N118);
   U4842 : NOR4_X1 port map( A1 => n3086, A2 => n3087, A3 => n3088, A4 => n3089
                           , ZN => n3085);
   U4843 : OAI221_X1 port map( B1 => n304, B2 => n2248, C1 => n270, C2 => n2249
                           , A => n3090, ZN => n3089);
   U4844 : AOI22_X1 port map( A1 => n2251, A2 => pc_target_26_9_port, B1 => 
                           n2252, B2 => pc_target_27_9_port, ZN => n3090);
   U4847 : OAI221_X1 port map( B1 => n164, B2 => n2253, C1 => n118_port, C2 => 
                           n2254, A => n3091, ZN => n3088);
   U4848 : AOI22_X1 port map( A1 => n2256, A2 => pc_target_30_9_port, B1 => 
                           n2257, B2 => pc_target_31_9_port, ZN => n3091);
   U4851 : OAI221_X1 port map( B1 => n580, B2 => n2258, C1 => n546, C2 => n2259
                           , A => n3092, ZN => n3087);
   U4852 : AOI22_X1 port map( A1 => n2261, A2 => pc_target_18_9_port, B1 => 
                           n2262, B2 => pc_target_19_9_port, ZN => n3092);
   U4855 : OAI221_X1 port map( B1 => n374, B2 => n2263, C1 => n339, C2 => n2264
                           , A => n3093, ZN => n3086);
   U4856 : AOI22_X1 port map( A1 => n2266, A2 => pc_target_20_9_port, B1 => 
                           n2267, B2 => pc_target_21_9_port, ZN => n3093);
   U4859 : NOR4_X1 port map( A1 => n3094, A2 => n3095, A3 => n3096, A4 => n3097
                           , ZN => n3084);
   U4860 : OAI221_X1 port map( B1 => n857, B2 => n2272, C1 => n823, C2 => n2273
                           , A => n3098, ZN => n3097);
   U4861 : AOI22_X1 port map( A1 => n2275, A2 => pc_target_10_9_port, B1 => 
                           n2276, B2 => pc_target_11_9_port, ZN => n3098);
   U4864 : OAI221_X1 port map( B1 => n719, B2 => n2277, C1 => n685, C2 => n2278
                           , A => n3099, ZN => n3096);
   U4865 : AOI22_X1 port map( A1 => n2280, A2 => pc_target_14_9_port, B1 => 
                           n2281, B2 => pc_target_15_9_port, ZN => n3099);
   U4868 : OAI221_X1 port map( B1 => n1131, B2 => n2282, C1 => n1097, C2 => 
                           n2283, A => n3100, ZN => n3095);
   U4869 : AOI22_X1 port map( A1 => n2285, A2 => pc_target_2_9_port, B1 => 
                           n2286, B2 => pc_target_3_9_port, ZN => n3100);
   U4872 : OAI221_X1 port map( B1 => n994, B2 => n2287, C1 => n960, C2 => n2288
                           , A => n3101, ZN => n3094);
   U4873 : AOI22_X1 port map( A1 => n2290, A2 => pc_target_6_9_port, B1 => 
                           n2291, B2 => pc_target_7_9_port, ZN => n3101);
   U4876 : NAND2_X1 port map( A1 => n3102, A2 => n3103, ZN => N117);
   U4877 : NOR4_X1 port map( A1 => n3104, A2 => n3105, A3 => n3106, A4 => n3107
                           , ZN => n3103);
   U4878 : OAI221_X1 port map( B1 => n294, B2 => n2248, C1 => n260, C2 => n2249
                           , A => n3108, ZN => n3107);
   U4879 : AOI22_X1 port map( A1 => n2251, A2 => pc_target_26_10_port, B1 => 
                           n2252, B2 => pc_target_27_10_port, ZN => n3108);
   U4882 : OAI221_X1 port map( B1 => n154, B2 => n2253, C1 => n98_port, C2 => 
                           n2254, A => n3109, ZN => n3106);
   U4883 : AOI22_X1 port map( A1 => n2256, A2 => pc_target_30_10_port, B1 => 
                           n2257, B2 => pc_target_31_10_port, ZN => n3109);
   U4886 : OAI221_X1 port map( B1 => n570, B2 => n2258, C1 => n536, C2 => n2259
                           , A => n3110, ZN => n3105);
   U4887 : AOI22_X1 port map( A1 => n2261, A2 => pc_target_18_10_port, B1 => 
                           n2262, B2 => pc_target_19_10_port, ZN => n3110);
   U4890 : OAI221_X1 port map( B1 => n364, B2 => n2263, C1 => n329, C2 => n2264
                           , A => n3111, ZN => n3104);
   U4891 : AOI22_X1 port map( A1 => n2266, A2 => pc_target_20_10_port, B1 => 
                           n2267, B2 => pc_target_21_10_port, ZN => n3111);
   U4894 : NOR4_X1 port map( A1 => n3112, A2 => n3113, A3 => n3114, A4 => n3115
                           , ZN => n3102);
   U4895 : OAI221_X1 port map( B1 => n847, B2 => n2272, C1 => n813, C2 => n2273
                           , A => n3116, ZN => n3115);
   U4896 : AOI22_X1 port map( A1 => n2275, A2 => pc_target_10_10_port, B1 => 
                           n2276, B2 => pc_target_11_10_port, ZN => n3116);
   U4899 : OAI221_X1 port map( B1 => n709, B2 => n2277, C1 => n675, C2 => n2278
                           , A => n3117, ZN => n3114);
   U4900 : AOI22_X1 port map( A1 => n2280, A2 => pc_target_14_10_port, B1 => 
                           n2281, B2 => pc_target_15_10_port, ZN => n3117);
   U4903 : OAI221_X1 port map( B1 => n1121, B2 => n2282, C1 => n1087, C2 => 
                           n2283, A => n3118, ZN => n3113);
   U4904 : AOI22_X1 port map( A1 => n2285, A2 => pc_target_2_10_port, B1 => 
                           n2286, B2 => pc_target_3_10_port, ZN => n3118);
   U4907 : OAI221_X1 port map( B1 => n984, B2 => n2287, C1 => n950, C2 => n2288
                           , A => n3119, ZN => n3112);
   U4908 : AOI22_X1 port map( A1 => n2290, A2 => pc_target_6_10_port, B1 => 
                           n2291, B2 => pc_target_7_10_port, ZN => n3119);
   U4911 : NAND2_X1 port map( A1 => n3120, A2 => n3121, ZN => N116);
   U4912 : NOR4_X1 port map( A1 => n3122, A2 => n3123, A3 => n3124, A4 => n3125
                           , ZN => n3121);
   U4913 : OAI221_X1 port map( B1 => n305, B2 => n2248, C1 => n271, C2 => n2249
                           , A => n3126, ZN => n3125);
   U4914 : AOI22_X1 port map( A1 => n2251, A2 => pc_target_26_11_port, B1 => 
                           n2252, B2 => pc_target_27_11_port, ZN => n3126);
   U4917 : OAI221_X1 port map( B1 => n165, B2 => n2253, C1 => n120_port, C2 => 
                           n2254, A => n3127, ZN => n3124);
   U4918 : AOI22_X1 port map( A1 => n2256, A2 => pc_target_30_11_port, B1 => 
                           n2257, B2 => pc_target_31_11_port, ZN => n3127);
   U4921 : OAI221_X1 port map( B1 => n581, B2 => n2258, C1 => n547, C2 => n2259
                           , A => n3128, ZN => n3123);
   U4922 : AOI22_X1 port map( A1 => n2261, A2 => pc_target_18_11_port, B1 => 
                           n2262, B2 => pc_target_19_11_port, ZN => n3128);
   U4925 : OAI221_X1 port map( B1 => n375, B2 => n2263, C1 => n340, C2 => n2264
                           , A => n3129, ZN => n3122);
   U4926 : AOI22_X1 port map( A1 => n2266, A2 => pc_target_20_11_port, B1 => 
                           n2267, B2 => pc_target_21_11_port, ZN => n3129);
   U4929 : NOR4_X1 port map( A1 => n3130, A2 => n3131, A3 => n3132, A4 => n3133
                           , ZN => n3120);
   U4930 : OAI221_X1 port map( B1 => n858, B2 => n2272, C1 => n824, C2 => n2273
                           , A => n3134, ZN => n3133);
   U4931 : AOI22_X1 port map( A1 => n2275, A2 => pc_target_10_11_port, B1 => 
                           n2276, B2 => pc_target_11_11_port, ZN => n3134);
   U4934 : OAI221_X1 port map( B1 => n720, B2 => n2277, C1 => n686, C2 => n2278
                           , A => n3135, ZN => n3132);
   U4935 : AOI22_X1 port map( A1 => n2280, A2 => pc_target_14_11_port, B1 => 
                           n2281, B2 => pc_target_15_11_port, ZN => n3135);
   U4938 : OAI221_X1 port map( B1 => n1132, B2 => n2282, C1 => n1098, C2 => 
                           n2283, A => n3136, ZN => n3131);
   U4939 : AOI22_X1 port map( A1 => n2285, A2 => pc_target_2_11_port, B1 => 
                           n2286, B2 => pc_target_3_11_port, ZN => n3136);
   U4942 : OAI221_X1 port map( B1 => n995, B2 => n2287, C1 => n961, C2 => n2288
                           , A => n3137, ZN => n3130);
   U4943 : AOI22_X1 port map( A1 => n2290, A2 => pc_target_6_11_port, B1 => 
                           n2291, B2 => pc_target_7_11_port, ZN => n3137);
   U4946 : NAND2_X1 port map( A1 => n3138, A2 => n3139, ZN => N115);
   U4947 : NOR4_X1 port map( A1 => n3140, A2 => n3141, A3 => n3142, A4 => n3143
                           , ZN => n3139);
   U4948 : OAI221_X1 port map( B1 => n293, B2 => n2248, C1 => n259, C2 => n2249
                           , A => n3144, ZN => n3143);
   U4949 : AOI22_X1 port map( A1 => n2251, A2 => pc_target_26_12_port, B1 => 
                           n2252, B2 => pc_target_27_12_port, ZN => n3144);
   U4952 : OAI221_X1 port map( B1 => n153, B2 => n2253, C1 => n96_port, C2 => 
                           n2254, A => n3145, ZN => n3142);
   U4953 : AOI22_X1 port map( A1 => n2256, A2 => pc_target_30_12_port, B1 => 
                           n2257, B2 => pc_target_31_12_port, ZN => n3145);
   U4956 : OAI221_X1 port map( B1 => n569, B2 => n2258, C1 => n535, C2 => n2259
                           , A => n3146, ZN => n3141);
   U4957 : AOI22_X1 port map( A1 => n2261, A2 => pc_target_18_12_port, B1 => 
                           n2262, B2 => pc_target_19_12_port, ZN => n3146);
   U4960 : OAI221_X1 port map( B1 => n363, B2 => n2263, C1 => n328, C2 => n2264
                           , A => n3147, ZN => n3140);
   U4961 : AOI22_X1 port map( A1 => n2266, A2 => pc_target_20_12_port, B1 => 
                           n2267, B2 => pc_target_21_12_port, ZN => n3147);
   U4964 : NOR4_X1 port map( A1 => n3148, A2 => n3149, A3 => n3150, A4 => n3151
                           , ZN => n3138);
   U4965 : OAI221_X1 port map( B1 => n846, B2 => n2272, C1 => n812, C2 => n2273
                           , A => n3152, ZN => n3151);
   U4966 : AOI22_X1 port map( A1 => n2275, A2 => pc_target_10_12_port, B1 => 
                           n2276, B2 => pc_target_11_12_port, ZN => n3152);
   U4969 : OAI221_X1 port map( B1 => n708, B2 => n2277, C1 => n674, C2 => n2278
                           , A => n3153, ZN => n3150);
   U4970 : AOI22_X1 port map( A1 => n2280, A2 => pc_target_14_12_port, B1 => 
                           n2281, B2 => pc_target_15_12_port, ZN => n3153);
   U4973 : OAI221_X1 port map( B1 => n1120, B2 => n2282, C1 => n1086, C2 => 
                           n2283, A => n3154, ZN => n3149);
   U4974 : AOI22_X1 port map( A1 => n2285, A2 => pc_target_2_12_port, B1 => 
                           n2286, B2 => pc_target_3_12_port, ZN => n3154);
   U4977 : OAI221_X1 port map( B1 => n983, B2 => n2287, C1 => n949, C2 => n2288
                           , A => n3155, ZN => n3148);
   U4978 : AOI22_X1 port map( A1 => n2290, A2 => pc_target_6_12_port, B1 => 
                           n2291, B2 => pc_target_7_12_port, ZN => n3155);
   U4981 : NAND2_X1 port map( A1 => n3156, A2 => n3157, ZN => N114);
   U4982 : NOR4_X1 port map( A1 => n3158, A2 => n3159, A3 => n3160, A4 => n3161
                           , ZN => n3157);
   U4983 : OAI221_X1 port map( B1 => n306, B2 => n2248, C1 => n272, C2 => n2249
                           , A => n3162, ZN => n3161);
   U4984 : AOI22_X1 port map( A1 => n2251, A2 => pc_target_26_13_port, B1 => 
                           n2252, B2 => pc_target_27_13_port, ZN => n3162);
   U4987 : OAI221_X1 port map( B1 => n166, B2 => n2253, C1 => n122_port, C2 => 
                           n2254, A => n3163, ZN => n3160);
   U4988 : AOI22_X1 port map( A1 => n2256, A2 => pc_target_30_13_port, B1 => 
                           n2257, B2 => pc_target_31_13_port, ZN => n3163);
   U4991 : OAI221_X1 port map( B1 => n582, B2 => n2258, C1 => n548, C2 => n2259
                           , A => n3164, ZN => n3159);
   U4992 : AOI22_X1 port map( A1 => n2261, A2 => pc_target_18_13_port, B1 => 
                           n2262, B2 => pc_target_19_13_port, ZN => n3164);
   U4995 : OAI221_X1 port map( B1 => n376, B2 => n2263, C1 => n341, C2 => n2264
                           , A => n3165, ZN => n3158);
   U4996 : AOI22_X1 port map( A1 => n2266, A2 => pc_target_20_13_port, B1 => 
                           n2267, B2 => pc_target_21_13_port, ZN => n3165);
   U4999 : NOR4_X1 port map( A1 => n3166, A2 => n3167, A3 => n3168, A4 => n3169
                           , ZN => n3156);
   U5000 : OAI221_X1 port map( B1 => n859, B2 => n2272, C1 => n825, C2 => n2273
                           , A => n3170, ZN => n3169);
   U5001 : AOI22_X1 port map( A1 => n2275, A2 => pc_target_10_13_port, B1 => 
                           n2276, B2 => pc_target_11_13_port, ZN => n3170);
   U5004 : OAI221_X1 port map( B1 => n721, B2 => n2277, C1 => n687, C2 => n2278
                           , A => n3171, ZN => n3168);
   U5005 : AOI22_X1 port map( A1 => n2280, A2 => pc_target_14_13_port, B1 => 
                           n2281, B2 => pc_target_15_13_port, ZN => n3171);
   U5008 : OAI221_X1 port map( B1 => n1133, B2 => n2282, C1 => n1099, C2 => 
                           n2283, A => n3172, ZN => n3167);
   U5009 : AOI22_X1 port map( A1 => n2285, A2 => pc_target_2_13_port, B1 => 
                           n2286, B2 => pc_target_3_13_port, ZN => n3172);
   U5012 : OAI221_X1 port map( B1 => n996, B2 => n2287, C1 => n962, C2 => n2288
                           , A => n3173, ZN => n3166);
   U5013 : AOI22_X1 port map( A1 => n2290, A2 => pc_target_6_13_port, B1 => 
                           n2291, B2 => pc_target_7_13_port, ZN => n3173);
   U5016 : NAND2_X1 port map( A1 => n3174, A2 => n3175, ZN => N113);
   U5017 : NOR4_X1 port map( A1 => n3176, A2 => n3177, A3 => n3178, A4 => n3179
                           , ZN => n3175);
   U5018 : OAI221_X1 port map( B1 => n292, B2 => n2248, C1 => n258, C2 => n2249
                           , A => n3180, ZN => n3179);
   U5019 : AOI22_X1 port map( A1 => n2251, A2 => pc_target_26_14_port, B1 => 
                           n2252, B2 => pc_target_27_14_port, ZN => n3180);
   U5022 : OAI221_X1 port map( B1 => n152, B2 => n2253, C1 => n94, C2 => n2254,
                           A => n3181, ZN => n3178);
   U5023 : AOI22_X1 port map( A1 => n2256, A2 => pc_target_30_14_port, B1 => 
                           n2257, B2 => pc_target_31_14_port, ZN => n3181);
   U5026 : OAI221_X1 port map( B1 => n568, B2 => n2258, C1 => n534, C2 => n2259
                           , A => n3182, ZN => n3177);
   U5027 : AOI22_X1 port map( A1 => n2261, A2 => pc_target_18_14_port, B1 => 
                           n2262, B2 => pc_target_19_14_port, ZN => n3182);
   U5030 : OAI221_X1 port map( B1 => n362, B2 => n2263, C1 => n327, C2 => n2264
                           , A => n3183, ZN => n3176);
   U5031 : AOI22_X1 port map( A1 => n2266, A2 => pc_target_20_14_port, B1 => 
                           n2267, B2 => pc_target_21_14_port, ZN => n3183);
   U5034 : NOR4_X1 port map( A1 => n3184, A2 => n3185, A3 => n3186, A4 => n3187
                           , ZN => n3174);
   U5035 : OAI221_X1 port map( B1 => n845, B2 => n2272, C1 => n811, C2 => n2273
                           , A => n3188, ZN => n3187);
   U5036 : AOI22_X1 port map( A1 => n2275, A2 => pc_target_10_14_port, B1 => 
                           n2276, B2 => pc_target_11_14_port, ZN => n3188);
   U5039 : OAI221_X1 port map( B1 => n707, B2 => n2277, C1 => n673, C2 => n2278
                           , A => n3189, ZN => n3186);
   U5040 : AOI22_X1 port map( A1 => n2280, A2 => pc_target_14_14_port, B1 => 
                           n2281, B2 => pc_target_15_14_port, ZN => n3189);
   U5043 : OAI221_X1 port map( B1 => n1119, B2 => n2282, C1 => n1085, C2 => 
                           n2283, A => n3190, ZN => n3185);
   U5044 : AOI22_X1 port map( A1 => n2285, A2 => pc_target_2_14_port, B1 => 
                           n2286, B2 => pc_target_3_14_port, ZN => n3190);
   U5047 : OAI221_X1 port map( B1 => n982, B2 => n2287, C1 => n948, C2 => n2288
                           , A => n3191, ZN => n3184);
   U5048 : AOI22_X1 port map( A1 => n2290, A2 => pc_target_6_14_port, B1 => 
                           n2291, B2 => pc_target_7_14_port, ZN => n3191);
   U5051 : NAND2_X1 port map( A1 => n3192, A2 => n3193, ZN => N112);
   U5052 : NOR4_X1 port map( A1 => n3194, A2 => n3195, A3 => n3196, A4 => n3197
                           , ZN => n3193);
   U5053 : OAI221_X1 port map( B1 => n307, B2 => n2248, C1 => n273, C2 => n2249
                           , A => n3198, ZN => n3197);
   U5054 : AOI22_X1 port map( A1 => n2251, A2 => pc_target_26_15_port, B1 => 
                           n2252, B2 => pc_target_27_15_port, ZN => n3198);
   U5057 : OAI221_X1 port map( B1 => n167, B2 => n2253, C1 => n124_port, C2 => 
                           n2254, A => n3199, ZN => n3196);
   U5058 : AOI22_X1 port map( A1 => n2256, A2 => pc_target_30_15_port, B1 => 
                           n2257, B2 => pc_target_31_15_port, ZN => n3199);
   U5061 : OAI221_X1 port map( B1 => n583, B2 => n2258, C1 => n549, C2 => n2259
                           , A => n3200, ZN => n3195);
   U5062 : AOI22_X1 port map( A1 => n2261, A2 => pc_target_18_15_port, B1 => 
                           n2262, B2 => pc_target_19_15_port, ZN => n3200);
   U5065 : OAI221_X1 port map( B1 => n377, B2 => n2263, C1 => n342, C2 => n2264
                           , A => n3201, ZN => n3194);
   U5066 : AOI22_X1 port map( A1 => n2266, A2 => pc_target_20_15_port, B1 => 
                           n2267, B2 => pc_target_21_15_port, ZN => n3201);
   U5069 : NOR4_X1 port map( A1 => n3202, A2 => n3203, A3 => n3204, A4 => n3205
                           , ZN => n3192);
   U5070 : OAI221_X1 port map( B1 => n860, B2 => n2272, C1 => n826, C2 => n2273
                           , A => n3206, ZN => n3205);
   U5071 : AOI22_X1 port map( A1 => n2275, A2 => pc_target_10_15_port, B1 => 
                           n2276, B2 => pc_target_11_15_port, ZN => n3206);
   U5074 : OAI221_X1 port map( B1 => n722, B2 => n2277, C1 => n688, C2 => n2278
                           , A => n3207, ZN => n3204);
   U5075 : AOI22_X1 port map( A1 => n2280, A2 => pc_target_14_15_port, B1 => 
                           n2281, B2 => pc_target_15_15_port, ZN => n3207);
   U5078 : OAI221_X1 port map( B1 => n1134, B2 => n2282, C1 => n1100, C2 => 
                           n2283, A => n3208, ZN => n3203);
   U5079 : AOI22_X1 port map( A1 => n2285, A2 => pc_target_2_15_port, B1 => 
                           n2286, B2 => pc_target_3_15_port, ZN => n3208);
   U5082 : OAI221_X1 port map( B1 => n997, B2 => n2287, C1 => n963, C2 => n2288
                           , A => n3209, ZN => n3202);
   U5083 : AOI22_X1 port map( A1 => n2290, A2 => pc_target_6_15_port, B1 => 
                           n2291, B2 => pc_target_7_15_port, ZN => n3209);
   U5086 : NAND2_X1 port map( A1 => n3210, A2 => n3211, ZN => N111);
   U5087 : NOR4_X1 port map( A1 => n3212, A2 => n3213, A3 => n3214, A4 => n3215
                           , ZN => n3211);
   U5088 : OAI221_X1 port map( B1 => n291, B2 => n2248, C1 => n257, C2 => n2249
                           , A => n3216, ZN => n3215);
   U5089 : AOI22_X1 port map( A1 => n2251, A2 => pc_target_26_16_port, B1 => 
                           n2252, B2 => pc_target_27_16_port, ZN => n3216);
   U5092 : OAI221_X1 port map( B1 => n151, B2 => n2253, C1 => n92, C2 => n2254,
                           A => n3217, ZN => n3214);
   U5093 : AOI22_X1 port map( A1 => n2256, A2 => pc_target_30_16_port, B1 => 
                           n2257, B2 => pc_target_31_16_port, ZN => n3217);
   U5096 : OAI221_X1 port map( B1 => n567, B2 => n2258, C1 => n533, C2 => n2259
                           , A => n3218, ZN => n3213);
   U5097 : AOI22_X1 port map( A1 => n2261, A2 => pc_target_18_16_port, B1 => 
                           n2262, B2 => pc_target_19_16_port, ZN => n3218);
   U5100 : OAI221_X1 port map( B1 => n361, B2 => n2263, C1 => n326, C2 => n2264
                           , A => n3219, ZN => n3212);
   U5101 : AOI22_X1 port map( A1 => n2266, A2 => pc_target_20_16_port, B1 => 
                           n2267, B2 => pc_target_21_16_port, ZN => n3219);
   U5104 : NOR4_X1 port map( A1 => n3220, A2 => n3221, A3 => n3222, A4 => n3223
                           , ZN => n3210);
   U5105 : OAI221_X1 port map( B1 => n844, B2 => n2272, C1 => n810, C2 => n2273
                           , A => n3224, ZN => n3223);
   U5106 : AOI22_X1 port map( A1 => n2275, A2 => pc_target_10_16_port, B1 => 
                           n2276, B2 => pc_target_11_16_port, ZN => n3224);
   U5109 : OAI221_X1 port map( B1 => n706, B2 => n2277, C1 => n672, C2 => n2278
                           , A => n3225, ZN => n3222);
   U5110 : AOI22_X1 port map( A1 => n2280, A2 => pc_target_14_16_port, B1 => 
                           n2281, B2 => pc_target_15_16_port, ZN => n3225);
   U5113 : OAI221_X1 port map( B1 => n1118, B2 => n2282, C1 => n1084, C2 => 
                           n2283, A => n3226, ZN => n3221);
   U5114 : AOI22_X1 port map( A1 => n2285, A2 => pc_target_2_16_port, B1 => 
                           n2286, B2 => pc_target_3_16_port, ZN => n3226);
   U5117 : OAI221_X1 port map( B1 => n981, B2 => n2287, C1 => n947, C2 => n2288
                           , A => n3227, ZN => n3220);
   U5118 : AOI22_X1 port map( A1 => n2290, A2 => pc_target_6_16_port, B1 => 
                           n2291, B2 => pc_target_7_16_port, ZN => n3227);
   U5121 : NAND2_X1 port map( A1 => n3228, A2 => n3229, ZN => N110);
   U5122 : NOR4_X1 port map( A1 => n3230, A2 => n3231, A3 => n3232, A4 => n3233
                           , ZN => n3229);
   U5123 : OAI221_X1 port map( B1 => n308, B2 => n2248, C1 => n274, C2 => n2249
                           , A => n3234, ZN => n3233);
   U5124 : AOI22_X1 port map( A1 => n2251, A2 => pc_target_26_17_port, B1 => 
                           n2252, B2 => pc_target_27_17_port, ZN => n3234);
   U5127 : OAI221_X1 port map( B1 => n168, B2 => n2253, C1 => n126_port, C2 => 
                           n2254, A => n3235, ZN => n3232);
   U5128 : AOI22_X1 port map( A1 => n2256, A2 => pc_target_30_17_port, B1 => 
                           n2257, B2 => pc_target_31_17_port, ZN => n3235);
   U5131 : OAI221_X1 port map( B1 => n584, B2 => n2258, C1 => n550, C2 => n2259
                           , A => n3236, ZN => n3231);
   U5132 : AOI22_X1 port map( A1 => n2261, A2 => pc_target_18_17_port, B1 => 
                           n2262, B2 => pc_target_19_17_port, ZN => n3236);
   U5135 : OAI221_X1 port map( B1 => n378, B2 => n2263, C1 => n343, C2 => n2264
                           , A => n3237, ZN => n3230);
   U5136 : AOI22_X1 port map( A1 => n2266, A2 => pc_target_20_17_port, B1 => 
                           n2267, B2 => pc_target_21_17_port, ZN => n3237);
   U5139 : NOR4_X1 port map( A1 => n3238, A2 => n3239, A3 => n3240, A4 => n3241
                           , ZN => n3228);
   U5140 : OAI221_X1 port map( B1 => n861, B2 => n2272, C1 => n827, C2 => n2273
                           , A => n3242, ZN => n3241);
   U5141 : AOI22_X1 port map( A1 => n2275, A2 => pc_target_10_17_port, B1 => 
                           n2276, B2 => pc_target_11_17_port, ZN => n3242);
   U5144 : OAI221_X1 port map( B1 => n723, B2 => n2277, C1 => n689, C2 => n2278
                           , A => n3243, ZN => n3240);
   U5145 : AOI22_X1 port map( A1 => n2280, A2 => pc_target_14_17_port, B1 => 
                           n2281, B2 => pc_target_15_17_port, ZN => n3243);
   U5148 : OAI221_X1 port map( B1 => n1135, B2 => n2282, C1 => n1101, C2 => 
                           n2283, A => n3244, ZN => n3239);
   U5149 : AOI22_X1 port map( A1 => n2285, A2 => pc_target_2_17_port, B1 => 
                           n2286, B2 => pc_target_3_17_port, ZN => n3244);
   U5152 : OAI221_X1 port map( B1 => n998, B2 => n2287, C1 => n964, C2 => n2288
                           , A => n3245, ZN => n3238);
   U5153 : AOI22_X1 port map( A1 => n2290, A2 => pc_target_6_17_port, B1 => 
                           n2291, B2 => pc_target_7_17_port, ZN => n3245);
   U5156 : NAND2_X1 port map( A1 => n3246, A2 => n3247, ZN => N109);
   U5157 : NOR4_X1 port map( A1 => n3248, A2 => n3249, A3 => n3250, A4 => n3251
                           , ZN => n3247);
   U5158 : OAI221_X1 port map( B1 => n290, B2 => n2248, C1 => n256, C2 => n2249
                           , A => n3252, ZN => n3251);
   U5159 : AOI22_X1 port map( A1 => n2251, A2 => pc_target_26_18_port, B1 => 
                           n2252, B2 => pc_target_27_18_port, ZN => n3252);
   U5162 : OAI221_X1 port map( B1 => n150, B2 => n2253, C1 => n90, C2 => n2254,
                           A => n3253, ZN => n3250);
   U5163 : AOI22_X1 port map( A1 => n2256, A2 => pc_target_30_18_port, B1 => 
                           n2257, B2 => pc_target_31_18_port, ZN => n3253);
   U5166 : OAI221_X1 port map( B1 => n566, B2 => n2258, C1 => n532, C2 => n2259
                           , A => n3254, ZN => n3249);
   U5167 : AOI22_X1 port map( A1 => n2261, A2 => pc_target_18_18_port, B1 => 
                           n2262, B2 => pc_target_19_18_port, ZN => n3254);
   U5170 : OAI221_X1 port map( B1 => n360, B2 => n2263, C1 => n325, C2 => n2264
                           , A => n3255, ZN => n3248);
   U5171 : AOI22_X1 port map( A1 => n2266, A2 => pc_target_20_18_port, B1 => 
                           n2267, B2 => pc_target_21_18_port, ZN => n3255);
   U5174 : NOR4_X1 port map( A1 => n3256, A2 => n3257, A3 => n3258, A4 => n3259
                           , ZN => n3246);
   U5175 : OAI221_X1 port map( B1 => n843, B2 => n2272, C1 => n809, C2 => n2273
                           , A => n3260, ZN => n3259);
   U5176 : AOI22_X1 port map( A1 => n2275, A2 => pc_target_10_18_port, B1 => 
                           n2276, B2 => pc_target_11_18_port, ZN => n3260);
   U5179 : OAI221_X1 port map( B1 => n705, B2 => n2277, C1 => n671, C2 => n2278
                           , A => n3261, ZN => n3258);
   U5180 : AOI22_X1 port map( A1 => n2280, A2 => pc_target_14_18_port, B1 => 
                           n2281, B2 => pc_target_15_18_port, ZN => n3261);
   U5183 : OAI221_X1 port map( B1 => n1117, B2 => n2282, C1 => n1083, C2 => 
                           n2283, A => n3262, ZN => n3257);
   U5184 : AOI22_X1 port map( A1 => n2285, A2 => pc_target_2_18_port, B1 => 
                           n2286, B2 => pc_target_3_18_port, ZN => n3262);
   U5187 : OAI221_X1 port map( B1 => n980, B2 => n2287, C1 => n946, C2 => n2288
                           , A => n3263, ZN => n3256);
   U5188 : AOI22_X1 port map( A1 => n2290, A2 => pc_target_6_18_port, B1 => 
                           n2291, B2 => pc_target_7_18_port, ZN => n3263);
   U5191 : NAND2_X1 port map( A1 => n3264, A2 => n3265, ZN => N108);
   U5192 : NOR4_X1 port map( A1 => n3266, A2 => n3267, A3 => n3268, A4 => n3269
                           , ZN => n3265);
   U5193 : OAI221_X1 port map( B1 => n309, B2 => n2248, C1 => n275, C2 => n2249
                           , A => n3270, ZN => n3269);
   U5194 : AOI22_X1 port map( A1 => n2251, A2 => pc_target_26_19_port, B1 => 
                           n2252, B2 => pc_target_27_19_port, ZN => n3270);
   U5197 : OAI221_X1 port map( B1 => n169, B2 => n2253, C1 => n128, C2 => n2254
                           , A => n3271, ZN => n3268);
   U5198 : AOI22_X1 port map( A1 => n2256, A2 => pc_target_30_19_port, B1 => 
                           n2257, B2 => pc_target_31_19_port, ZN => n3271);
   U5201 : OAI221_X1 port map( B1 => n585, B2 => n2258, C1 => n551, C2 => n2259
                           , A => n3272, ZN => n3267);
   U5202 : AOI22_X1 port map( A1 => n2261, A2 => pc_target_18_19_port, B1 => 
                           n2262, B2 => pc_target_19_19_port, ZN => n3272);
   U5205 : OAI221_X1 port map( B1 => n379, B2 => n2263, C1 => n344, C2 => n2264
                           , A => n3273, ZN => n3266);
   U5206 : AOI22_X1 port map( A1 => n2266, A2 => pc_target_20_19_port, B1 => 
                           n2267, B2 => pc_target_21_19_port, ZN => n3273);
   U5209 : NOR4_X1 port map( A1 => n3274, A2 => n3275, A3 => n3276, A4 => n3277
                           , ZN => n3264);
   U5210 : OAI221_X1 port map( B1 => n862, B2 => n2272, C1 => n828, C2 => n2273
                           , A => n3278, ZN => n3277);
   U5211 : AOI22_X1 port map( A1 => n2275, A2 => pc_target_10_19_port, B1 => 
                           n2276, B2 => pc_target_11_19_port, ZN => n3278);
   U5214 : OAI221_X1 port map( B1 => n724, B2 => n2277, C1 => n690, C2 => n2278
                           , A => n3279, ZN => n3276);
   U5215 : AOI22_X1 port map( A1 => n2280, A2 => pc_target_14_19_port, B1 => 
                           n2281, B2 => pc_target_15_19_port, ZN => n3279);
   U5218 : OAI221_X1 port map( B1 => n1136, B2 => n2282, C1 => n1102, C2 => 
                           n2283, A => n3280, ZN => n3275);
   U5219 : AOI22_X1 port map( A1 => n2285, A2 => pc_target_2_19_port, B1 => 
                           n2286, B2 => pc_target_3_19_port, ZN => n3280);
   U5222 : OAI221_X1 port map( B1 => n999, B2 => n2287, C1 => n965, C2 => n2288
                           , A => n3281, ZN => n3274);
   U5223 : AOI22_X1 port map( A1 => n2290, A2 => pc_target_6_19_port, B1 => 
                           n2291, B2 => pc_target_7_19_port, ZN => n3281);
   U5226 : NAND2_X1 port map( A1 => n3282, A2 => n3283, ZN => N107);
   U5227 : NOR4_X1 port map( A1 => n3284, A2 => n3285, A3 => n3286, A4 => n3287
                           , ZN => n3283);
   U5228 : OAI221_X1 port map( B1 => n289, B2 => n2248, C1 => n255, C2 => n2249
                           , A => n3288, ZN => n3287);
   U5229 : AOI22_X1 port map( A1 => n2251, A2 => pc_target_26_20_port, B1 => 
                           n2252, B2 => pc_target_27_20_port, ZN => n3288);
   U5232 : OAI221_X1 port map( B1 => n149, B2 => n2253, C1 => n88, C2 => n2254,
                           A => n3289, ZN => n3286);
   U5233 : AOI22_X1 port map( A1 => n2256, A2 => pc_target_30_20_port, B1 => 
                           n2257, B2 => pc_target_31_20_port, ZN => n3289);
   U5236 : OAI221_X1 port map( B1 => n565, B2 => n2258, C1 => n531, C2 => n2259
                           , A => n3290, ZN => n3285);
   U5237 : AOI22_X1 port map( A1 => n2261, A2 => pc_target_18_20_port, B1 => 
                           n2262, B2 => pc_target_19_20_port, ZN => n3290);
   U5240 : OAI221_X1 port map( B1 => n359, B2 => n2263, C1 => n324, C2 => n2264
                           , A => n3291, ZN => n3284);
   U5241 : AOI22_X1 port map( A1 => n2266, A2 => pc_target_20_20_port, B1 => 
                           n2267, B2 => pc_target_21_20_port, ZN => n3291);
   U5244 : NOR4_X1 port map( A1 => n3292, A2 => n3293, A3 => n3294, A4 => n3295
                           , ZN => n3282);
   U5245 : OAI221_X1 port map( B1 => n842, B2 => n2272, C1 => n808, C2 => n2273
                           , A => n3296, ZN => n3295);
   U5246 : AOI22_X1 port map( A1 => n2275, A2 => pc_target_10_20_port, B1 => 
                           n2276, B2 => pc_target_11_20_port, ZN => n3296);
   U5249 : OAI221_X1 port map( B1 => n704, B2 => n2277, C1 => n670, C2 => n2278
                           , A => n3297, ZN => n3294);
   U5250 : AOI22_X1 port map( A1 => n2280, A2 => pc_target_14_20_port, B1 => 
                           n2281, B2 => pc_target_15_20_port, ZN => n3297);
   U5253 : OAI221_X1 port map( B1 => n1116, B2 => n2282, C1 => n1082, C2 => 
                           n2283, A => n3298, ZN => n3293);
   U5254 : AOI22_X1 port map( A1 => n2285, A2 => pc_target_2_20_port, B1 => 
                           n2286, B2 => pc_target_3_20_port, ZN => n3298);
   U5257 : OAI221_X1 port map( B1 => n979, B2 => n2287, C1 => n945, C2 => n2288
                           , A => n3299, ZN => n3292);
   U5258 : AOI22_X1 port map( A1 => n2290, A2 => pc_target_6_20_port, B1 => 
                           n2291, B2 => pc_target_7_20_port, ZN => n3299);
   U5261 : NAND2_X1 port map( A1 => n3300, A2 => n3301, ZN => N106);
   U5262 : NOR4_X1 port map( A1 => n3302, A2 => n3303, A3 => n3304, A4 => n3305
                           , ZN => n3301);
   U5263 : OAI221_X1 port map( B1 => n310, B2 => n2248, C1 => n276, C2 => n2249
                           , A => n3306, ZN => n3305);
   U5264 : AOI22_X1 port map( A1 => n2251, A2 => pc_target_26_21_port, B1 => 
                           n2252, B2 => pc_target_27_21_port, ZN => n3306);
   U5267 : OAI221_X1 port map( B1 => n170, B2 => n2253, C1 => n130, C2 => n2254
                           , A => n3307, ZN => n3304);
   U5268 : AOI22_X1 port map( A1 => n2256, A2 => pc_target_30_21_port, B1 => 
                           n2257, B2 => pc_target_31_21_port, ZN => n3307);
   U5271 : OAI221_X1 port map( B1 => n586, B2 => n2258, C1 => n552, C2 => n2259
                           , A => n3308, ZN => n3303);
   U5272 : AOI22_X1 port map( A1 => n2261, A2 => pc_target_18_21_port, B1 => 
                           n2262, B2 => pc_target_19_21_port, ZN => n3308);
   U5275 : OAI221_X1 port map( B1 => n380, B2 => n2263, C1 => n345, C2 => n2264
                           , A => n3309, ZN => n3302);
   U5276 : AOI22_X1 port map( A1 => n2266, A2 => pc_target_20_21_port, B1 => 
                           n2267, B2 => pc_target_21_21_port, ZN => n3309);
   U5279 : NOR4_X1 port map( A1 => n3310, A2 => n3311, A3 => n3312, A4 => n3313
                           , ZN => n3300);
   U5280 : OAI221_X1 port map( B1 => n863, B2 => n2272, C1 => n829, C2 => n2273
                           , A => n3314, ZN => n3313);
   U5281 : AOI22_X1 port map( A1 => n2275, A2 => pc_target_10_21_port, B1 => 
                           n2276, B2 => pc_target_11_21_port, ZN => n3314);
   U5284 : OAI221_X1 port map( B1 => n725, B2 => n2277, C1 => n691, C2 => n2278
                           , A => n3315, ZN => n3312);
   U5285 : AOI22_X1 port map( A1 => n2280, A2 => pc_target_14_21_port, B1 => 
                           n2281, B2 => pc_target_15_21_port, ZN => n3315);
   U5288 : OAI221_X1 port map( B1 => n1137, B2 => n2282, C1 => n1103, C2 => 
                           n2283, A => n3316, ZN => n3311);
   U5289 : AOI22_X1 port map( A1 => n2285, A2 => pc_target_2_21_port, B1 => 
                           n2286, B2 => pc_target_3_21_port, ZN => n3316);
   U5292 : OAI221_X1 port map( B1 => n1000, B2 => n2287, C1 => n966, C2 => 
                           n2288, A => n3317, ZN => n3310);
   U5293 : AOI22_X1 port map( A1 => n2290, A2 => pc_target_6_21_port, B1 => 
                           n2291, B2 => pc_target_7_21_port, ZN => n3317);
   U5296 : NAND2_X1 port map( A1 => n3318, A2 => n3319, ZN => N105);
   U5297 : NOR4_X1 port map( A1 => n3320, A2 => n3321, A3 => n3322, A4 => n3323
                           , ZN => n3319);
   U5298 : OAI221_X1 port map( B1 => n288, B2 => n2248, C1 => n254, C2 => n2249
                           , A => n3324, ZN => n3323);
   U5299 : AOI22_X1 port map( A1 => n2251, A2 => pc_target_26_22_port, B1 => 
                           n2252, B2 => pc_target_27_22_port, ZN => n3324);
   U5302 : OAI221_X1 port map( B1 => n148, B2 => n2253, C1 => n86, C2 => n2254,
                           A => n3325, ZN => n3322);
   U5303 : AOI22_X1 port map( A1 => n2256, A2 => pc_target_30_22_port, B1 => 
                           n2257, B2 => pc_target_31_22_port, ZN => n3325);
   U5306 : OAI221_X1 port map( B1 => n564, B2 => n2258, C1 => n530, C2 => n2259
                           , A => n3326, ZN => n3321);
   U5307 : AOI22_X1 port map( A1 => n2261, A2 => pc_target_18_22_port, B1 => 
                           n2262, B2 => pc_target_19_22_port, ZN => n3326);
   U5310 : OAI221_X1 port map( B1 => n358, B2 => n2263, C1 => n323, C2 => n2264
                           , A => n3327, ZN => n3320);
   U5311 : AOI22_X1 port map( A1 => n2266, A2 => pc_target_20_22_port, B1 => 
                           n2267, B2 => pc_target_21_22_port, ZN => n3327);
   U5314 : NOR4_X1 port map( A1 => n3328, A2 => n3329, A3 => n3330, A4 => n3331
                           , ZN => n3318);
   U5315 : OAI221_X1 port map( B1 => n841, B2 => n2272, C1 => n807, C2 => n2273
                           , A => n3332, ZN => n3331);
   U5316 : AOI22_X1 port map( A1 => n2275, A2 => pc_target_10_22_port, B1 => 
                           n2276, B2 => pc_target_11_22_port, ZN => n3332);
   U5319 : OAI221_X1 port map( B1 => n703, B2 => n2277, C1 => n669, C2 => n2278
                           , A => n3333, ZN => n3330);
   U5320 : AOI22_X1 port map( A1 => n2280, A2 => pc_target_14_22_port, B1 => 
                           n2281, B2 => pc_target_15_22_port, ZN => n3333);
   U5323 : OAI221_X1 port map( B1 => n1115, B2 => n2282, C1 => n1081, C2 => 
                           n2283, A => n3334, ZN => n3329);
   U5324 : AOI22_X1 port map( A1 => n2285, A2 => pc_target_2_22_port, B1 => 
                           n2286, B2 => pc_target_3_22_port, ZN => n3334);
   U5327 : OAI221_X1 port map( B1 => n978, B2 => n2287, C1 => n944, C2 => n2288
                           , A => n3335, ZN => n3328);
   U5328 : AOI22_X1 port map( A1 => n2290, A2 => pc_target_6_22_port, B1 => 
                           n2291, B2 => pc_target_7_22_port, ZN => n3335);
   U5331 : NAND2_X1 port map( A1 => n3336, A2 => n3337, ZN => N104);
   U5332 : NOR4_X1 port map( A1 => n3338, A2 => n3339, A3 => n3340, A4 => n3341
                           , ZN => n3337);
   U5333 : OAI221_X1 port map( B1 => n311, B2 => n2248, C1 => n277, C2 => n2249
                           , A => n3342, ZN => n3341);
   U5334 : AOI22_X1 port map( A1 => n2251, A2 => pc_target_26_23_port, B1 => 
                           n2252, B2 => pc_target_27_23_port, ZN => n3342);
   U5337 : OAI221_X1 port map( B1 => n171, B2 => n2253, C1 => n132, C2 => n2254
                           , A => n3343, ZN => n3340);
   U5338 : AOI22_X1 port map( A1 => n2256, A2 => pc_target_30_23_port, B1 => 
                           n2257, B2 => pc_target_31_23_port, ZN => n3343);
   U5341 : OAI221_X1 port map( B1 => n587, B2 => n2258, C1 => n553, C2 => n2259
                           , A => n3344, ZN => n3339);
   U5342 : AOI22_X1 port map( A1 => n2261, A2 => pc_target_18_23_port, B1 => 
                           n2262, B2 => pc_target_19_23_port, ZN => n3344);
   U5345 : OAI221_X1 port map( B1 => n381, B2 => n2263, C1 => n346, C2 => n2264
                           , A => n3345, ZN => n3338);
   U5346 : AOI22_X1 port map( A1 => n2266, A2 => pc_target_20_23_port, B1 => 
                           n2267, B2 => pc_target_21_23_port, ZN => n3345);
   U5349 : NOR4_X1 port map( A1 => n3346, A2 => n3347, A3 => n3348, A4 => n3349
                           , ZN => n3336);
   U5350 : OAI221_X1 port map( B1 => n864, B2 => n2272, C1 => n830, C2 => n2273
                           , A => n3350, ZN => n3349);
   U5351 : AOI22_X1 port map( A1 => n2275, A2 => pc_target_10_23_port, B1 => 
                           n2276, B2 => pc_target_11_23_port, ZN => n3350);
   U5354 : OAI221_X1 port map( B1 => n726, B2 => n2277, C1 => n692, C2 => n2278
                           , A => n3351, ZN => n3348);
   U5355 : AOI22_X1 port map( A1 => n2280, A2 => pc_target_14_23_port, B1 => 
                           n2281, B2 => pc_target_15_23_port, ZN => n3351);
   U5358 : OAI221_X1 port map( B1 => n1138, B2 => n2282, C1 => n1104, C2 => 
                           n2283, A => n3352, ZN => n3347);
   U5359 : AOI22_X1 port map( A1 => n2285, A2 => pc_target_2_23_port, B1 => 
                           n2286, B2 => pc_target_3_23_port, ZN => n3352);
   U5362 : OAI221_X1 port map( B1 => n1001, B2 => n2287, C1 => n967, C2 => 
                           n2288, A => n3353, ZN => n3346);
   U5363 : AOI22_X1 port map( A1 => n2290, A2 => pc_target_6_23_port, B1 => 
                           n2291, B2 => pc_target_7_23_port, ZN => n3353);
   U5366 : NAND2_X1 port map( A1 => n3354, A2 => n3355, ZN => N103);
   U5367 : NOR4_X1 port map( A1 => n3356, A2 => n3357, A3 => n3358, A4 => n3359
                           , ZN => n3355);
   U5368 : OAI221_X1 port map( B1 => n287, B2 => n2248, C1 => n253, C2 => n2249
                           , A => n3360, ZN => n3359);
   U5369 : AOI22_X1 port map( A1 => n2251, A2 => pc_target_26_24_port, B1 => 
                           n2252, B2 => pc_target_27_24_port, ZN => n3360);
   U5372 : OAI221_X1 port map( B1 => n147, B2 => n2253, C1 => n84, C2 => n2254,
                           A => n3361, ZN => n3358);
   U5373 : AOI22_X1 port map( A1 => n2256, A2 => pc_target_30_24_port, B1 => 
                           n2257, B2 => pc_target_31_24_port, ZN => n3361);
   U5376 : OAI221_X1 port map( B1 => n563, B2 => n2258, C1 => n529, C2 => n2259
                           , A => n3362, ZN => n3357);
   U5377 : AOI22_X1 port map( A1 => n2261, A2 => pc_target_18_24_port, B1 => 
                           n2262, B2 => pc_target_19_24_port, ZN => n3362);
   U5380 : OAI221_X1 port map( B1 => n357, B2 => n2263, C1 => n322, C2 => n2264
                           , A => n3363, ZN => n3356);
   U5381 : AOI22_X1 port map( A1 => n2266, A2 => pc_target_20_24_port, B1 => 
                           n2267, B2 => pc_target_21_24_port, ZN => n3363);
   U5384 : NOR4_X1 port map( A1 => n3364, A2 => n3365, A3 => n3366, A4 => n3367
                           , ZN => n3354);
   U5385 : OAI221_X1 port map( B1 => n840, B2 => n2272, C1 => n806, C2 => n2273
                           , A => n3368, ZN => n3367);
   U5386 : AOI22_X1 port map( A1 => n2275, A2 => pc_target_10_24_port, B1 => 
                           n2276, B2 => pc_target_11_24_port, ZN => n3368);
   U5389 : OAI221_X1 port map( B1 => n702, B2 => n2277, C1 => n668, C2 => n2278
                           , A => n3369, ZN => n3366);
   U5390 : AOI22_X1 port map( A1 => n2280, A2 => pc_target_14_24_port, B1 => 
                           n2281, B2 => pc_target_15_24_port, ZN => n3369);
   U5393 : OAI221_X1 port map( B1 => n1114, B2 => n2282, C1 => n1080, C2 => 
                           n2283, A => n3370, ZN => n3365);
   U5394 : AOI22_X1 port map( A1 => n2285, A2 => pc_target_2_24_port, B1 => 
                           n2286, B2 => pc_target_3_24_port, ZN => n3370);
   U5397 : OAI221_X1 port map( B1 => n977, B2 => n2287, C1 => n943, C2 => n2288
                           , A => n3371, ZN => n3364);
   U5398 : AOI22_X1 port map( A1 => n2290, A2 => pc_target_6_24_port, B1 => 
                           n2291, B2 => pc_target_7_24_port, ZN => n3371);
   U5401 : NAND2_X1 port map( A1 => n3372, A2 => n3373, ZN => N102);
   U5402 : NOR4_X1 port map( A1 => n3374, A2 => n3375, A3 => n3376, A4 => n3377
                           , ZN => n3373);
   U5403 : OAI221_X1 port map( B1 => n312, B2 => n2248, C1 => n278, C2 => n2249
                           , A => n3378, ZN => n3377);
   U5404 : AOI22_X1 port map( A1 => n2251, A2 => pc_target_26_25_port, B1 => 
                           n2252, B2 => pc_target_27_25_port, ZN => n3378);
   U5407 : OAI221_X1 port map( B1 => n172, B2 => n2253, C1 => n134, C2 => n2254
                           , A => n3379, ZN => n3376);
   U5408 : AOI22_X1 port map( A1 => n2256, A2 => pc_target_30_25_port, B1 => 
                           n2257, B2 => pc_target_31_25_port, ZN => n3379);
   U5411 : OAI221_X1 port map( B1 => n588, B2 => n2258, C1 => n554, C2 => n2259
                           , A => n3380, ZN => n3375);
   U5412 : AOI22_X1 port map( A1 => n2261, A2 => pc_target_18_25_port, B1 => 
                           n2262, B2 => pc_target_19_25_port, ZN => n3380);
   U5415 : OAI221_X1 port map( B1 => n382, B2 => n2263, C1 => n347, C2 => n2264
                           , A => n3381, ZN => n3374);
   U5416 : AOI22_X1 port map( A1 => n2266, A2 => pc_target_20_25_port, B1 => 
                           n2267, B2 => pc_target_21_25_port, ZN => n3381);
   U5419 : NOR4_X1 port map( A1 => n3382, A2 => n3383, A3 => n3384, A4 => n3385
                           , ZN => n3372);
   U5420 : OAI221_X1 port map( B1 => n865, B2 => n2272, C1 => n831, C2 => n2273
                           , A => n3386, ZN => n3385);
   U5421 : AOI22_X1 port map( A1 => n2275, A2 => pc_target_10_25_port, B1 => 
                           n2276, B2 => pc_target_11_25_port, ZN => n3386);
   U5424 : OAI221_X1 port map( B1 => n727, B2 => n2277, C1 => n693, C2 => n2278
                           , A => n3387, ZN => n3384);
   U5425 : AOI22_X1 port map( A1 => n2280, A2 => pc_target_14_25_port, B1 => 
                           n2281, B2 => pc_target_15_25_port, ZN => n3387);
   U5428 : OAI221_X1 port map( B1 => n1139, B2 => n2282, C1 => n1105, C2 => 
                           n2283, A => n3388, ZN => n3383);
   U5429 : AOI22_X1 port map( A1 => n2285, A2 => pc_target_2_25_port, B1 => 
                           n2286, B2 => pc_target_3_25_port, ZN => n3388);
   U5432 : OAI221_X1 port map( B1 => n1002, B2 => n2287, C1 => n968, C2 => 
                           n2288, A => n3389, ZN => n3382);
   U5433 : AOI22_X1 port map( A1 => n2290, A2 => pc_target_6_25_port, B1 => 
                           n2291, B2 => pc_target_7_25_port, ZN => n3389);
   U5436 : NAND2_X1 port map( A1 => n3390, A2 => n3391, ZN => N101);
   U5437 : NOR4_X1 port map( A1 => n3392, A2 => n3393, A3 => n3394, A4 => n3395
                           , ZN => n3391);
   U5438 : OAI221_X1 port map( B1 => n286, B2 => n2248, C1 => n252, C2 => n2249
                           , A => n3396, ZN => n3395);
   U5439 : AOI22_X1 port map( A1 => n2251, A2 => pc_target_26_26_port, B1 => 
                           n2252, B2 => pc_target_27_26_port, ZN => n3396);
   U5442 : OAI221_X1 port map( B1 => n146, B2 => n2253, C1 => n82, C2 => n2254,
                           A => n3397, ZN => n3394);
   U5443 : AOI22_X1 port map( A1 => n2256, A2 => pc_target_30_26_port, B1 => 
                           n2257, B2 => pc_target_31_26_port, ZN => n3397);
   U5446 : OAI221_X1 port map( B1 => n562, B2 => n2258, C1 => n528, C2 => n2259
                           , A => n3398, ZN => n3393);
   U5447 : AOI22_X1 port map( A1 => n2261, A2 => pc_target_18_26_port, B1 => 
                           n2262, B2 => pc_target_19_26_port, ZN => n3398);
   U5450 : OAI221_X1 port map( B1 => n356, B2 => n2263, C1 => n321, C2 => n2264
                           , A => n3399, ZN => n3392);
   U5451 : AOI22_X1 port map( A1 => n2266, A2 => pc_target_20_26_port, B1 => 
                           n2267, B2 => pc_target_21_26_port, ZN => n3399);
   U5454 : NOR4_X1 port map( A1 => n3400, A2 => n3401, A3 => n3402, A4 => n3403
                           , ZN => n3390);
   U5455 : OAI221_X1 port map( B1 => n839, B2 => n2272, C1 => n805, C2 => n2273
                           , A => n3404, ZN => n3403);
   U5456 : AOI22_X1 port map( A1 => n2275, A2 => pc_target_10_26_port, B1 => 
                           n2276, B2 => pc_target_11_26_port, ZN => n3404);
   U5459 : OAI221_X1 port map( B1 => n701, B2 => n2277, C1 => n667, C2 => n2278
                           , A => n3405, ZN => n3402);
   U5460 : AOI22_X1 port map( A1 => n2280, A2 => pc_target_14_26_port, B1 => 
                           n2281, B2 => pc_target_15_26_port, ZN => n3405);
   U5463 : OAI221_X1 port map( B1 => n1113, B2 => n2282, C1 => n1079, C2 => 
                           n2283, A => n3406, ZN => n3401);
   U5464 : AOI22_X1 port map( A1 => n2285, A2 => pc_target_2_26_port, B1 => 
                           n2286, B2 => pc_target_3_26_port, ZN => n3406);
   U5467 : OAI221_X1 port map( B1 => n976, B2 => n2287, C1 => n942, C2 => n2288
                           , A => n3407, ZN => n3400);
   U5468 : AOI22_X1 port map( A1 => n2290, A2 => pc_target_6_26_port, B1 => 
                           n2291, B2 => pc_target_7_26_port, ZN => n3407);
   U5471 : NAND2_X1 port map( A1 => n3408, A2 => n3409, ZN => N100);
   U5472 : NOR4_X1 port map( A1 => n3410, A2 => n3411, A3 => n3412, A4 => n3413
                           , ZN => n3409);
   U5473 : OAI221_X1 port map( B1 => n313, B2 => n2248, C1 => n279, C2 => n2249
                           , A => n3414, ZN => n3413);
   U5474 : AOI22_X1 port map( A1 => n2251, A2 => pc_target_26_27_port, B1 => 
                           n2252, B2 => pc_target_27_27_port, ZN => n3414);
   U5481 : OAI221_X1 port map( B1 => n173, B2 => n2253, C1 => n136, C2 => n2254
                           , A => n3419, ZN => n3412);
   U5482 : AOI22_X1 port map( A1 => n2256, A2 => pc_target_30_27_port, B1 => 
                           n2257, B2 => pc_target_31_27_port, ZN => n3419);
   U5486 : AND3_X1 port map( A1 => PC_read(0), A2 => PC_read(4), A3 => 
                           PC_read(3), ZN => n3415);
   U5489 : AND3_X1 port map( A1 => PC_read(4), A2 => n3422, A3 => PC_read(3), 
                           ZN => n3417);
   U5491 : OAI221_X1 port map( B1 => n589, B2 => n2258, C1 => n555, C2 => n2259
                           , A => n3423, ZN => n3411);
   U5492 : AOI22_X1 port map( A1 => n2261, A2 => pc_target_18_27_port, B1 => 
                           n2262, B2 => pc_target_19_27_port, ZN => n3423);
   U5499 : OAI221_X1 port map( B1 => n383, B2 => n2263, C1 => n348, C2 => n2264
                           , A => n3426, ZN => n3410);
   U5500 : AOI22_X1 port map( A1 => n2266, A2 => pc_target_20_27_port, B1 => 
                           n2267, B2 => pc_target_21_27_port, ZN => n3426);
   U5504 : AND3_X1 port map( A1 => PC_read(4), A2 => n3427, A3 => PC_read(0), 
                           ZN => n3424);
   U5507 : AND3_X1 port map( A1 => n3422, A2 => n3427, A3 => PC_read(4), ZN => 
                           n3425);
   U5509 : NOR4_X1 port map( A1 => n3428, A2 => n3429, A3 => n3430, A4 => n3431
                           , ZN => n3408);
   U5510 : OAI221_X1 port map( B1 => n866, B2 => n2272, C1 => n832, C2 => n2273
                           , A => n3432, ZN => n3431);
   U5511 : AOI22_X1 port map( A1 => n2275, A2 => pc_target_10_27_port, B1 => 
                           n2276, B2 => pc_target_11_27_port, ZN => n3432);
   U5518 : OAI221_X1 port map( B1 => n728, B2 => n2277, C1 => n694, C2 => n2278
                           , A => n3435, ZN => n3430);
   U5519 : AOI22_X1 port map( A1 => n2280, A2 => pc_target_14_27_port, B1 => 
                           n2281, B2 => pc_target_15_27_port, ZN => n3435);
   U5527 : INV_X1 port map( A => PC_read(3), ZN => n3427);
   U5529 : OAI221_X1 port map( B1 => n1140, B2 => n2282, C1 => n1106, C2 => 
                           n2283, A => n3436, ZN => n3429);
   U5530 : AOI22_X1 port map( A1 => n2285, A2 => pc_target_2_27_port, B1 => 
                           n2286, B2 => pc_target_3_27_port, ZN => n3436);
   U5539 : OAI221_X1 port map( B1 => n1003, B2 => n2287, C1 => n969, C2 => 
                           n2288, A => n3440, ZN => n3428);
   U5540 : AOI22_X1 port map( A1 => n2290, A2 => pc_target_6_27_port, B1 => 
                           n2291, B2 => pc_target_7_27_port, ZN => n3440);
   U5544 : INV_X1 port map( A => PC_read(1), ZN => n3439);
   U5547 : INV_X1 port map( A => PC_read(0), ZN => n3422);
   U5551 : INV_X1 port map( A => PC_read(2), ZN => n3441);
   pc_target_reg_6_30_inst : DFFR_X2 port map( D => n6290, CK => Clk, RN => 
                           n3824, Q => pc_target_6_30_port, QN => n3502);
   pc_target_reg_6_28_inst : DFFR_X2 port map( D => n6291, CK => Clk, RN => 
                           n3825, Q => pc_target_6_28_port, QN => n3501);
   pc_target_reg_6_26_inst : DFFR_X2 port map( D => n6292, CK => Clk, RN => 
                           n3824, Q => pc_target_6_26_port, QN => n3500);
   pc_target_reg_6_24_inst : DFFR_X2 port map( D => n6293, CK => Clk, RN => 
                           n3823, Q => pc_target_6_24_port, QN => n3499);
   pc_target_reg_6_22_inst : DFFR_X2 port map( D => n6294, CK => Clk, RN => 
                           n3825, Q => pc_target_6_22_port, QN => n3498);
   pc_target_reg_6_20_inst : DFFR_X2 port map( D => n6295, CK => Clk, RN => 
                           n3825, Q => pc_target_6_20_port, QN => n3497);
   pc_target_reg_6_18_inst : DFFR_X2 port map( D => n6296, CK => Clk, RN => 
                           n3825, Q => pc_target_6_18_port, QN => n3496);
   pc_target_reg_6_16_inst : DFFR_X2 port map( D => n6297, CK => Clk, RN => 
                           n3824, Q => pc_target_6_16_port, QN => n3495);
   pc_target_reg_6_14_inst : DFFR_X2 port map( D => n6298, CK => Clk, RN => 
                           n3825, Q => pc_target_6_14_port, QN => n3494);
   pc_target_reg_6_12_inst : DFFR_X2 port map( D => n6299, CK => Clk, RN => 
                           n3825, Q => pc_target_6_12_port, QN => n3493);
   pc_target_reg_6_10_inst : DFFR_X2 port map( D => n6300, CK => Clk, RN => 
                           n3824, Q => pc_target_6_10_port, QN => n3492);
   pc_target_reg_6_8_inst : DFFR_X2 port map( D => n6301, CK => Clk, RN => 
                           n3825, Q => pc_target_6_8_port, QN => n3491);
   pc_target_reg_6_6_inst : DFFR_X2 port map( D => n6302, CK => Clk, RN => 
                           n3823, Q => pc_target_6_6_port, QN => n3490);
   pc_target_reg_6_4_inst : DFFR_X2 port map( D => n6303, CK => Clk, RN => 
                           n3824, Q => pc_target_6_4_port, QN => n3489);
   pc_target_reg_6_2_inst : DFFR_X2 port map( D => n6304, CK => Clk, RN => 
                           n3825, Q => pc_target_6_2_port, QN => n3488);
   pc_target_reg_6_0_inst : DFFR_X2 port map( D => n6305, CK => Clk, RN => 
                           n3824, Q => pc_target_6_0_port, QN => n3487);
   pc_target_reg_6_1_inst : DFFR_X2 port map( D => n6306, CK => Clk, RN => 
                           n3824, Q => pc_target_6_1_port, QN => n3486);
   pc_target_reg_6_3_inst : DFFR_X2 port map( D => n6307, CK => Clk, RN => 
                           n3824, Q => pc_target_6_3_port, QN => n3485);
   pc_target_reg_6_5_inst : DFFR_X2 port map( D => n6308, CK => Clk, RN => 
                           n3825, Q => pc_target_6_5_port, QN => n3484);
   pc_target_reg_6_7_inst : DFFR_X2 port map( D => n6309, CK => Clk, RN => 
                           n3826, Q => pc_target_6_7_port, QN => n3483);
   pc_target_reg_6_9_inst : DFFR_X2 port map( D => n6310, CK => Clk, RN => 
                           n3824, Q => pc_target_6_9_port, QN => n3482);
   pc_target_reg_6_11_inst : DFFR_X2 port map( D => n6311, CK => Clk, RN => 
                           n3826, Q => pc_target_6_11_port, QN => n3481);
   pc_target_reg_6_13_inst : DFFR_X2 port map( D => n6312, CK => Clk, RN => 
                           n3826, Q => pc_target_6_13_port, QN => n3480);
   pc_target_reg_6_15_inst : DFFR_X2 port map( D => n6313, CK => Clk, RN => 
                           n3824, Q => pc_target_6_15_port, QN => n3479);
   pc_target_reg_6_17_inst : DFFR_X2 port map( D => n6314, CK => Clk, RN => 
                           n3824, Q => pc_target_6_17_port, QN => n3478);
   pc_target_reg_6_19_inst : DFFR_X2 port map( D => n6315, CK => Clk, RN => 
                           n3826, Q => pc_target_6_19_port, QN => n3477);
   pc_target_reg_6_21_inst : DFFR_X2 port map( D => n6316, CK => Clk, RN => 
                           n3825, Q => pc_target_6_21_port, QN => n3476);
   pc_target_reg_6_23_inst : DFFR_X2 port map( D => n6317, CK => Clk, RN => 
                           n3826, Q => pc_target_6_23_port, QN => n3475);
   pc_target_reg_6_25_inst : DFFR_X2 port map( D => n6318, CK => Clk, RN => 
                           n3826, Q => pc_target_6_25_port, QN => n3474);
   pc_target_reg_6_27_inst : DFFR_X2 port map( D => n6319, CK => Clk, RN => 
                           n3825, Q => pc_target_6_27_port, QN => n3473);
   pc_target_reg_6_29_inst : DFFR_X2 port map( D => n6320, CK => Clk, RN => 
                           n3825, Q => pc_target_6_29_port, QN => n3472);
   pc_target_reg_6_31_inst : DFFR_X2 port map( D => n6321, CK => Clk, RN => 
                           n3822, Q => pc_target_6_31_port, QN => n3471);
   pc_target_reg_2_30_inst : DFFR_X2 port map( D => n6418, CK => Clk, RN => 
                           n3822, Q => pc_target_2_30_port, QN => n3470);
   pc_target_reg_2_28_inst : DFFR_X2 port map( D => n6419, CK => Clk, RN => 
                           n3822, Q => pc_target_2_28_port, QN => n3469);
   pc_target_reg_2_26_inst : DFFR_X2 port map( D => n6420, CK => Clk, RN => 
                           n3822, Q => pc_target_2_26_port, QN => n3468);
   pc_target_reg_2_24_inst : DFFR_X2 port map( D => n6421, CK => Clk, RN => 
                           n3822, Q => pc_target_2_24_port, QN => n3467);
   pc_target_reg_2_22_inst : DFFR_X2 port map( D => n6422, CK => Clk, RN => 
                           n3822, Q => pc_target_2_22_port, QN => n3466);
   pc_target_reg_2_20_inst : DFFR_X2 port map( D => n6423, CK => Clk, RN => 
                           n3822, Q => pc_target_2_20_port, QN => n3465);
   pc_target_reg_2_18_inst : DFFR_X2 port map( D => n6424, CK => Clk, RN => 
                           n3822, Q => pc_target_2_18_port, QN => n3464);
   pc_target_reg_2_16_inst : DFFR_X2 port map( D => n6425, CK => Clk, RN => 
                           n3822, Q => pc_target_2_16_port, QN => n3463);
   pc_target_reg_2_14_inst : DFFR_X2 port map( D => n6426, CK => Clk, RN => 
                           n3822, Q => pc_target_2_14_port, QN => n3462);
   pc_target_reg_2_12_inst : DFFR_X2 port map( D => n6427, CK => Clk, RN => 
                           n3822, Q => pc_target_2_12_port, QN => n3461);
   pc_target_reg_2_7_inst : DFFR_X2 port map( D => n6437, CK => Clk, RN => 
                           n3823, Q => pc_target_2_7_port, QN => n3460);
   pc_target_reg_2_11_inst : DFFR_X2 port map( D => n6439, CK => Clk, RN => 
                           n3823, Q => pc_target_2_11_port, QN => n3459);
   pc_target_reg_2_13_inst : DFFR_X2 port map( D => n6440, CK => Clk, RN => 
                           n3823, Q => pc_target_2_13_port, QN => n3458);
   pc_target_reg_2_15_inst : DFFR_X2 port map( D => n6441, CK => Clk, RN => 
                           n3822, Q => pc_target_2_15_port, QN => n3457);
   pc_target_reg_2_17_inst : DFFR_X2 port map( D => n6442, CK => Clk, RN => 
                           n3823, Q => pc_target_2_17_port, QN => n3456);
   pc_target_reg_2_19_inst : DFFR_X2 port map( D => n6443, CK => Clk, RN => 
                           n3823, Q => pc_target_2_19_port, QN => n3455);
   pc_target_reg_2_21_inst : DFFR_X2 port map( D => n6444, CK => Clk, RN => 
                           n3823, Q => pc_target_2_21_port, QN => n3454);
   pc_target_reg_2_23_inst : DFFR_X2 port map( D => n6445, CK => Clk, RN => 
                           n3823, Q => pc_target_2_23_port, QN => n3453);
   pc_target_reg_2_25_inst : DFFR_X2 port map( D => n6446, CK => Clk, RN => 
                           n3823, Q => pc_target_2_25_port, QN => n3452);
   pc_target_reg_2_27_inst : DFFR_X2 port map( D => n6447, CK => Clk, RN => 
                           n3823, Q => pc_target_2_27_port, QN => n3451);
   pc_target_reg_2_29_inst : DFFR_X2 port map( D => n6448, CK => Clk, RN => 
                           n3824, Q => pc_target_2_29_port, QN => n3450);
   pc_target_reg_2_31_inst : DFFR_X2 port map( D => n6449, CK => Clk, RN => 
                           n3823, Q => pc_target_2_31_port, QN => n3449);
   pc_target_reg_2_6_inst : DFFR_X1 port map( D => n6430, CK => Clk, RN => 
                           n3910, Q => pc_target_2_6_port, QN => n2435);
   pc_target_reg_2_5_inst : DFFR_X1 port map( D => n6436, CK => Clk, RN => 
                           n3910, Q => pc_target_2_5_port, QN => n2434);
   pc_target_reg_2_4_inst : DFFR_X1 port map( D => n6431, CK => Clk, RN => 
                           n3910, Q => pc_target_2_4_port, QN => n2433);
   pc_target_reg_2_2_inst : DFFR_X1 port map( D => n6432, CK => Clk, RN => 
                           n3910, Q => pc_target_2_2_port, QN => n2432);
   pc_target_reg_2_1_inst : DFFR_X1 port map( D => n6434, CK => Clk, RN => 
                           n3910, Q => pc_target_2_1_port, QN => n2431);
   pc_target_reg_2_0_inst : DFFR_X1 port map( D => n6433, CK => Clk, RN => 
                           n3827, Q => pc_target_2_0_port, QN => n2430);
   pc_lut_reg_14_3_inst : DFFR_X1 port map( D => n7075, CK => Clk, RN => n3911,
                           Q => pc_lut_14_3_port, QN => n2429);
   pc_lut_reg_14_2_inst : DFFR_X1 port map( D => n7072, CK => Clk, RN => n3911,
                           Q => pc_lut_14_2_port, QN => n2428);
   pc_lut_reg_14_1_inst : DFFR_X1 port map( D => n7074, CK => Clk, RN => n3911,
                           Q => pc_lut_14_1_port, QN => n2418);
   pc_lut_reg_15_3_inst : DFFR_X1 port map( D => n7043, CK => Clk, RN => n3911,
                           Q => pc_lut_15_3_port, QN => n2417);
   pc_lut_reg_15_2_inst : DFFR_X1 port map( D => n7040, CK => Clk, RN => n3912,
                           Q => pc_lut_15_2_port, QN => n2416);
   pc_lut_reg_15_1_inst : DFFR_X1 port map( D => n7042, CK => Clk, RN => n3911,
                           Q => pc_lut_15_1_port, QN => n2411);
   pc_lut_reg_15_0_inst : DFFR_X1 port map( D => n7041, CK => Clk, RN => n3912,
                           Q => pc_lut_15_0_port, QN => n2410);
   pc_lut_reg_26_4_inst : DFFR_X1 port map( D => n6687, CK => Clk, RN => n3912,
                           Q => pc_lut_26_4_port, QN => n2409);
   pc_lut_reg_26_3_inst : DFFR_X1 port map( D => n6691, CK => Clk, RN => n3912,
                           Q => pc_lut_26_3_port, QN => n2408);
   pc_lut_reg_26_1_inst : DFFR_X1 port map( D => n6690, CK => Clk, RN => n3912,
                           Q => pc_lut_26_1_port, QN => n2403);
   pc_lut_reg_28_4_inst : DFFR_X1 port map( D => n6623, CK => Clk, RN => n3912,
                           Q => n2402, QN => n1290);
   pc_lut_reg_28_3_inst : DFFR_X1 port map( D => n6627, CK => Clk, RN => n3912,
                           Q => n2398, QN => n1294);
   pc_lut_reg_28_2_inst : DFFR_X1 port map( D => n6624, CK => Clk, RN => n3912,
                           Q => n2396, QN => n1291);
   pc_lut_reg_29_4_inst : DFFR_X1 port map( D => n6591, CK => Clk, RN => n3912,
                           Q => n2395, QN => n1255);
   pc_lut_reg_29_3_inst : DFFR_X1 port map( D => n6595, CK => Clk, RN => n3912,
                           Q => n2393, QN => n1260);
   pc_lut_reg_29_2_inst : DFFR_X1 port map( D => n6592, CK => Clk, RN => n3912,
                           Q => n2390, QN => n1257);
   pc_lut_reg_29_0_inst : DFFR_X1 port map( D => n6593, CK => Clk, RN => n3912,
                           Q => n2388, QN => n1258);
   pc_target_reg_24_5_inst : DFFR_X1 port map( D => n5732, CK => Clk, RN => 
                           n3910, Q => n2387, QN => n302);
   pc_target_reg_24_4_inst : DFFR_X1 port map( D => n5727, CK => Clk, RN => 
                           n3911, Q => n2385, QN => n297);
   pc_target_reg_17_5_inst : DFFR_X1 port map( D => n5956, CK => Clk, RN => 
                           n3911, Q => n2373, QN => n544);
   pc_target_reg_17_4_inst : DFFR_X1 port map( D => n5951, CK => Clk, RN => 
                           n3911, Q => n2227, QN => n539);
   pc_target_reg_9_5_inst : DFFR_X1 port map( D => n6212, CK => Clk, RN => 
                           n3908, Q => n2226, QN => n821);
   pc_target_reg_9_4_inst : DFFR_X1 port map( D => n6207, CK => Clk, RN => 
                           n3908, Q => n2225, QN => n816);
   pc_target_reg_4_5_inst : DFFR_X1 port map( D => n6372, CK => Clk, RN => 
                           n3909, Q => n2224, QN => n992);
   pc_target_reg_4_4_inst : DFFR_X1 port map( D => n6367, CK => Clk, RN => 
                           n3909, Q => n2223, QN => n987);
   pc_target_reg_2_10_inst : DFFR_X1 port map( D => n6428, CK => Clk, RN => 
                           n3910, Q => pc_target_2_10_port, QN => n2193);
   pc_target_reg_2_9_inst : DFFR_X1 port map( D => n6438, CK => Clk, RN => 
                           n3910, Q => pc_target_2_9_port, QN => n2192);
   pc_target_reg_2_8_inst : DFFR_X1 port map( D => n6429, CK => Clk, RN => 
                           n3910, Q => pc_target_2_8_port, QN => n2190);
   pc_target_reg_10_10_inst : DFFR_X1 port map( D => n6172, CK => Clk, RN => 
                           n3908, Q => pc_target_10_10_port, QN => n2189);
   pc_target_reg_10_9_inst : DFFR_X1 port map( D => n6182, CK => Clk, RN => 
                           n3908, Q => pc_target_10_9_port, QN => n2146);
   pc_target_reg_10_8_inst : DFFR_X1 port map( D => n6173, CK => Clk, RN => 
                           n3908, Q => pc_target_10_8_port, QN => n2112);
   pc_target_reg_10_3_inst : DFFR_X1 port map( D => n6179, CK => Clk, RN => 
                           n3908, Q => pc_target_10_3_port, QN => n2095);
   pc_target_reg_15_10_inst : DFFR_X1 port map( D => n6012, CK => Clk, RN => 
                           n3909, Q => pc_target_15_10_port, QN => n2094);
   pc_target_reg_15_9_inst : DFFR_X1 port map( D => n6022, CK => Clk, RN => 
                           n3909, Q => pc_target_15_9_port, QN => n2093);
   pc_target_reg_15_8_inst : DFFR_X1 port map( D => n6013, CK => Clk, RN => 
                           n3909, Q => pc_target_15_8_port, QN => n2091);
   pc_target_reg_15_6_inst : DFFR_X1 port map( D => n6014, CK => Clk, RN => 
                           n3909, Q => pc_target_15_6_port, QN => n2061);
   pc_target_reg_15_5_inst : DFFR_X1 port map( D => n6020, CK => Clk, RN => 
                           n3909, Q => pc_target_15_5_port, QN => n2060);
   pc_target_reg_15_4_inst : DFFR_X1 port map( D => n6015, CK => Clk, RN => 
                           n3909, Q => pc_target_15_4_port, QN => n2057);
   pc_target_reg_15_2_inst : DFFR_X1 port map( D => n6016, CK => Clk, RN => 
                           n3909, Q => pc_target_15_2_port, QN => n2013);
   pc_target_reg_15_1_inst : DFFR_X1 port map( D => n6018, CK => Clk, RN => 
                           n3909, Q => pc_target_15_1_port, QN => n1962);
   pc_target_reg_15_0_inst : DFFR_X1 port map( D => n6017, CK => Clk, RN => 
                           n3912, Q => pc_target_15_0_port, QN => n1961);
   pc_target_reg_15_3_inst : DFFR_X1 port map( D => n6019, CK => Clk, RN => 
                           n3909, Q => pc_target_15_3_port, QN => n1960);
   pc_target_reg_2_3_inst : DFFR_X1 port map( D => n6435, CK => Clk, RN => 
                           n3910, Q => pc_target_2_3_port, QN => n1959);
   pc_target_reg_3_10_inst : DFFR_X1 port map( D => n6396, CK => Clk, RN => 
                           n3910, Q => pc_target_3_10_port, QN => n1928);
   pc_target_reg_3_9_inst : DFFR_X1 port map( D => n6406, CK => Clk, RN => 
                           n3909, Q => pc_target_3_9_port, QN => n1926);
   pc_target_reg_3_8_inst : DFFR_X1 port map( D => n6397, CK => Clk, RN => 
                           n3910, Q => pc_target_3_8_port, QN => n1925);
   pc_target_reg_3_6_inst : DFFR_X1 port map( D => n6398, CK => Clk, RN => 
                           n3910, Q => pc_target_3_6_port, QN => n1881);
   pc_target_reg_3_5_inst : DFFR_X1 port map( D => n6404, CK => Clk, RN => 
                           n3909, Q => pc_target_3_5_port, QN => n1827);
   pc_target_reg_3_4_inst : DFFR_X1 port map( D => n6399, CK => Clk, RN => 
                           n3910, Q => pc_target_3_4_port, QN => n1826);
   pc_target_reg_3_3_inst : DFFR_X1 port map( D => n6403, CK => Clk, RN => 
                           n3909, Q => pc_target_3_3_port, QN => n1824);
   pc_target_reg_3_2_inst : DFFR_X1 port map( D => n6400, CK => Clk, RN => 
                           n3910, Q => pc_target_3_2_port, QN => n1793);
   pc_target_reg_3_1_inst : DFFR_X1 port map( D => n6402, CK => Clk, RN => 
                           n3909, Q => pc_target_3_1_port, QN => n1790);
   pc_target_reg_3_0_inst : DFFR_X1 port map( D => n6401, CK => Clk, RN => 
                           n3921, Q => pc_target_3_0_port, QN => n1743);
   pc_target_reg_21_10_inst : DFFR_X1 port map( D => n5820, CK => Clk, RN => 
                           n3911, Q => pc_target_21_10_port, QN => n1709);
   pc_target_reg_21_9_inst : DFFR_X1 port map( D => n5830, CK => Clk, RN => 
                           n3911, Q => pc_target_21_9_port, QN => n1693);
   pc_target_reg_21_8_inst : DFFR_X1 port map( D => n5821, CK => Clk, RN => 
                           n3911, Q => pc_target_21_8_port, QN => n1692);
   pc_target_reg_21_6_inst : DFFR_X1 port map( D => n5822, CK => Clk, RN => 
                           n3911, Q => pc_target_21_6_port, QN => n1691);
   pc_target_reg_21_5_inst : DFFR_X1 port map( D => n5828, CK => Clk, RN => 
                           n3911, Q => pc_target_21_5_port, QN => n1690);
   pc_target_reg_21_4_inst : DFFR_X1 port map( D => n5823, CK => Clk, RN => 
                           n3911, Q => pc_target_21_4_port, QN => n1659);
   pc_target_reg_24_30_inst : DFFR_X1 port map( D => n5714, CK => Clk, RN => 
                           n3911, Q => n1658, QN => n284);
   U68 : NOR2_X1 port map( A1 => n2404, A2 => n2405, ZN => n2401);
   U69 : NOR2_X1 port map( A1 => n2412, A2 => n2413, ZN => n2400);
   U134 : INV_X1 port map( A => n2419, ZN => N215);
   U135 : OAI21_X1 port map( B1 => n1393, B2 => n2249, A => n2352, ZN => n2351)
                           ;
   U168 : NAND2_X1 port map( A1 => n2252, A2 => pc_lut_27_0_port, ZN => n2352);
   U169 : OAI21_X1 port map( B1 => n1258, B2 => n2254, A => n2353, ZN => n2350)
                           ;
   U202 : NAND2_X1 port map( A1 => n2257, A2 => pc_lut_31_0_port, ZN => n2353);
   U203 : OAI21_X1 port map( B1 => n1657, B2 => n2259, A => n2354, ZN => n2349)
                           ;
   U204 : NAND2_X1 port map( A1 => n2262, A2 => pc_lut_19_0_port, ZN => n2354);
   U269 : OAI21_X1 port map( B1 => n1461, B2 => n2264, A => n2355, ZN => n2348)
                           ;
   U270 : NAND2_X1 port map( A1 => n2267, A2 => pc_lut_21_0_port, ZN => n2355);
   U335 : OAI21_X1 port map( B1 => n1927, B2 => n2273, A => n2360, ZN => n2359)
                           ;
   U336 : NAND2_X1 port map( A1 => n2276, A2 => pc_lut_11_0_port, ZN => n2360);
   U369 : OAI21_X1 port map( B1 => n1792, B2 => n2278, A => n2361, ZN => n2358)
                           ;
   U370 : NAND2_X1 port map( A1 => n2281, A2 => pc_lut_15_0_port, ZN => n2361);
   U403 : OAI21_X1 port map( B1 => n2191, B2 => n2283, A => n2362, ZN => n2357)
                           ;
   U404 : NAND2_X1 port map( A1 => n2286, A2 => pc_lut_3_0_port, ZN => n2362);
   U405 : OAI21_X1 port map( B1 => n2059, B2 => n2288, A => n2363, ZN => n2356)
                           ;
   U438 : NAND2_X1 port map( A1 => n2291, A2 => pc_lut_7_0_port, ZN => n2363);
   U439 : INV_X1 port map( A => n2370, ZN => n2369);
   U472 : INV_X1 port map( A => n2371, ZN => n2368);
   U473 : INV_X1 port map( A => n2372, ZN => n2367);
   U538 : OAI22_X1 port map( A1 => n1497, A2 => n2263, B1 => n1462, B2 => n2264
                           , ZN => n2366);
   U539 : INV_X1 port map( A => n2378, ZN => n2377);
   U604 : INV_X1 port map( A => n2379, ZN => n2376);
   U605 : INV_X1 port map( A => n2380, ZN => n2375);
   U606 : INV_X1 port map( A => n2381, ZN => n2374);
   U671 : NOR2_X1 port map( A1 => n2384, A2 => n2386, ZN => n2383);
   U672 : NOR2_X1 port map( A1 => n2392, A2 => n2394, ZN => n2382);
   U737 : INV_X2 port map( A => Set_target(15), ZN => n123_port);
   U738 : INV_X2 port map( A => Set_target(13), ZN => n121_port);
   U771 : INV_X2 port map( A => Set_target(12), ZN => n95);
   U772 : INV_X2 port map( A => Set_target(14), ZN => n93);
   U777 : INV_X2 port map( A => n2210, ZN => n2208);
   U805 : NAND2_X4 port map( A1 => n2141, A2 => n176, ZN => n2210);
   U806 : INV_X2 port map( A => n1946, ZN => n1944);
   U808 : INV_X2 port map( A => n1676, ZN => n1674);
   U873 : INV_X2 port map( A => n2078, ZN => n2076);
   U874 : INV_X2 port map( A => n2176, ZN => n2174);
   U939 : NAND2_X4 port map( A1 => n2141, A2 => n141, ZN => n2176);
   U940 : AND2_X1 port map( A1 => n2141, A2 => n74, ZN => n2);
   U973 : INV_X1 port map( A => n2, ZN => n3);
   U974 : INV_X1 port map( A => n2, ZN => n283);
   U1007 : NAND2_X4 port map( A1 => n2010, A2 => n141, ZN => n2044);
   U1008 : NAND2_X4 port map( A1 => n1608, A2 => n141, ZN => n1642);
   U1009 : NAND2_X4 port map( A1 => n1878, A2 => n141, ZN => n1912);
   U1074 : NAND2_X4 port map( A1 => n2010, A2 => n176, ZN => n2078);
   U1075 : NAND2_X4 port map( A1 => n1878, A2 => n176, ZN => n1946);
   U1140 : NAND2_X4 port map( A1 => n1608, A2 => n176, ZN => n1676);
   U1174 : NAND2_X4 port map( A1 => n1742, A2 => n176, ZN => n1811);
   U1175 : NOR2_X4 port map( A1 => PC_write(0), A2 => PC_write(1), ZN => n176);
   U1209 : AND2_X1 port map( A1 => n1608, A2 => n74, ZN => n525);
   U1210 : INV_X1 port map( A => n525, ZN => n558);
   U1275 : INV_X1 port map( A => n525, ZN => n768);
   U1276 : AND2_X1 port map( A1 => n2141, A2 => n38, ZN => n802);
   U1341 : INV_X1 port map( A => n802, ZN => n871);
   U1342 : INV_X1 port map( A => n802, ZN => n973);
   U1375 : AND2_X1 port map( A1 => n1878, A2 => n74, ZN => n1240);
   U1376 : INV_X1 port map( A => n1240, ZN => n1256);
   U1409 : INV_X1 port map( A => n1240, ZN => n1259);
   U1410 : AND2_X1 port map( A1 => n2010, A2 => n74, ZN => n1275);
   U1411 : INV_X1 port map( A => n1275, ZN => n1292);
   U1476 : INV_X1 port map( A => n1275, ZN => n1293);
   U1543 : NAND2_X4 port map( A1 => n1742, A2 => n141, ZN => n1777);
   U1576 : AND2_X1 port map( A1 => n1478, A2 => n74, ZN => n1344);
   U1577 : INV_X1 port map( A => n1344, ZN => n1392);
   U1579 : INV_X1 port map( A => n1344, ZN => n1394);
   U1591 : INV_X2 port map( A => n697, ZN => n698);
   U1593 : NAND2_X2 port map( A1 => n628, A2 => n176, ZN => n697);
   U1595 : INV_X2 port map( A => n1109, ZN => n1110);
   U1621 : INV_X2 port map( A => n1075, ZN => n1076);
   U1623 : INV_X2 port map( A => n317, ZN => n318);
   U1625 : INV_X2 port map( A => n352, ZN => n353);
   U1627 : INV_X2 port map( A => n76, ZN => n77);
   U1629 : NOR2_X4 port map( A1 => n2143, A2 => PC_write(1), ZN => n141);
   U1631 : INV_X2 port map( A => n663, ZN => n664);
   U1633 : NOR2_X4 port map( A1 => n2142, A2 => n2143, ZN => n38);
   U1635 : INV_X2 port map( A => n631, ZN => n630);
   U1637 : NAND2_X2 port map( A1 => PC_write(23), A2 => n3521, ZN => n1197);
   U1639 : NAND2_X2 port map( A1 => PC_write(25), A2 => n3521, ZN => n1199);
   U1641 : NAND2_X2 port map( A1 => PC_write(27), A2 => n3521, ZN => n1201);
   U1642 : NAND2_X2 port map( A1 => PC_write(21), A2 => n3521, ZN => n1195);
   U1643 : NAND2_X2 port map( A1 => PC_write(19), A2 => n3521, ZN => n1193);
   U1644 : NAND2_X2 port map( A1 => PC_write(29), A2 => n3521, ZN => n1203);
   U1645 : NAND2_X2 port map( A1 => PC_write(31), A2 => n3521, ZN => n1205);
   U1648 : NAND2_X2 port map( A1 => PC_write(17), A2 => n3521, ZN => n1191);
   U1650 : NAND2_X2 port map( A1 => PC_write(15), A2 => n3521, ZN => n1189);
   U1652 : NAND2_X2 port map( A1 => PC_write(28), A2 => n3521, ZN => n1150);
   U1654 : NAND2_X2 port map( A1 => PC_write(26), A2 => n3521, ZN => n1152);
   U1656 : NAND2_X2 port map( A1 => PC_write(13), A2 => n3521, ZN => n1187);
   U1658 : NAND2_X2 port map( A1 => PC_write(11), A2 => n3521, ZN => n1185);
   U1660 : NAND2_X2 port map( A1 => PC_write(24), A2 => n3521, ZN => n1154);
   U1662 : NAND2_X2 port map( A1 => PC_write(22), A2 => n3521, ZN => n1156);
   U1664 : NAND2_X2 port map( A1 => PC_write(9), A2 => n3521, ZN => n1183);
   U1666 : NAND2_X2 port map( A1 => PC_write(7), A2 => n3521, ZN => n1181);
   U1668 : NAND2_X2 port map( A1 => PC_write(20), A2 => n3521, ZN => n1158);
   U1670 : NAND2_X2 port map( A1 => PC_write(18), A2 => n3521, ZN => n1160);
   U1672 : NAND2_X2 port map( A1 => PC_write(5), A2 => n3521, ZN => n1179);
   U1684 : NAND2_X2 port map( A1 => PC_write(6), A2 => n3521, ZN => n1172);
   U1686 : NAND2_X2 port map( A1 => PC_write(16), A2 => n3521, ZN => n1162);
   U1688 : NAND2_X2 port map( A1 => PC_write(14), A2 => n3521, ZN => n1164);
   U1690 : NAND2_X2 port map( A1 => PC_write(8), A2 => n3521, ZN => n1170);
   U1692 : NAND2_X2 port map( A1 => PC_write(10), A2 => n3521, ZN => n1168);
   U1694 : NAND2_X2 port map( A1 => PC_write(12), A2 => n3521, ZN => n1166);
   U1696 : NAND2_X2 port map( A1 => PC_write(30), A2 => n3521, ZN => n1147);
   U1698 : AND2_X1 port map( A1 => n1478, A2 => n38, ZN => n1426);
   U1700 : INV_X1 port map( A => n1426, ZN => n1427);
   U1702 : INV_X1 port map( A => n1426, ZN => n1428);
   U1706 : NOR2_X4 port map( A1 => n2142, A2 => PC_write(0), ZN => n74);
   U1710 : AND2_X2 port map( A1 => n316, A2 => n177, ZN => n213_port);
   U1712 : AND2_X1 port map( A1 => n489, A2 => n176, ZN => n1446);
   U1714 : INV_X1 port map( A => n1446, ZN => n1463);
   U1716 : INV_X1 port map( A => n1446, ZN => n1481);
   U1720 : INV_X1 port map( A => n3521, ZN => n1496);
   U1722 : BUF_X8 port map( A => n3518, Z => n3521);
   U1724 : INV_X2 port map( A => n906, ZN => n905);
   U1728 : AND2_X1 port map( A1 => n903, A2 => n38, ZN => n1498);
   U1730 : INV_X1 port map( A => n1498, ZN => n1611);
   U1732 : INV_X1 port map( A => n1498, ZN => n1656);
   U1734 : INV_X2 port map( A => n734, ZN => n733);
   U1738 : INV_X2 port map( A => n248, ZN => n249);
   U1749 : INV_X2 port map( A => n835, ZN => n836);
   U1751 : NAND2_X2 port map( A1 => n766, A2 => n176, ZN => n835);
   U1755 : AND2_X2 port map( A1 => n731, A2 => n454, ZN => n903);
   U1757 : AND2_X4 port map( A1 => n3437, A2 => n3420, ZN => n2291);
   U1759 : AND2_X4 port map( A1 => n3415, A2 => n3416, ZN => n2252);
   U1761 : AND2_X4 port map( A1 => n3415, A2 => n3420, ZN => n2257);
   U1763 : AND2_X4 port map( A1 => n3421, A2 => n3424, ZN => n2267);
   U1765 : AND2_X4 port map( A1 => n3433, A2 => n3416, ZN => n2276);
   U1767 : NOR3_X2 port map( A1 => n3422, A2 => PC_read(4), A3 => n3427, ZN => 
                           n3433);
   U1769 : AND2_X4 port map( A1 => n3437, A2 => n3416, ZN => n2286);
   U1771 : NOR2_X2 port map( A1 => n3439, A2 => PC_read(2), ZN => n3416);
   U1773 : NOR3_X2 port map( A1 => PC_read(3), A2 => PC_read(4), A3 => n3422, 
                           ZN => n3437);
   U1775 : AND2_X4 port map( A1 => n3433, A2 => n3420, ZN => n2281);
   U1776 : AND2_X4 port map( A1 => n3416, A2 => n3424, ZN => n2262);
   U1777 : NAND2_X4 port map( A1 => n3415, A2 => n3421, ZN => n2254);
   U1794 : NAND2_X4 port map( A1 => n3424, A2 => n3420, ZN => n2264);
   U1810 : NOR2_X2 port map( A1 => n3441, A2 => n3439, ZN => n3420);
   U1811 : NAND2_X4 port map( A1 => n3433, A2 => n3418, ZN => n2273);
   U1827 : NAND2_X4 port map( A1 => n3437, A2 => n3418, ZN => n2283);
   U1828 : NAND2_X4 port map( A1 => n3415, A2 => n3418, ZN => n2249);
   U1844 : NAND2_X4 port map( A1 => n3437, A2 => n3421, ZN => n2288);
   U1845 : NAND2_X4 port map( A1 => n3433, A2 => n3421, ZN => n2278);
   U1848 : NAND2_X4 port map( A1 => n3418, A2 => n3424, ZN => n2259);
   U1850 : NAND2_X4 port map( A1 => n3434, A2 => n3418, ZN => n2272);
   U1852 : NOR2_X2 port map( A1 => PC_read(1), A2 => PC_read(2), ZN => n3418);
   U1854 : NOR3_X2 port map( A1 => PC_read(0), A2 => PC_read(4), A3 => n3427, 
                           ZN => n3434);
   U1856 : NAND2_X4 port map( A1 => n3417, A2 => n3421, ZN => n2253);
   U1858 : NAND2_X4 port map( A1 => n3420, A2 => n3425, ZN => n2263);
   U1860 : NAND2_X4 port map( A1 => n3438, A2 => n3418, ZN => n2282);
   U1862 : NOR3_X2 port map( A1 => PC_read(3), A2 => PC_read(4), A3 => 
                           PC_read(0), ZN => n3438);
   U1864 : NAND2_X4 port map( A1 => n3418, A2 => n3425, ZN => n2258);
   U1866 : NAND2_X4 port map( A1 => n3434, A2 => n3421, ZN => n2277);
   U1868 : NAND2_X4 port map( A1 => n3438, A2 => n3421, ZN => n2287);
   U1870 : NOR2_X2 port map( A1 => n3441, A2 => PC_read(1), ZN => n3421);
   U1872 : NAND2_X4 port map( A1 => n3417, A2 => n3418, ZN => n2248);
   U1875 : AND2_X4 port map( A1 => n3421, A2 => n3425, ZN => n2266);
   U1883 : AND2_X4 port map( A1 => n3434, A2 => n3416, ZN => n2275);
   U1885 : AND2_X4 port map( A1 => n3416, A2 => n3425, ZN => n2261);
   U1887 : AND2_X4 port map( A1 => n3434, A2 => n3420, ZN => n2280);
   U1889 : AND2_X4 port map( A1 => n3417, A2 => n3420, ZN => n2256);
   U1891 : AND2_X4 port map( A1 => n3438, A2 => n3420, ZN => n2290);
   U1893 : AND2_X4 port map( A1 => n3438, A2 => n3416, ZN => n2285);
   U1895 : AND2_X4 port map( A1 => n3417, A2 => n3416, ZN => n2251);
   U1897 : NAND2_X4 port map( A1 => n628, A2 => n141, ZN => n663);
   U1901 : AND2_X4 port map( A1 => n766, A2 => n141, ZN => n3442);
   U1903 : INV_X4 port map( A => n3442, ZN => n801);
   U1905 : NAND2_X4 port map( A1 => n1040, A2 => n141, ZN => n1075);
   U1909 : AND2_X4 port map( A1 => n731, A2 => n592, ZN => n1040);
   U1910 : AND2_X4 port map( A1 => n903, A2 => n176, ZN => n3443);
   U1911 : INV_X4 port map( A => n3443, ZN => n972);
   U1940 : INV_X2 port map( A => Set_target(22), ZN => n85);
   U1974 : INV_X2 port map( A => Set_target(17), ZN => n125_port);
   U1975 : INV_X2 port map( A => Set_target(16), ZN => n91);
   U1990 : INV_X2 port map( A => Set_target(18), ZN => n89);
   U1992 : NAND2_X4 port map( A1 => n141, A2 => n39, ZN => n76);
   U2009 : AND2_X4 port map( A1 => n177, A2 => n178, ZN => n39);
   U2024 : AND2_X4 port map( A1 => n213_port, A2 => n176, ZN => n3444);
   U2025 : INV_X4 port map( A => n3444, ZN => n282);
   U2026 : NAND2_X4 port map( A1 => n351, A2 => n74, ZN => n352);
   U2042 : NAND2_X4 port map( A1 => n351, A2 => n38, ZN => n317);
   U2077 : AND2_X4 port map( A1 => n489, A2 => n141, ZN => n3445);
   U2078 : INV_X4 port map( A => n3445, ZN => n524);
   U2094 : AND2_X4 port map( A1 => n766, A2 => n74, ZN => n3446);
   U2096 : INV_X4 port map( A => n3446, ZN => n769);
   U2111 : OR2_X4 port map( A1 => n3447, A2 => n3448, ZN => n631);
   U2112 : INV_X1 port map( A => n628, ZN => n3447);
   U2114 : INV_X1 port map( A => n74, ZN => n3448);
   U2116 : MUX2_X1 port map( A => Set_target(22), B => pc_target_16_22_port, S 
                           => n1463, Z => n5974);
   U2118 : INV_X2 port map( A => n1043, ZN => n1042);
   U2120 : NAND2_X4 port map( A1 => n1040, A2 => n74, ZN => n1043);
   U2122 : INV_X2 port map( A => Set_target(30), ZN => n75);
   U2158 : INV_X2 port map( A => Set_target(11), ZN => n119_port);
   U2160 : CLKBUF_X1 port map( A => SetT_NT, Z => n3518);
   U2162 : INV_X2 port map( A => Set_target(21), ZN => n129);
   U2164 : INV_X2 port map( A => Set_target(25), ZN => n133);
   U2166 : INV_X2 port map( A => Set_target(24), ZN => n83);
   U2168 : INV_X2 port map( A => Set_target(26), ZN => n81);
   U2170 : INV_X2 port map( A => Set_target(29), ZN => n137);
   U2172 : AND2_X2 port map( A1 => n3519, A2 => n316, ZN => n766);
   U2174 : AND2_X1 port map( A1 => n3520, A2 => n1143, ZN => n3519);
   U2175 : AND2_X1 port map( A1 => n3520, A2 => n1143, ZN => n731);
   U2180 : INV_X2 port map( A => n422, ZN => n421);
   U2186 : AND4_X1 port map( A1 => WR, A2 => SetT_NT, A3 => Enable, A4 => n1144
                           , ZN => n593);
   U2188 : AND2_X2 port map( A1 => n3519, A2 => n178, ZN => n628);
   U2192 : INV_X4 port map( A => n1611, ZN => n870);
   U2196 : AND2_X2 port map( A1 => n593, A2 => PC_write(4), ZN => n177);
   U2198 : INV_X2 port map( A => Set_target(19), ZN => n127_port);
   U2200 : INV_X1 port map( A => n3518, ZN => n3529);
   U2202 : INV_X2 port map( A => Set_target(23), ZN => n131);
   U2207 : INV_X2 port map( A => Set_target(20), ZN => n87);
   U2208 : INV_X2 port map( A => Set_target(28), ZN => n79);
   U2209 : INV_X2 port map( A => Set_target(27), ZN => n135);
   U2211 : INV_X1 port map( A => n1980, ZN => n3522);
   U2213 : INV_X1 port map( A => n3522, ZN => n3523);
   U2215 : INV_X2 port map( A => n3522, ZN => n3524);
   U2217 : INV_X1 port map( A => n1848, ZN => n3525);
   U2219 : INV_X1 port map( A => n3525, ZN => n3526);
   U2221 : INV_X2 port map( A => n3525, ZN => n3527);
   U2223 : INV_X2 port map( A => n1463, ZN => n559);
   U2227 : INV_X2 port map( A => n216_port, ZN => n215_port);
   U2229 : INV_X2 port map( A => n457, ZN => n456);
   U2233 : INV_X2 port map( A => n6, ZN => n5);
   U2237 : INV_X1 port map( A => SetT_NT, ZN => n3528);
   U2238 : INV_X1 port map( A => n1578, ZN => n3530);
   U2239 : INV_X1 port map( A => n3530, ZN => n3531);
   U2269 : INV_X1 port map( A => n3530, ZN => n3533);
   U2274 : INV_X1 port map( A => n3530, ZN => n3532);
   U2303 : AND2_X4 port map( A1 => n1206, A2 => n176, ZN => n3534);
   U2306 : INV_X4 port map( A => n3534, ZN => n1277);
   U2308 : AND2_X4 port map( A1 => n1742, A2 => n74, ZN => n3535);
   U2310 : INV_X4 port map( A => n3535, ZN => n1745);
   U2312 : AND2_X4 port map( A1 => n1206, A2 => n141, ZN => n3536);
   U2314 : INV_X4 port map( A => n3536, ZN => n1242);
   U2316 : AND2_X4 port map( A1 => n1742, A2 => n38, ZN => n3537);
   U2318 : INV_X4 port map( A => n3537, ZN => n1711);
   U2320 : AND2_X4 port map( A1 => n1343, A2 => n74, ZN => n3538);
   U2324 : INV_X2 port map( A => n2044, ZN => n2042);
   U2326 : INV_X2 port map( A => n1912, ZN => n1910);
   U2328 : INV_X2 port map( A => n1811, ZN => n1809);
   U2330 : INV_X2 port map( A => n1642, ZN => n1640);
   U2333 : INV_X2 port map( A => n1777, ZN => n1775);
   U2334 : INV_X2 port map( A => n1412, ZN => n1410);
   U2337 : INV_X2 port map( A => n1392, ZN => n1479);
   U2339 : INV_X2 port map( A => n3, ZN => n2144);
   U2341 : INV_X2 port map( A => n1378, ZN => n1376);
   U2343 : INV_X2 port map( A => n1427, ZN => n1444);
   U2347 : INV_X2 port map( A => n1292, ZN => n2011);
   U2349 : INV_X2 port map( A => n1256, ZN => n1879);
   U2351 : INV_X2 port map( A => n558, ZN => n1609);
   U2353 : INV_X2 port map( A => n871, ZN => n2110);
   U2357 : INV_X2 port map( A => n3523, ZN => n1978);
   U2359 : INV_X2 port map( A => n3526, ZN => n1846);
   U2361 : INV_X2 port map( A => n3531, ZN => n1576);
   eq_43 : BTB_PC_SIZE32_BTBSIZE5_DW01_cmp6_0 port map( A(31) => N188, A(30) =>
                           N189, A(29) => N190, A(28) => N191, A(27) => N192, 
                           A(26) => N193, A(25) => N194, A(24) => N195, A(23) 
                           => N196, A(22) => N197, A(21) => N198, A(20) => N199
                           , A(19) => N200, A(18) => N201, A(17) => N202, A(16)
                           => N203, A(15) => N204, A(14) => N205, A(13) => N206
                           , A(12) => N207, A(11) => N208, A(10) => N209, A(9) 
                           => N210, A(8) => N211, A(7) => N212, A(6) => N213, 
                           A(5) => N214, A(4) => N215, A(3) => N216, A(2) => 
                           N217, A(1) => N218, A(0) => N219, B(31) => 
                           PC_read(31), B(30) => PC_read(30), B(29) => 
                           PC_read(29), B(28) => PC_read(28), B(27) => 
                           PC_read(27), B(26) => PC_read(26), B(25) => 
                           PC_read(25), B(24) => PC_read(24), B(23) => 
                           PC_read(23), B(22) => PC_read(22), B(21) => 
                           PC_read(21), B(20) => PC_read(20), B(19) => 
                           PC_read(19), B(18) => PC_read(18), B(17) => 
                           PC_read(17), B(16) => PC_read(16), B(15) => 
                           PC_read(15), B(14) => PC_read(14), B(13) => 
                           PC_read(13), B(12) => PC_read(12), B(11) => 
                           PC_read(11), B(10) => PC_read(10), B(9) => 
                           PC_read(9), B(8) => PC_read(8), B(7) => PC_read(7), 
                           B(6) => PC_read(6), B(5) => PC_read(5), B(4) => 
                           PC_read(4), B(3) => PC_read(3), B(2) => PC_read(2), 
                           B(1) => PC_read(1), B(0) => PC_read(0), TC => n1, LT
                           => n_1112, GT => n_1113, EQ => N220, LE => n_1114, 
                           GE => n_1115, NE => n_1116);
   pc_target_reg_16_30_inst : DFFR_X1 port map( D => n5970, CK => Clk, RN => 
                           Reset, Q => n3792, QN => n560);
   pc_target_reg_9_30_inst : DFFR_X1 port map( D => n6194, CK => Clk, RN => 
                           Reset, Q => n3791, QN => n803);
   pc_target_reg_4_30_inst : DFFR_X1 port map( D => n6354, CK => Clk, RN => 
                           Reset, Q => n3790, QN => n974);
   pc_target_reg_17_30_inst : DFFR_X1 port map( D => n5938, CK => Clk, RN => 
                           Reset, Q => n3789, QN => n526);
   pc_target_reg_13_30_inst : DFFR_X1 port map( D => n6066, CK => Clk, RN => 
                           Reset, Q => n3788, QN => n665);
   pc_target_reg_5_30_inst : DFFR_X1 port map( D => n6322, CK => Clk, RN => 
                           Reset, Q => n3787, QN => n940);
   pc_target_reg_0_30_inst : DFFR_X1 port map( D => n6482, CK => Clk, RN => 
                           Reset, Q => n3786, QN => n1111);
   pc_target_reg_1_30_inst : DFFR_X1 port map( D => n6450, CK => Clk, RN => 
                           Reset, Q => n3785, QN => n1077);
   pc_target_reg_23_30_inst : DFFR_X1 port map( D => n5746, CK => Clk, RN => 
                           Reset, Q => n3784, QN => n319);
   pc_target_reg_22_30_inst : DFFR_X1 port map( D => n5778, CK => Clk, RN => 
                           Reset, Q => n3783, QN => n354);
   pc_target_reg_25_30_inst : DFFR_X1 port map( D => n5682, CK => Clk, RN => 
                           Reset, Q => n3782, QN => n250);
   pc_target_reg_28_30_inst : DFFR_X1 port map( D => n5586, CK => Clk, RN => 
                           Reset, Q => n3781, QN => n144);
   pc_target_reg_29_30_inst : DFFR_X1 port map( D => n5554, CK => Clk, RN => 
                           Reset, Q => n3780, QN => n78);
   pc_target_reg_8_30_inst : DFFR_X1 port map( D => n6226, CK => Clk, RN => 
                           Reset, Q => n3779, QN => n837);
   pc_target_reg_12_30_inst : DFFR_X1 port map( D => n6098, CK => Clk, RN => 
                           Reset, Q => n3778, QN => n699);
   pc_target_reg_16_22_inst : DFFR_X1 port map( D => n5974, CK => Clk, RN => 
                           Reset, Q => pc_target_16_22_port, QN => n564);
   pc_lut_reg_31_3_inst : DFFR_X1 port map( D => n6531, CK => Clk, RN => Reset,
                           Q => pc_lut_31_3_port, QN => n3777);
   pc_lut_reg_31_2_inst : DFFR_X1 port map( D => n6528, CK => Clk, RN => Reset,
                           Q => pc_lut_31_2_port, QN => n3776);
   pc_lut_reg_31_1_inst : DFFR_X1 port map( D => n6530, CK => Clk, RN => Reset,
                           Q => pc_lut_31_1_port, QN => n3775);
   pc_lut_reg_31_0_inst : DFFR_X1 port map( D => n6529, CK => Clk, RN => Reset,
                           Q => pc_lut_31_0_port, QN => n3774);
   pc_lut_reg_27_3_inst : DFFR_X1 port map( D => n6659, CK => Clk, RN => Reset,
                           Q => pc_lut_27_3_port, QN => n3773);
   pc_lut_reg_27_1_inst : DFFR_X1 port map( D => n6658, CK => Clk, RN => Reset,
                           Q => pc_lut_27_1_port, QN => n3772);
   pc_lut_reg_27_0_inst : DFFR_X1 port map( D => n6657, CK => Clk, RN => Reset,
                           Q => pc_lut_27_0_port, QN => n3771);
   pc_lut_reg_31_4_inst : DFFR_X1 port map( D => n6527, CK => Clk, RN => Reset,
                           Q => pc_lut_31_4_port, QN => n3770);
   pc_lut_reg_27_4_inst : DFFR_X1 port map( D => n6655, CK => Clk, RN => Reset,
                           Q => pc_lut_27_4_port, QN => n3769);
   pc_target_reg_7_31_inst : DFFR_X1 port map( D => n6289, CK => Clk, RN => 
                           Reset, Q => pc_target_7_31_port, QN => n3768);
   pc_target_reg_7_23_inst : DFFR_X1 port map( D => n6285, CK => Clk, RN => 
                           Reset, Q => pc_target_7_23_port, QN => n3767);
   pc_target_reg_7_26_inst : DFFR_X1 port map( D => n6260, CK => Clk, RN => 
                           Reset, Q => pc_target_7_26_port, QN => n3766);
   pc_target_reg_7_19_inst : DFFR_X1 port map( D => n6283, CK => Clk, RN => 
                           Reset, Q => pc_target_7_19_port, QN => n3765);
   pc_target_reg_7_14_inst : DFFR_X1 port map( D => n6266, CK => Clk, RN => 
                           Reset, Q => pc_target_7_14_port, QN => n3764);
   pc_target_reg_7_11_inst : DFFR_X1 port map( D => n6279, CK => Clk, RN => 
                           Reset, Q => pc_target_7_11_port, QN => n3763);
   pc_target_reg_7_30_inst : DFFR_X1 port map( D => n6258, CK => Clk, RN => 
                           Reset, Q => pc_target_7_30_port, QN => n3762);
   pc_target_reg_7_29_inst : DFFR_X1 port map( D => n6288, CK => Clk, RN => 
                           Reset, Q => pc_target_7_29_port, QN => n3761);
   pc_target_reg_7_28_inst : DFFR_X1 port map( D => n6259, CK => Clk, RN => 
                           Reset, Q => pc_target_7_28_port, QN => n3760);
   pc_target_reg_7_27_inst : DFFR_X1 port map( D => n6287, CK => Clk, RN => 
                           Reset, Q => pc_target_7_27_port, QN => n3759);
   pc_target_reg_7_25_inst : DFFR_X1 port map( D => n6286, CK => Clk, RN => 
                           Reset, Q => pc_target_7_25_port, QN => n3758);
   pc_target_reg_7_24_inst : DFFR_X1 port map( D => n6261, CK => Clk, RN => 
                           Reset, Q => pc_target_7_24_port, QN => n3757);
   pc_target_reg_7_22_inst : DFFR_X1 port map( D => n6262, CK => Clk, RN => 
                           Reset, Q => pc_target_7_22_port, QN => n3756);
   pc_target_reg_7_21_inst : DFFR_X1 port map( D => n6284, CK => Clk, RN => 
                           Reset, Q => pc_target_7_21_port, QN => n3755);
   pc_target_reg_7_20_inst : DFFR_X1 port map( D => n6263, CK => Clk, RN => 
                           Reset, Q => pc_target_7_20_port, QN => n3754);
   pc_target_reg_7_18_inst : DFFR_X1 port map( D => n6264, CK => Clk, RN => 
                           Reset, Q => pc_target_7_18_port, QN => n3753);
   pc_target_reg_7_17_inst : DFFR_X1 port map( D => n6282, CK => Clk, RN => 
                           Reset, Q => pc_target_7_17_port, QN => n3752);
   pc_target_reg_7_16_inst : DFFR_X1 port map( D => n6265, CK => Clk, RN => 
                           Reset, Q => pc_target_7_16_port, QN => n3751);
   pc_target_reg_7_15_inst : DFFR_X1 port map( D => n6281, CK => Clk, RN => 
                           Reset, Q => pc_target_7_15_port, QN => n3750);
   pc_target_reg_7_13_inst : DFFR_X1 port map( D => n6280, CK => Clk, RN => 
                           Reset, Q => pc_target_7_13_port, QN => n3749);
   pc_target_reg_7_12_inst : DFFR_X1 port map( D => n6267, CK => Clk, RN => 
                           Reset, Q => pc_target_7_12_port, QN => n3748);
   pc_target_reg_7_10_inst : DFFR_X1 port map( D => n6268, CK => Clk, RN => 
                           Reset, Q => pc_target_7_10_port, QN => n3747);
   pc_target_reg_7_9_inst : DFFR_X1 port map( D => n6278, CK => Clk, RN => 
                           Reset, Q => pc_target_7_9_port, QN => n3746);
   pc_target_reg_7_8_inst : DFFR_X1 port map( D => n6269, CK => Clk, RN => 
                           Reset, Q => pc_target_7_8_port, QN => n3745);
   pc_target_reg_7_7_inst : DFFR_X1 port map( D => n6277, CK => Clk, RN => 
                           Reset, Q => pc_target_7_7_port, QN => n3744);
   U807 : INV_X2 port map( A => n938, ZN => n939);
   U1141 : NAND2_X4 port map( A1 => n903, A2 => n141, ZN => n938);
   U1208 : INV_X2 port map( A => n3810, ZN => n1515);
   U1477 : NAND2_X4 port map( A1 => n1040, A2 => n176, ZN => n1109);
   U1542 : NAND2_X4 port map( A1 => n766, A2 => n38, ZN => n734);
   U1581 : OAI211_X1 port map( C1 => n3528, C2 => n1144, A => Enable, B => WR, 
                           ZN => n3793);
   U1583 : NOR2_X1 port map( A1 => n1708, A2 => PC_write(4), ZN => n3794);
   U1585 : NAND2_X4 port map( A1 => n903, A2 => n74, ZN => n906);
   U1587 : NAND2_X4 port map( A1 => n213_port, A2 => n141, ZN => n248);
   U1589 : INV_X2 port map( A => n3538, ZN => n1346);
   U1597 : INV_X2 port map( A => n596, ZN => n595);
   U1704 : NAND2_X4 port map( A1 => n628, A2 => n38, ZN => n596);
   U1708 : AND2_X1 port map( A1 => n1206, A2 => n38, ZN => n3795);
   U1711 : INV_X4 port map( A => n3795, ZN => n1148);
   U1718 : AND4_X1 port map( A1 => WR, A2 => SetT_NT, A3 => Enable, A4 => n1144
                           , ZN => n3520);
   U1726 : INV_X2 port map( A => n3805, ZN => n1209);
   U1736 : AND2_X2 port map( A1 => n1309, A2 => n592, ZN => n1608);
   U1743 : AND2_X1 port map( A1 => n1343, A2 => n38, ZN => n3796);
   U1753 : INV_X4 port map( A => n3796, ZN => n1312);
   U1846 : INV_X2 port map( A => n1008, ZN => n1007);
   U1899 : NAND2_X4 port map( A1 => n1040, A2 => n38, ZN => n1008);
   U1907 : INV_X2 port map( A => n142, ZN => n143);
   U1913 : NAND2_X4 port map( A1 => n176, A2 => n39, ZN => n142);
   U1915 : NAND2_X4 port map( A1 => n213_port, A2 => n74, ZN => n216_port);
   U1917 : AND2_X4 port map( A1 => n213_port, A2 => n38, ZN => n3797);
   U1919 : INV_X4 port map( A => n3797, ZN => n181);
   U1921 : NAND2_X4 port map( A1 => n489, A2 => n38, ZN => n457);
   U1923 : NAND2_X4 port map( A1 => n38, A2 => n39, ZN => n6);
   U1925 : AND2_X4 port map( A1 => n74, A2 => n39, ZN => n3798);
   U1927 : INV_X4 port map( A => n3798, ZN => n42);
   U1929 : NAND2_X4 port map( A1 => n351, A2 => n176, ZN => n422);
   U1931 : AND2_X4 port map( A1 => n454, A2 => n177, ZN => n351);
   U1933 : NAND2_X4 port map( A1 => n1343, A2 => n176, ZN => n1412);
   U1935 : AND2_X4 port map( A1 => n351, A2 => n141, ZN => n3799);
   U1937 : INV_X4 port map( A => n3799, ZN => n388);
   U1941 : INV_X2 port map( A => n492, ZN => n491);
   U1947 : NAND2_X4 port map( A1 => n489, A2 => n74, ZN => n492);
   U1949 : AND2_X2 port map( A1 => n592, A2 => n177, ZN => n489);
   U1951 : AND2_X4 port map( A1 => n1478, A2 => n176, ZN => n3800);
   U1953 : INV_X4 port map( A => n3800, ZN => n1547);
   U1955 : AND2_X2 port map( A1 => n1843, A2 => n178, ZN => n1742);
   U1957 : INV_X1 port map( A => n3796, ZN => n3801);
   U1959 : INV_X1 port map( A => n3801, ZN => n3802);
   U1961 : INV_X2 port map( A => n3801, ZN => n3804);
   U1963 : INV_X2 port map( A => n3801, ZN => n3803);
   U1965 : AND2_X4 port map( A1 => n1206, A2 => n74, ZN => n3805);
   U1967 : INV_X1 port map( A => n3795, ZN => n3806);
   U1969 : INV_X1 port map( A => n3806, ZN => n3807);
   U1971 : INV_X2 port map( A => n3806, ZN => n3809);
   U1973 : INV_X2 port map( A => n3806, ZN => n3808);
   U2008 : AND2_X4 port map( A1 => n1478, A2 => n141, ZN => n3810);
   U2043 : NAND2_X4 port map( A1 => n1343, A2 => n141, ZN => n1378);
   U2044 : AND2_X2 port map( A1 => n1309, A2 => n316, ZN => n1343);
   U2062 : AND2_X2 port map( A1 => n1309, A2 => n178, ZN => n1206);
   U2124 : CLKBUF_X3 port map( A => n3821, Z => n3811);
   U2126 : CLKBUF_X3 port map( A => n3821, Z => n3812);
   U2128 : CLKBUF_X3 port map( A => n3820, Z => n3813);
   U2130 : CLKBUF_X3 port map( A => n3820, Z => n3814);
   U2132 : CLKBUF_X3 port map( A => n3820, Z => n3815);
   U2134 : CLKBUF_X3 port map( A => n3819, Z => n3816);
   U2136 : CLKBUF_X3 port map( A => n3819, Z => n3817);
   U2138 : CLKBUF_X3 port map( A => n3819, Z => n3818);
   U2145 : CLKBUF_X3 port map( A => Reset, Z => n3819);
   U2146 : CLKBUF_X3 port map( A => Reset, Z => n3820);
   U2148 : CLKBUF_X3 port map( A => Reset, Z => n3821);
   U2150 : CLKBUF_X1 port map( A => n3976, Z => n3822);
   U2152 : CLKBUF_X1 port map( A => n3975, Z => n3823);
   U2154 : CLKBUF_X1 port map( A => n3975, Z => n3824);
   U2156 : CLKBUF_X1 port map( A => n3975, Z => n3825);
   U2176 : CLKBUF_X1 port map( A => n3975, Z => n3826);
   U2178 : CLKBUF_X1 port map( A => n3975, Z => n3827);
   U2182 : CLKBUF_X1 port map( A => n3975, Z => n3828);
   U2184 : CLKBUF_X1 port map( A => n3974, Z => n3829);
   U2190 : CLKBUF_X1 port map( A => n3974, Z => n3830);
   U2194 : CLKBUF_X1 port map( A => n3974, Z => n3831);
   U2225 : CLKBUF_X1 port map( A => n3974, Z => n3832);
   U2231 : CLKBUF_X1 port map( A => n3974, Z => n3833);
   U2235 : CLKBUF_X1 port map( A => n3974, Z => n3834);
   U2242 : CLKBUF_X1 port map( A => n3973, Z => n3835);
   U2244 : CLKBUF_X1 port map( A => n3973, Z => n3836);
   U2246 : CLKBUF_X1 port map( A => n3973, Z => n3837);
   U2248 : CLKBUF_X1 port map( A => n3973, Z => n3838);
   U2250 : CLKBUF_X1 port map( A => n3973, Z => n3839);
   U2252 : CLKBUF_X1 port map( A => n3973, Z => n3840);
   U2254 : CLKBUF_X1 port map( A => n3972, Z => n3841);
   U2256 : CLKBUF_X1 port map( A => n3972, Z => n3842);
   U2258 : CLKBUF_X1 port map( A => n3972, Z => n3843);
   U2260 : CLKBUF_X1 port map( A => n3972, Z => n3844);
   U2262 : CLKBUF_X1 port map( A => n3972, Z => n3845);
   U2264 : CLKBUF_X1 port map( A => n3972, Z => n3846);
   U2266 : CLKBUF_X1 port map( A => n3971, Z => n3847);
   U2276 : CLKBUF_X1 port map( A => n3971, Z => n3848);
   U2278 : CLKBUF_X1 port map( A => n3971, Z => n3849);
   U2280 : CLKBUF_X1 port map( A => n3971, Z => n3850);
   U2282 : CLKBUF_X1 port map( A => n3971, Z => n3851);
   U2284 : CLKBUF_X1 port map( A => n3971, Z => n3852);
   U2286 : CLKBUF_X1 port map( A => n3970, Z => n3853);
   U2288 : CLKBUF_X1 port map( A => n3970, Z => n3854);
   U2290 : CLKBUF_X1 port map( A => n3970, Z => n3855);
   U2292 : CLKBUF_X1 port map( A => n3970, Z => n3856);
   U2294 : CLKBUF_X1 port map( A => n3970, Z => n3857);
   U2296 : CLKBUF_X1 port map( A => n3970, Z => n3858);
   U2298 : CLKBUF_X1 port map( A => n3969, Z => n3859);
   U2300 : CLKBUF_X1 port map( A => n3969, Z => n3860);
   U2302 : CLKBUF_X1 port map( A => n3969, Z => n3861);
   U2322 : CLKBUF_X1 port map( A => n3969, Z => n3862);
   U2345 : CLKBUF_X1 port map( A => n3969, Z => n3863);
   U2355 : CLKBUF_X1 port map( A => n3969, Z => n3864);
   U2363 : CLKBUF_X1 port map( A => n3968, Z => n3865);
   U2365 : CLKBUF_X1 port map( A => n3968, Z => n3866);
   U2366 : CLKBUF_X1 port map( A => n3968, Z => n3867);
   U2367 : CLKBUF_X1 port map( A => n3968, Z => n3868);
   U2382 : CLKBUF_X1 port map( A => n3968, Z => n3869);
   U2384 : CLKBUF_X1 port map( A => n3968, Z => n3870);
   U2385 : CLKBUF_X1 port map( A => n3967, Z => n3871);
   U2400 : CLKBUF_X1 port map( A => n3967, Z => n3872);
   U2401 : CLKBUF_X1 port map( A => n3967, Z => n3873);
   U2416 : CLKBUF_X1 port map( A => n3967, Z => n3874);
   U2417 : CLKBUF_X1 port map( A => n3967, Z => n3875);
   U2418 : CLKBUF_X1 port map( A => n3967, Z => n3876);
   U2419 : CLKBUF_X1 port map( A => n3966, Z => n3877);
   U2434 : CLKBUF_X1 port map( A => n3966, Z => n3878);
   U2435 : CLKBUF_X1 port map( A => n3966, Z => n3879);
   U2436 : CLKBUF_X1 port map( A => n3966, Z => n3880);
   U2440 : CLKBUF_X1 port map( A => n3966, Z => n3881);
   U2442 : CLKBUF_X1 port map( A => n3966, Z => n3882);
   U2444 : CLKBUF_X1 port map( A => n3965, Z => n3883);
   U2446 : CLKBUF_X1 port map( A => n3965, Z => n3884);
   U2448 : CLKBUF_X1 port map( A => n3965, Z => n3885);
   U2450 : CLKBUF_X1 port map( A => n3965, Z => n3886);
   U2452 : CLKBUF_X1 port map( A => n3965, Z => n3887);
   U2454 : CLKBUF_X1 port map( A => n3965, Z => n3888);
   U2456 : CLKBUF_X1 port map( A => n3964, Z => n3889);
   U2458 : CLKBUF_X1 port map( A => n3964, Z => n3890);
   U2460 : CLKBUF_X1 port map( A => n3964, Z => n3891);
   U2462 : CLKBUF_X1 port map( A => n3964, Z => n3892);
   U2464 : CLKBUF_X1 port map( A => n3964, Z => n3893);
   U2465 : CLKBUF_X1 port map( A => n3964, Z => n3894);
   U2475 : CLKBUF_X1 port map( A => n3963, Z => n3895);
   U2477 : CLKBUF_X1 port map( A => n3963, Z => n3896);
   U2479 : CLKBUF_X1 port map( A => n3963, Z => n3897);
   U2481 : CLKBUF_X1 port map( A => n3963, Z => n3898);
   U2483 : CLKBUF_X1 port map( A => n3963, Z => n3899);
   U2485 : CLKBUF_X1 port map( A => n3963, Z => n3900);
   U2487 : CLKBUF_X1 port map( A => n3962, Z => n3901);
   U2489 : CLKBUF_X1 port map( A => n3962, Z => n3902);
   U2491 : CLKBUF_X1 port map( A => n3962, Z => n3903);
   U2493 : CLKBUF_X1 port map( A => n3962, Z => n3904);
   U2495 : CLKBUF_X1 port map( A => n3962, Z => n3905);
   U2497 : CLKBUF_X1 port map( A => n3962, Z => n3906);
   U2499 : CLKBUF_X1 port map( A => n3961, Z => n3907);
   U2501 : CLKBUF_X1 port map( A => n3961, Z => n3908);
   U2502 : CLKBUF_X1 port map( A => n3961, Z => n3909);
   U2503 : CLKBUF_X1 port map( A => n3961, Z => n3910);
   U2505 : CLKBUF_X1 port map( A => n3961, Z => n3911);
   U2507 : CLKBUF_X1 port map( A => n3961, Z => n3912);
   U2509 : CLKBUF_X1 port map( A => n3960, Z => n3913);
   U2511 : CLKBUF_X1 port map( A => n3960, Z => n3914);
   U2513 : CLKBUF_X1 port map( A => n3960, Z => n3915);
   U2515 : CLKBUF_X1 port map( A => n3960, Z => n3916);
   U2517 : CLKBUF_X1 port map( A => n3960, Z => n3917);
   U2519 : CLKBUF_X1 port map( A => n3960, Z => n3918);
   U2521 : CLKBUF_X1 port map( A => n3959, Z => n3919);
   U2523 : CLKBUF_X1 port map( A => n3959, Z => n3920);
   U2525 : CLKBUF_X1 port map( A => n3959, Z => n3921);
   U2527 : CLKBUF_X1 port map( A => n3959, Z => n3922);
   U2529 : CLKBUF_X1 port map( A => n3959, Z => n3923);
   U2530 : CLKBUF_X1 port map( A => n3959, Z => n3924);
   U2533 : CLKBUF_X1 port map( A => n3958, Z => n3925);
   U2539 : CLKBUF_X1 port map( A => n3958, Z => n3926);
   U2541 : CLKBUF_X1 port map( A => n3958, Z => n3927);
   U2543 : CLKBUF_X1 port map( A => n3958, Z => n3928);
   U2545 : CLKBUF_X1 port map( A => n3958, Z => n3929);
   U2547 : CLKBUF_X1 port map( A => n3958, Z => n3930);
   U2549 : CLKBUF_X1 port map( A => n3957, Z => n3931);
   U2551 : CLKBUF_X1 port map( A => n3957, Z => n3932);
   U2553 : CLKBUF_X1 port map( A => n3957, Z => n3933);
   U2555 : CLKBUF_X1 port map( A => n3957, Z => n3934);
   U2557 : CLKBUF_X1 port map( A => n3957, Z => n3935);
   U2559 : CLKBUF_X1 port map( A => n3957, Z => n3936);
   U2561 : CLKBUF_X1 port map( A => n3956, Z => n3937);
   U2563 : CLKBUF_X1 port map( A => n3956, Z => n3938);
   U2565 : CLKBUF_X1 port map( A => n3956, Z => n3939);
   U2566 : CLKBUF_X1 port map( A => n3956, Z => n3940);
   U2567 : CLKBUF_X1 port map( A => n3956, Z => n3941);
   U2581 : CLKBUF_X1 port map( A => n3956, Z => n3942);
   U2584 : CLKBUF_X1 port map( A => n3955, Z => n3943);
   U2600 : CLKBUF_X1 port map( A => n3955, Z => n3944);
   U2601 : CLKBUF_X1 port map( A => n3955, Z => n3945);
   U2615 : CLKBUF_X1 port map( A => n3955, Z => n3946);
   U2617 : CLKBUF_X1 port map( A => n3955, Z => n3947);
   U2618 : CLKBUF_X1 port map( A => n3955, Z => n3948);
   U2634 : CLKBUF_X1 port map( A => n3954, Z => n3949);
   U2635 : CLKBUF_X1 port map( A => n3954, Z => n3950);
   U2636 : CLKBUF_X1 port map( A => n3954, Z => n3951);
   U2639 : CLKBUF_X1 port map( A => n3954, Z => n3952);
   U2641 : CLKBUF_X1 port map( A => n3954, Z => n3953);
   U2643 : CLKBUF_X3 port map( A => n3811, Z => n3954);
   U2645 : CLKBUF_X3 port map( A => n3811, Z => n3955);
   U2647 : CLKBUF_X3 port map( A => n3811, Z => n3956);
   U2649 : CLKBUF_X3 port map( A => n3812, Z => n3957);
   U2651 : CLKBUF_X3 port map( A => n3812, Z => n3958);
   U2653 : CLKBUF_X3 port map( A => n3812, Z => n3959);
   U2655 : CLKBUF_X3 port map( A => n3813, Z => n3960);
   U2657 : CLKBUF_X3 port map( A => n3813, Z => n3961);
   U2659 : CLKBUF_X3 port map( A => n3813, Z => n3962);
   U2661 : CLKBUF_X3 port map( A => n3814, Z => n3963);
   U2663 : CLKBUF_X3 port map( A => n3814, Z => n3964);
   U2664 : CLKBUF_X3 port map( A => n3814, Z => n3965);
   U2665 : CLKBUF_X3 port map( A => n3815, Z => n3966);
   U2673 : CLKBUF_X3 port map( A => n3815, Z => n3967);
   U2675 : CLKBUF_X3 port map( A => n3815, Z => n3968);
   U2677 : CLKBUF_X3 port map( A => n3816, Z => n3969);
   U2679 : CLKBUF_X3 port map( A => n3816, Z => n3970);
   U2681 : CLKBUF_X3 port map( A => n3816, Z => n3971);
   U2683 : CLKBUF_X3 port map( A => n3817, Z => n3972);
   U2685 : CLKBUF_X3 port map( A => n3817, Z => n3973);
   U2687 : CLKBUF_X3 port map( A => n3817, Z => n3974);
   U2689 : CLKBUF_X3 port map( A => n3818, Z => n3975);
   U2691 : CLKBUF_X3 port map( A => n3818, Z => n3976);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity datapath_NUMBIT32_ADDRESS_WIDTH_RF5_ADDRESS_WIDTH_DM32 is

   port( CLK, RST : in std_logic;  INP1 : in std_logic_vector (31 downto 0);  
         INP2 : in std_logic_vector (15 downto 0);  IMM26 : in std_logic_vector
         (25 downto 0);  RS1, RS2, RD : in std_logic_vector (4 downto 0);  
         REGF_LATCH_EN, RegA_LATCH_EN, RegB_LATCH_EN, RegIMM_LATCH_EN, 
         RegRD1_LATCH_EN, SIGN_UNSIGN, RFR1_EN, RFR2_EN, MUX_IMM_SEL, JUMP, 
         JUMP_EN, EQ_COND, MUXA_SEL, MUXB_SEL, RALUOUT_LATCH_EN, REGME_LATCH_EN
         , RegRD2_LATCH_EN : in std_logic;  ALU_OPCODE : in std_logic_vector (0
         to 4);  ADDR_DRAM, DATAIN_DRAM : out std_logic_vector (31 downto 0);  
         DATAOUT_DRAM : in std_logic_vector (31 downto 0);  LMD_LATCH_EN, 
         RALUOUT2_LATCH_EN, RegRD3_LATCH_EN, RPCplus8_LATCH_EN, WB_MUX_SEL, 
         RF_WE, ROUT_LATCH_EN, JandL : in std_logic;  BRANCH_CTRL_SIG : out 
         std_logic;  BRANCH_ALU_OUT, Data_out : out std_logic_vector (31 downto
         0);  REGWRITE_XM, REGWRITE_MW : in std_logic);

end datapath_NUMBIT32_ADDRESS_WIDTH_RF5_ADDRESS_WIDTH_DM32;

architecture SYN_Struct of 
   datapath_NUMBIT32_ADDRESS_WIDTH_RF5_ADDRESS_WIDTH_DM32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X2
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component ForwardingUnit_NUMBIT32_ADDRESS_WIDTH_RF5
      port( CLK, RST : in std_logic;  RS1, RS2, RD_XM, RD_MW : in 
            std_logic_vector (4 downto 0);  REGWRITE_XM, REGWRITE_MW : in 
            std_logic;  ForwardA, forwardB : out std_logic_vector (1 downto 0);
            ForwardC : out std_logic;  ForwardD : out std_logic_vector (1 
            downto 0));
   end component;
   
   component MUX21_GENERIC_N32_1
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_N5
      port( A, B : in std_logic_vector (4 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (4 downto 0));
   end component;
   
   component reg_NUMBIT32_1
      port( clk, en, rst : in std_logic;  d : in std_logic_vector (31 downto 0)
            ;  q : out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_N32_2
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_N32_3
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component reg_NUMBIT32_2
      port( clk, en, rst : in std_logic;  d : in std_logic_vector (31 downto 0)
            ;  q : out std_logic_vector (31 downto 0));
   end component;
   
   component reg_NUMBIT5_1
      port( clk, en, rst : in std_logic;  d : in std_logic_vector (4 downto 0);
            q : out std_logic_vector (4 downto 0));
   end component;
   
   component reg_NUMBIT32_3
      port( clk, en, rst : in std_logic;  d : in std_logic_vector (31 downto 0)
            ;  q : out std_logic_vector (31 downto 0));
   end component;
   
   component reg_NUMBIT32_4
      port( clk, en, rst : in std_logic;  d : in std_logic_vector (31 downto 0)
            ;  q : out std_logic_vector (31 downto 0));
   end component;
   
   component reg_NUMBIT5_2
      port( clk, en, rst : in std_logic;  d : in std_logic_vector (4 downto 0);
            q : out std_logic_vector (4 downto 0));
   end component;
   
   component reg_NUMBIT32_5
      port( clk, en, rst : in std_logic;  d : in std_logic_vector (31 downto 0)
            ;  q : out std_logic_vector (31 downto 0));
   end component;
   
   component reg_NUMBIT32_6
      port( clk, en, rst : in std_logic;  d : in std_logic_vector (31 downto 0)
            ;  q : out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_N32_4
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_N32_5
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21
      port( A, B, SEL : in std_logic;  Y : out std_logic);
   end component;
   
   component BranchMgmt_NUMBIT32
      port( Rin : in std_logic_vector (31 downto 0);  Cond, Jump : in std_logic
            ;  Branch : out std_logic);
   end component;
   
   component reg_NUMBIT5_0
      port( clk, en, rst : in std_logic;  d : in std_logic_vector (4 downto 0);
            q : out std_logic_vector (4 downto 0));
   end component;
   
   component reg_NUMBIT32_7
      port( clk, en, rst : in std_logic;  d : in std_logic_vector (31 downto 0)
            ;  q : out std_logic_vector (31 downto 0));
   end component;
   
   component reg_NUMBIT32_8
      port( clk, en, rst : in std_logic;  d : in std_logic_vector (31 downto 0)
            ;  q : out std_logic_vector (31 downto 0));
   end component;
   
   component reg_NUMBIT32_9
      port( clk, en, rst : in std_logic;  d : in std_logic_vector (31 downto 0)
            ;  q : out std_logic_vector (31 downto 0));
   end component;
   
   component reg_NUMBIT32_0
      port( clk, en, rst : in std_logic;  d : in std_logic_vector (31 downto 0)
            ;  q : out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_N32_0
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component signExtend_NUMBIT_in26_NUMBIT_out32
      port( in_s : in std_logic_vector (25 downto 0);  sign_unsign : in 
            std_logic;  out_s : out std_logic_vector (31 downto 0));
   end component;
   
   component signExtend_NUMBIT_in16_NUMBIT_out32
      port( in_s : in std_logic_vector (15 downto 0);  sign_unsign : in 
            std_logic;  out_s : out std_logic_vector (31 downto 0));
   end component;
   
   component register_file_NUMBIT32_BITADDR5
      port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
            ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
            std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X4
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component alu_NUMBIT32
      port( DATA1, DATA2 : in std_logic_vector (31 downto 0);  FUNC : in 
            std_logic_vector (0 to 4);  OUTALU : out std_logic_vector (31 
            downto 0));
   end component;
   
   component P4addersub_N32
      port( A, B : in std_logic_vector (31 downto 0);  sub_add : in std_logic; 
            Y : out std_logic_vector (31 downto 0);  Cout : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, ADDR_DRAM_31_port, ADDR_DRAM_30_port, 
      ADDR_DRAM_29_port, ADDR_DRAM_28_port, ADDR_DRAM_27_port, 
      ADDR_DRAM_26_port, ADDR_DRAM_25_port, ADDR_DRAM_24_port, 
      ADDR_DRAM_23_port, ADDR_DRAM_22_port, ADDR_DRAM_21_port, 
      ADDR_DRAM_20_port, ADDR_DRAM_19_port, ADDR_DRAM_18_port, 
      ADDR_DRAM_17_port, ADDR_DRAM_16_port, ADDR_DRAM_15_port, 
      ADDR_DRAM_14_port, ADDR_DRAM_13_port, ADDR_DRAM_12_port, 
      ADDR_DRAM_11_port, ADDR_DRAM_10_port, ADDR_DRAM_9_port, ADDR_DRAM_8_port,
      ADDR_DRAM_7_port, ADDR_DRAM_6_port, ADDR_DRAM_5_port, ADDR_DRAM_4_port, 
      ADDR_DRAM_3_port, ADDR_DRAM_2_port, ADDR_DRAM_1_port, ADDR_DRAM_0_port, 
      n214, n215, n216, MUX_WRaddr_OUT_4_port, MUX_WRaddr_OUT_3_port, 
      MUX_WRaddr_OUT_2_port, MUX_WRaddr_OUT_1_port, MUX_WRaddr_OUT_0_port, 
      MUX_WRdata_OUT_31_port, MUX_WRdata_OUT_30_port, MUX_WRdata_OUT_29_port, 
      MUX_WRdata_OUT_28_port, MUX_WRdata_OUT_27_port, MUX_WRdata_OUT_26_port, 
      MUX_WRdata_OUT_25_port, MUX_WRdata_OUT_24_port, MUX_WRdata_OUT_23_port, 
      MUX_WRdata_OUT_22_port, MUX_WRdata_OUT_21_port, MUX_WRdata_OUT_20_port, 
      MUX_WRdata_OUT_19_port, MUX_WRdata_OUT_18_port, MUX_WRdata_OUT_17_port, 
      MUX_WRdata_OUT_16_port, MUX_WRdata_OUT_15_port, MUX_WRdata_OUT_14_port, 
      MUX_WRdata_OUT_13_port, MUX_WRdata_OUT_12_port, MUX_WRdata_OUT_11_port, 
      MUX_WRdata_OUT_10_port, MUX_WRdata_OUT_9_port, MUX_WRdata_OUT_8_port, 
      MUX_WRdata_OUT_7_port, MUX_WRdata_OUT_6_port, MUX_WRdata_OUT_5_port, 
      MUX_WRdata_OUT_4_port, MUX_WRdata_OUT_3_port, MUX_WRdata_OUT_2_port, 
      MUX_WRdata_OUT_1_port, MUX_WRdata_OUT_0_port, RA_IN_31_port, 
      RA_IN_30_port, RA_IN_29_port, RA_IN_28_port, RA_IN_27_port, RA_IN_26_port
      , RA_IN_25_port, RA_IN_24_port, RA_IN_23_port, RA_IN_22_port, 
      RA_IN_21_port, RA_IN_20_port, RA_IN_19_port, RA_IN_18_port, RA_IN_17_port
      , RA_IN_16_port, RA_IN_15_port, RA_IN_14_port, RA_IN_13_port, 
      RA_IN_12_port, RA_IN_11_port, RA_IN_10_port, RA_IN_9_port, RA_IN_8_port, 
      RA_IN_7_port, RA_IN_6_port, RA_IN_5_port, RA_IN_4_port, RA_IN_3_port, 
      RA_IN_2_port, RA_IN_1_port, RA_IN_0_port, RB_IN_31_port, RB_IN_30_port, 
      RB_IN_29_port, RB_IN_28_port, RB_IN_27_port, RB_IN_26_port, RB_IN_25_port
      , RB_IN_24_port, RB_IN_23_port, RB_IN_22_port, RB_IN_21_port, 
      RB_IN_20_port, RB_IN_19_port, RB_IN_18_port, RB_IN_17_port, RB_IN_16_port
      , RB_IN_15_port, RB_IN_14_port, RB_IN_13_port, RB_IN_12_port, 
      RB_IN_11_port, RB_IN_10_port, RB_IN_9_port, RB_IN_8_port, RB_IN_7_port, 
      RB_IN_6_port, RB_IN_5_port, RB_IN_4_port, RB_IN_3_port, RB_IN_2_port, 
      RB_IN_1_port, RB_IN_0_port, SIGNEXT_IMP2_31_port, SIGNEXT_IMP2_30_port, 
      SIGNEXT_IMP2_29_port, SIGNEXT_IMP2_28_port, SIGNEXT_IMP2_27_port, 
      SIGNEXT_IMP2_26_port, SIGNEXT_IMP2_25_port, SIGNEXT_IMP2_24_port, 
      SIGNEXT_IMP2_23_port, SIGNEXT_IMP2_22_port, SIGNEXT_IMP2_21_port, 
      SIGNEXT_IMP2_20_port, SIGNEXT_IMP2_19_port, SIGNEXT_IMP2_18_port, 
      SIGNEXT_IMP2_17_port, SIGNEXT_IMP2_16_port, SIGNEXT_IMP2_15_port, 
      SIGNEXT_IMP2_14_port, SIGNEXT_IMP2_13_port, SIGNEXT_IMP2_12_port, 
      SIGNEXT_IMP2_11_port, SIGNEXT_IMP2_10_port, SIGNEXT_IMP2_9_port, 
      SIGNEXT_IMP2_8_port, SIGNEXT_IMP2_7_port, SIGNEXT_IMP2_6_port, 
      SIGNEXT_IMP2_5_port, SIGNEXT_IMP2_4_port, SIGNEXT_IMP2_3_port, 
      SIGNEXT_IMP2_2_port, SIGNEXT_IMP2_1_port, SIGNEXT_IMP2_0_port, 
      SIGNEXT_IMM26_31_port, SIGNEXT_IMM26_30_port, SIGNEXT_IMM26_29_port, 
      SIGNEXT_IMM26_28_port, SIGNEXT_IMM26_27_port, SIGNEXT_IMM26_26_port, 
      SIGNEXT_IMM26_25_port, SIGNEXT_IMM26_24_port, SIGNEXT_IMM26_23_port, 
      SIGNEXT_IMM26_22_port, SIGNEXT_IMM26_21_port, SIGNEXT_IMM26_20_port, 
      SIGNEXT_IMM26_19_port, SIGNEXT_IMM26_18_port, SIGNEXT_IMM26_17_port, 
      SIGNEXT_IMM26_16_port, SIGNEXT_IMM26_15_port, SIGNEXT_IMM26_14_port, 
      SIGNEXT_IMM26_13_port, SIGNEXT_IMM26_12_port, SIGNEXT_IMM26_11_port, 
      SIGNEXT_IMM26_10_port, SIGNEXT_IMM26_9_port, SIGNEXT_IMM26_8_port, 
      SIGNEXT_IMM26_7_port, SIGNEXT_IMM26_6_port, SIGNEXT_IMM26_5_port, 
      SIGNEXT_IMM26_4_port, SIGNEXT_IMM26_3_port, SIGNEXT_IMM26_2_port, 
      SIGNEXT_IMM26_1_port, SIGNEXT_IMM26_0_port, MUX_IMM_OUT_31_port, 
      MUX_IMM_OUT_30_port, MUX_IMM_OUT_29_port, MUX_IMM_OUT_28_port, 
      MUX_IMM_OUT_27_port, MUX_IMM_OUT_26_port, MUX_IMM_OUT_25_port, 
      MUX_IMM_OUT_24_port, MUX_IMM_OUT_23_port, MUX_IMM_OUT_22_port, 
      MUX_IMM_OUT_21_port, MUX_IMM_OUT_20_port, MUX_IMM_OUT_19_port, 
      MUX_IMM_OUT_18_port, MUX_IMM_OUT_17_port, MUX_IMM_OUT_16_port, 
      MUX_IMM_OUT_15_port, MUX_IMM_OUT_14_port, MUX_IMM_OUT_13_port, 
      MUX_IMM_OUT_12_port, MUX_IMM_OUT_11_port, MUX_IMM_OUT_10_port, 
      MUX_IMM_OUT_9_port, MUX_IMM_OUT_8_port, MUX_IMM_OUT_7_port, 
      MUX_IMM_OUT_6_port, MUX_IMM_OUT_5_port, MUX_IMM_OUT_4_port, 
      MUX_IMM_OUT_3_port, MUX_IMM_OUT_2_port, RA_OUT_31_port, RA_OUT_30_port, 
      RA_OUT_29_port, RA_OUT_28_port, RA_OUT_27_port, RA_OUT_26_port, 
      RA_OUT_25_port, RA_OUT_24_port, RA_OUT_23_port, RA_OUT_22_port, 
      RA_OUT_21_port, RA_OUT_20_port, RA_OUT_19_port, RA_OUT_18_port, 
      RA_OUT_17_port, RA_OUT_16_port, RA_OUT_15_port, RA_OUT_14_port, 
      RA_OUT_13_port, RA_OUT_12_port, RA_OUT_11_port, RA_OUT_10_port, 
      RA_OUT_9_port, RA_OUT_8_port, RA_OUT_7_port, RA_OUT_6_port, RA_OUT_5_port
      , RA_OUT_4_port, RA_OUT_3_port, RA_OUT_2_port, RA_OUT_1_port, 
      RA_OUT_0_port, RB_OUT_31_port, RB_OUT_30_port, RB_OUT_29_port, 
      RB_OUT_28_port, RB_OUT_27_port, RB_OUT_26_port, RB_OUT_25_port, 
      RB_OUT_24_port, RB_OUT_23_port, RB_OUT_22_port, RB_OUT_21_port, 
      RB_OUT_20_port, RB_OUT_19_port, RB_OUT_18_port, RB_OUT_17_port, 
      RB_OUT_16_port, RB_OUT_15_port, RB_OUT_14_port, RB_OUT_13_port, 
      RB_OUT_12_port, RB_OUT_11_port, RB_OUT_10_port, RB_OUT_9_port, 
      RB_OUT_8_port, RB_OUT_7_port, RB_OUT_6_port, RB_OUT_5_port, RB_OUT_4_port
      , RB_OUT_3_port, RB_OUT_2_port, RB_OUT_1_port, RB_OUT_0_port, 
      MUX_FORWARDING_BRANCH_OUT_31_port, MUX_FORWARDING_BRANCH_OUT_30_port, 
      MUX_FORWARDING_BRANCH_OUT_29_port, MUX_FORWARDING_BRANCH_OUT_28_port, 
      MUX_FORWARDING_BRANCH_OUT_27_port, MUX_FORWARDING_BRANCH_OUT_26_port, 
      MUX_FORWARDING_BRANCH_OUT_25_port, MUX_FORWARDING_BRANCH_OUT_24_port, 
      MUX_FORWARDING_BRANCH_OUT_23_port, MUX_FORWARDING_BRANCH_OUT_22_port, 
      MUX_FORWARDING_BRANCH_OUT_21_port, MUX_FORWARDING_BRANCH_OUT_20_port, 
      MUX_FORWARDING_BRANCH_OUT_19_port, MUX_FORWARDING_BRANCH_OUT_18_port, 
      MUX_FORWARDING_BRANCH_OUT_17_port, MUX_FORWARDING_BRANCH_OUT_16_port, 
      MUX_FORWARDING_BRANCH_OUT_15_port, MUX_FORWARDING_BRANCH_OUT_14_port, 
      MUX_FORWARDING_BRANCH_OUT_13_port, MUX_FORWARDING_BRANCH_OUT_12_port, 
      MUX_FORWARDING_BRANCH_OUT_11_port, MUX_FORWARDING_BRANCH_OUT_10_port, 
      MUX_FORWARDING_BRANCH_OUT_9_port, MUX_FORWARDING_BRANCH_OUT_8_port, 
      MUX_FORWARDING_BRANCH_OUT_7_port, MUX_FORWARDING_BRANCH_OUT_6_port, 
      MUX_FORWARDING_BRANCH_OUT_5_port, MUX_FORWARDING_BRANCH_OUT_4_port, 
      MUX_FORWARDING_BRANCH_OUT_3_port, MUX_FORWARDING_BRANCH_OUT_2_port, 
      MUX_FORWARDING_BRANCH_OUT_1_port, MUX_FORWARDING_BRANCH_OUT_0_port, 
      BRANCH_T_NT, MUXA_OUT_31_port, MUXA_OUT_30_port, MUXA_OUT_29_port, 
      MUXA_OUT_28_port, MUXA_OUT_27_port, MUXA_OUT_26_port, MUXA_OUT_25_port, 
      MUXA_OUT_24_port, MUXA_OUT_23_port, MUXA_OUT_22_port, MUXA_OUT_21_port, 
      MUXA_OUT_20_port, MUXA_OUT_19_port, MUXA_OUT_18_port, MUXA_OUT_17_port, 
      MUXA_OUT_16_port, MUXA_OUT_15_port, MUXA_OUT_14_port, MUXA_OUT_13_port, 
      MUXA_OUT_12_port, MUXA_OUT_11_port, MUXA_OUT_10_port, MUXA_OUT_9_port, 
      MUXA_OUT_8_port, MUXA_OUT_7_port, MUXA_OUT_6_port, MUXA_OUT_5_port, 
      MUXA_OUT_4_port, MUXA_OUT_3_port, MUXA_OUT_2_port, MUXA_OUT_1_port, 
      MUXA_OUT_0_port, ForwardD_1_port, ForwardD_0_port, MUXC_OUT_31_port, 
      MUXC_OUT_30_port, MUXC_OUT_29_port, MUXC_OUT_28_port, MUXC_OUT_27_port, 
      MUXC_OUT_26_port, MUXC_OUT_25_port, MUXC_OUT_24_port, MUXC_OUT_23_port, 
      MUXC_OUT_22_port, MUXC_OUT_21_port, MUXC_OUT_20_port, MUXC_OUT_19_port, 
      MUXC_OUT_18_port, MUXC_OUT_17_port, MUXC_OUT_16_port, MUXC_OUT_15_port, 
      MUXC_OUT_14_port, MUXC_OUT_13_port, MUXC_OUT_12_port, MUXC_OUT_11_port, 
      MUXC_OUT_10_port, MUXC_OUT_9_port, MUXC_OUT_8_port, MUXC_OUT_7_port, 
      MUXC_OUT_6_port, MUXC_OUT_5_port, MUXC_OUT_4_port, MUXC_OUT_3_port, 
      MUXC_OUT_2_port, MUXC_OUT_1_port, MUXC_OUT_0_port, ALU_inputB_31_port, 
      ALU_inputB_30_port, ALU_inputB_29_port, ALU_inputB_28_port, 
      ALU_inputB_27_port, ALU_inputB_26_port, ALU_inputB_25_port, 
      ALU_inputB_24_port, ALU_inputB_23_port, ALU_inputB_22_port, 
      ALU_inputB_21_port, ALU_inputB_20_port, ALU_inputB_19_port, 
      ALU_inputB_18_port, ALU_inputB_17_port, ALU_inputB_16_port, 
      ALU_inputB_15_port, ALU_inputB_14_port, ALU_inputB_13_port, 
      ALU_inputB_12_port, ALU_inputB_11_port, ALU_inputB_10_port, 
      ALU_inputB_9_port, ALU_inputB_8_port, ALU_inputB_7_port, 
      ALU_inputB_6_port, ALU_inputB_5_port, ALU_inputB_4_port, 
      ALU_inputB_3_port, ALU_inputB_2_port, ALU_inputB_1_port, 
      ALU_inputB_0_port, MUXB_OUT_31_port, MUXB_OUT_30_port, MUXB_OUT_29_port, 
      MUXB_OUT_28_port, MUXB_OUT_27_port, MUXB_OUT_26_port, MUXB_OUT_25_port, 
      MUXB_OUT_24_port, MUXB_OUT_23_port, MUXB_OUT_22_port, MUXB_OUT_21_port, 
      MUXB_OUT_20_port, MUXB_OUT_19_port, MUXB_OUT_18_port, MUXB_OUT_17_port, 
      MUXB_OUT_16_port, MUXB_OUT_15_port, MUXB_OUT_14_port, MUXB_OUT_13_port, 
      MUXB_OUT_12_port, MUXB_OUT_11_port, MUXB_OUT_10_port, MUXB_OUT_9_port, 
      MUXB_OUT_8_port, MUXB_OUT_7_port, MUXB_OUT_6_port, MUXB_OUT_5_port, 
      MUXB_OUT_4_port, MUXB_OUT_3_port, MUXB_OUT_2_port, MUXB_OUT_1_port, 
      MUXB_OUT_0_port, ALU_inputA_31_port, ALU_inputA_30_port, 
      ALU_inputA_29_port, ALU_inputA_28_port, ALU_inputA_27_port, 
      ALU_inputA_26_port, ALU_inputA_25_port, ALU_inputA_24_port, 
      ALU_inputA_23_port, ALU_inputA_22_port, ALU_inputA_21_port, 
      ALU_inputA_20_port, ALU_inputA_19_port, ALU_inputA_18_port, 
      ALU_inputA_17_port, ALU_inputA_16_port, ALU_inputA_15_port, 
      ALU_inputA_14_port, ALU_inputA_13_port, ALU_inputA_12_port, 
      ALU_inputA_11_port, ALU_inputA_10_port, ALU_inputA_9_port, 
      ALU_inputA_8_port, ALU_inputA_7_port, ALU_inputA_6_port, 
      ALU_inputA_5_port, ALU_inputA_4_port, ALU_inputA_3_port, 
      ALU_inputA_2_port, ALU_inputA_1_port, ALU_inputA_0_port, ALU_OUT_31_port,
      ALU_OUT_30_port, ALU_OUT_29_port, ALU_OUT_28_port, ALU_OUT_27_port, 
      ALU_OUT_26_port, ALU_OUT_25_port, ALU_OUT_24_port, ALU_OUT_23_port, 
      ALU_OUT_22_port, ALU_OUT_21_port, ALU_OUT_20_port, ALU_OUT_19_port, 
      ALU_OUT_18_port, ALU_OUT_17_port, ALU_OUT_16_port, ALU_OUT_15_port, 
      ALU_OUT_14_port, ALU_OUT_13_port, ALU_OUT_12_port, ALU_OUT_11_port, 
      ALU_OUT_10_port, ALU_OUT_9_port, ALU_OUT_8_port, ALU_OUT_7_port, 
      ALU_OUT_6_port, ALU_OUT_5_port, ALU_OUT_4_port, ALU_OUT_3_port, 
      ALU_OUT_2_port, ALU_OUT_1_port, ALU_OUT_0_port, RD2_OUT_4_port, 
      RD2_OUT_3_port, RD2_OUT_2_port, RD2_OUT_1_port, RD2_OUT_0_port, 
      ForwardA_1_port, ForwardA_0_port, forwardB_1_port, forwardB_0_port, 
      RD3_OUT_4_port, RD3_OUT_3_port, RD3_OUT_2_port, RD3_OUT_1_port, 
      RD3_OUT_0_port, ForwardC, net992, n2, n3, n4, n5, n6, n7, n8, n9, n10, 
      n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25
      , n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, 
      n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54
      , n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, 
      n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83
      , n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, 
      n99, n100, n101, n104, n106, n107, n108, n109, n110, n111, n112, n113, 
      n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, 
      n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n138, n139, 
      n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, net92960, 
      net92959, net92958, net94217, net94215, net94214, net95253, net95252, 
      net95311, net95310, net95343, net95342, net95411, net95416, net95415, 
      net95422, net95434, net95433, net95551, net95521, n98, n137, n136, n1, 
      n102, n103, n105, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n208, 
      n209, n210, RPCplus8_OUT_9_port, RPCplus8_OUT_8_port, RPCplus8_OUT_7_port
      , RPCplus8_OUT_6_port, RPCplus8_OUT_5_port, RPCplus8_OUT_4_port, 
      RPCplus8_OUT_3_port, RPCplus8_OUT_31_port, RPCplus8_OUT_30_port, 
      RPCplus8_OUT_2_port, RPCplus8_OUT_29_port, RPCplus8_OUT_28_port, 
      RPCplus8_OUT_27_port, RPCplus8_OUT_26_port, RPCplus8_OUT_25_port, 
      RPCplus8_OUT_24_port, RPCplus8_OUT_23_port, RPCplus8_OUT_22_port, 
      RPCplus8_OUT_21_port, RPCplus8_OUT_20_port, RPCplus8_OUT_1_port, 
      RPCplus8_OUT_19_port, RPCplus8_OUT_18_port, RPCplus8_OUT_17_port, 
      RPCplus8_OUT_16_port, RPCplus8_OUT_15_port, RPCplus8_OUT_14_port, 
      RPCplus8_OUT_13_port, RPCplus8_OUT_12_port, RPCplus8_OUT_11_port, 
      RPCplus8_OUT_10_port, RPCplus8_OUT_0_port, RME_OUT_9_port, RME_OUT_8_port
      , RME_OUT_7_port, RME_OUT_6_port, RME_OUT_5_port, RME_OUT_4_port, 
      RME_OUT_3_port, RME_OUT_31_port, RME_OUT_30_port, RME_OUT_2_port, 
      RME_OUT_29_port, RME_OUT_28_port, RME_OUT_27_port, RME_OUT_26_port, 
      RME_OUT_25_port, RME_OUT_24_port, RME_OUT_23_port, RME_OUT_22_port, 
      RME_OUT_21_port, RME_OUT_20_port, RME_OUT_1_port, RME_OUT_19_port, 
      RME_OUT_18_port, RME_OUT_17_port, RME_OUT_16_port, RME_OUT_15_port, 
      RME_OUT_14_port, RME_OUT_13_port, RME_OUT_12_port, RME_OUT_11_port, 
      RME_OUT_10_port, RME_OUT_0_port, RIMM2_OUT_9_port, RIMM2_OUT_8_port, 
      RIMM2_OUT_7_port, RIMM2_OUT_6_port, RIMM2_OUT_5_port, RIMM2_OUT_4_port, 
      RIMM2_OUT_3_port, RIMM2_OUT_31_port, RIMM2_OUT_30_port, RIMM2_OUT_2_port,
      RIMM2_OUT_29_port, RIMM2_OUT_28_port, RIMM2_OUT_27_port, 
      RIMM2_OUT_26_port, RIMM2_OUT_25_port, RIMM2_OUT_24_port, 
      RIMM2_OUT_23_port, RIMM2_OUT_22_port, RIMM2_OUT_21_port, 
      RIMM2_OUT_20_port, RIMM2_OUT_1_port, RIMM2_OUT_19_port, RIMM2_OUT_18_port
      , RIMM2_OUT_17_port, RIMM2_OUT_16_port, RIMM2_OUT_15_port, 
      RIMM2_OUT_14_port, RIMM2_OUT_13_port, RIMM2_OUT_12_port, 
      RIMM2_OUT_11_port, RIMM2_OUT_10_port, RIMM2_OUT_0_port, RIMM1_OUT_9_port,
      RIMM1_OUT_8_port, RIMM1_OUT_7_port, RIMM1_OUT_6_port, RIMM1_OUT_5_port, 
      RIMM1_OUT_4_port, RIMM1_OUT_3_port, RIMM1_OUT_31_port, RIMM1_OUT_30_port,
      RIMM1_OUT_2_port, RIMM1_OUT_29_port, RIMM1_OUT_28_port, RIMM1_OUT_27_port
      , RIMM1_OUT_26_port, RIMM1_OUT_25_port, RIMM1_OUT_24_port, 
      RIMM1_OUT_23_port, RIMM1_OUT_22_port, RIMM1_OUT_21_port, 
      RIMM1_OUT_20_port, RIMM1_OUT_1_port, RIMM1_OUT_19_port, RIMM1_OUT_18_port
      , RIMM1_OUT_17_port, RIMM1_OUT_16_port, RIMM1_OUT_15_port, 
      RIMM1_OUT_14_port, RIMM1_OUT_13_port, RIMM1_OUT_12_port, 
      RIMM1_OUT_11_port, RIMM1_OUT_10_port, RIMM1_OUT_0_port, RD1_OUT_4_port, 
      RD1_OUT_3_port, RD1_OUT_2_port, RD1_OUT_1_port, RD1_OUT_0_port, 
      RALUOUT2_OUT_9_port, RALUOUT2_OUT_8_port, RALUOUT2_OUT_7_port, 
      RALUOUT2_OUT_6_port, RALUOUT2_OUT_5_port, RALUOUT2_OUT_4_port, 
      RALUOUT2_OUT_3_port, RALUOUT2_OUT_31_port, RALUOUT2_OUT_30_port, 
      RALUOUT2_OUT_2_port, RALUOUT2_OUT_29_port, RALUOUT2_OUT_28_port, 
      RALUOUT2_OUT_27_port, RALUOUT2_OUT_26_port, RALUOUT2_OUT_25_port, 
      RALUOUT2_OUT_24_port, RALUOUT2_OUT_23_port, RALUOUT2_OUT_22_port, 
      RALUOUT2_OUT_21_port, RALUOUT2_OUT_20_port, RALUOUT2_OUT_1_port, 
      RALUOUT2_OUT_19_port, RALUOUT2_OUT_18_port, RALUOUT2_OUT_17_port, 
      RALUOUT2_OUT_16_port, RALUOUT2_OUT_15_port, RALUOUT2_OUT_14_port, 
      RALUOUT2_OUT_13_port, RALUOUT2_OUT_12_port, RALUOUT2_OUT_11_port, 
      RALUOUT2_OUT_10_port, RALUOUT2_OUT_0_port, MUX_IMM_OUT_1_port, 
      MUX_IMM_OUT_0_port, LMD_OUT_9_port, LMD_OUT_8_port, LMD_OUT_7_port, 
      LMD_OUT_6_port, LMD_OUT_5_port, LMD_OUT_4_port, LMD_OUT_3_port, 
      LMD_OUT_31_port, LMD_OUT_30_port, LMD_OUT_2_port, LMD_OUT_29_port, 
      LMD_OUT_28_port, LMD_OUT_27_port, LMD_OUT_26_port, LMD_OUT_25_port, 
      LMD_OUT_24_port, LMD_OUT_23_port, LMD_OUT_22_port, LMD_OUT_21_port, 
      LMD_OUT_20_port, LMD_OUT_1_port, LMD_OUT_19_port, LMD_OUT_18_port, 
      LMD_OUT_17_port, LMD_OUT_16_port, LMD_OUT_15_port, LMD_OUT_14_port, 
      LMD_OUT_13_port, LMD_OUT_12_port, LMD_OUT_11_port, LMD_OUT_10_port, 
      LMD_OUT_0_port, n217 : std_logic;

begin
   ADDR_DRAM <= ( ADDR_DRAM_31_port, ADDR_DRAM_30_port, ADDR_DRAM_29_port, 
      ADDR_DRAM_28_port, ADDR_DRAM_27_port, ADDR_DRAM_26_port, 
      ADDR_DRAM_25_port, ADDR_DRAM_24_port, ADDR_DRAM_23_port, 
      ADDR_DRAM_22_port, ADDR_DRAM_21_port, ADDR_DRAM_20_port, 
      ADDR_DRAM_19_port, ADDR_DRAM_18_port, ADDR_DRAM_17_port, 
      ADDR_DRAM_16_port, ADDR_DRAM_15_port, ADDR_DRAM_14_port, 
      ADDR_DRAM_13_port, ADDR_DRAM_12_port, ADDR_DRAM_11_port, 
      ADDR_DRAM_10_port, ADDR_DRAM_9_port, ADDR_DRAM_8_port, ADDR_DRAM_7_port, 
      ADDR_DRAM_6_port, ADDR_DRAM_5_port, ADDR_DRAM_4_port, ADDR_DRAM_3_port, 
      ADDR_DRAM_2_port, ADDR_DRAM_1_port, ADDR_DRAM_0_port );
   
   P4adder_branching : P4addersub_N32 port map( A(31) => MUXA_OUT_31_port, 
                           A(30) => MUXA_OUT_30_port, A(29) => MUXA_OUT_29_port
                           , A(28) => MUXA_OUT_28_port, A(27) => 
                           MUXA_OUT_27_port, A(26) => MUXA_OUT_26_port, A(25) 
                           => MUXA_OUT_25_port, A(24) => MUXA_OUT_24_port, 
                           A(23) => MUXA_OUT_23_port, A(22) => MUXA_OUT_22_port
                           , A(21) => MUXA_OUT_21_port, A(20) => 
                           MUXA_OUT_20_port, A(19) => MUXA_OUT_19_port, A(18) 
                           => MUXA_OUT_18_port, A(17) => MUXA_OUT_17_port, 
                           A(16) => MUXA_OUT_16_port, A(15) => MUXA_OUT_15_port
                           , A(14) => MUXA_OUT_14_port, A(13) => 
                           MUXA_OUT_13_port, A(12) => MUXA_OUT_12_port, A(11) 
                           => MUXA_OUT_11_port, A(10) => MUXA_OUT_10_port, A(9)
                           => MUXA_OUT_9_port, A(8) => MUXA_OUT_8_port, A(7) =>
                           MUXA_OUT_7_port, A(6) => MUXA_OUT_6_port, A(5) => 
                           MUXA_OUT_5_port, A(4) => MUXA_OUT_4_port, A(3) => 
                           MUXA_OUT_3_port, A(2) => MUXA_OUT_2_port, A(1) => 
                           MUXA_OUT_1_port, A(0) => MUXA_OUT_0_port, B(31) => 
                           MUX_IMM_OUT_31_port, B(30) => MUX_IMM_OUT_31_port, 
                           B(29) => MUX_IMM_OUT_31_port, B(28) => 
                           MUX_IMM_OUT_30_port, B(27) => MUX_IMM_OUT_29_port, 
                           B(26) => MUX_IMM_OUT_28_port, B(25) => 
                           MUX_IMM_OUT_27_port, B(24) => MUX_IMM_OUT_26_port, 
                           B(23) => MUX_IMM_OUT_25_port, B(22) => 
                           MUX_IMM_OUT_24_port, B(21) => MUX_IMM_OUT_23_port, 
                           B(20) => MUX_IMM_OUT_22_port, B(19) => 
                           MUX_IMM_OUT_21_port, B(18) => MUX_IMM_OUT_20_port, 
                           B(17) => MUX_IMM_OUT_19_port, B(16) => 
                           MUX_IMM_OUT_18_port, B(15) => MUX_IMM_OUT_17_port, 
                           B(14) => MUX_IMM_OUT_16_port, B(13) => 
                           MUX_IMM_OUT_15_port, B(12) => MUX_IMM_OUT_14_port, 
                           B(11) => MUX_IMM_OUT_13_port, B(10) => 
                           MUX_IMM_OUT_12_port, B(9) => MUX_IMM_OUT_11_port, 
                           B(8) => MUX_IMM_OUT_10_port, B(7) => 
                           MUX_IMM_OUT_9_port, B(6) => MUX_IMM_OUT_8_port, B(5)
                           => MUX_IMM_OUT_7_port, B(4) => MUX_IMM_OUT_6_port, 
                           B(3) => MUX_IMM_OUT_5_port, B(2) => 
                           MUX_IMM_OUT_4_port, B(1) => MUX_IMM_OUT_3_port, B(0)
                           => MUX_IMM_OUT_2_port, sub_add => X_Logic0_port, 
                           Y(31) => BRANCH_ALU_OUT(31), Y(30) => n214, Y(29) =>
                           BRANCH_ALU_OUT(29), Y(28) => BRANCH_ALU_OUT(28), 
                           Y(27) => BRANCH_ALU_OUT(27), Y(26) => 
                           BRANCH_ALU_OUT(26), Y(25) => n215, Y(24) => 
                           BRANCH_ALU_OUT(24), Y(23) => n216, Y(22) => 
                           BRANCH_ALU_OUT(22), Y(21) => BRANCH_ALU_OUT(21), 
                           Y(20) => BRANCH_ALU_OUT(20), Y(19) => 
                           BRANCH_ALU_OUT(19), Y(18) => BRANCH_ALU_OUT(18), 
                           Y(17) => BRANCH_ALU_OUT(17), Y(16) => 
                           BRANCH_ALU_OUT(16), Y(15) => BRANCH_ALU_OUT(15), 
                           Y(14) => BRANCH_ALU_OUT(14), Y(13) => 
                           BRANCH_ALU_OUT(13), Y(12) => BRANCH_ALU_OUT(12), 
                           Y(11) => BRANCH_ALU_OUT(11), Y(10) => 
                           BRANCH_ALU_OUT(10), Y(9) => BRANCH_ALU_OUT(9), Y(8) 
                           => BRANCH_ALU_OUT(8), Y(7) => BRANCH_ALU_OUT(7), 
                           Y(6) => BRANCH_ALU_OUT(6), Y(5) => BRANCH_ALU_OUT(5)
                           , Y(4) => BRANCH_ALU_OUT(4), Y(3) => 
                           BRANCH_ALU_OUT(3), Y(2) => BRANCH_ALU_OUT(2), Y(1) 
                           => BRANCH_ALU_OUT(1), Y(0) => BRANCH_ALU_OUT(0), 
                           Cout => net992);
   alu_0 : alu_NUMBIT32 port map( DATA1(31) => ALU_inputA_31_port, DATA1(30) =>
                           n186, DATA1(29) => ALU_inputA_29_port, DATA1(28) => 
                           ALU_inputA_28_port, DATA1(27) => ALU_inputA_27_port,
                           DATA1(26) => ALU_inputA_26_port, DATA1(25) => 
                           ALU_inputA_25_port, DATA1(24) => ALU_inputA_24_port,
                           DATA1(23) => ALU_inputA_23_port, DATA1(22) => 
                           ALU_inputA_22_port, DATA1(21) => ALU_inputA_21_port,
                           DATA1(20) => ALU_inputA_20_port, DATA1(19) => 
                           ALU_inputA_19_port, DATA1(18) => ALU_inputA_18_port,
                           DATA1(17) => ALU_inputA_17_port, DATA1(16) => 
                           ALU_inputA_16_port, DATA1(15) => ALU_inputA_15_port,
                           DATA1(14) => ALU_inputA_14_port, DATA1(13) => 
                           ALU_inputA_13_port, DATA1(12) => ALU_inputA_12_port,
                           DATA1(11) => ALU_inputA_11_port, DATA1(10) => 
                           ALU_inputA_10_port, DATA1(9) => ALU_inputA_9_port, 
                           DATA1(8) => ALU_inputA_8_port, DATA1(7) => 
                           ALU_inputA_7_port, DATA1(6) => ALU_inputA_6_port, 
                           DATA1(5) => ALU_inputA_5_port, DATA1(4) => 
                           ALU_inputA_4_port, DATA1(3) => ALU_inputA_3_port, 
                           DATA1(2) => ALU_inputA_2_port, DATA1(1) => 
                           ALU_inputA_1_port, DATA1(0) => ALU_inputA_0_port, 
                           DATA2(31) => MUXB_OUT_31_port, DATA2(30) => 
                           MUXB_OUT_30_port, DATA2(29) => MUXB_OUT_29_port, 
                           DATA2(28) => MUXB_OUT_28_port, DATA2(27) => 
                           MUXB_OUT_27_port, DATA2(26) => MUXB_OUT_26_port, 
                           DATA2(25) => MUXB_OUT_25_port, DATA2(24) => 
                           MUXB_OUT_24_port, DATA2(23) => MUXB_OUT_23_port, 
                           DATA2(22) => MUXB_OUT_22_port, DATA2(21) => 
                           MUXB_OUT_21_port, DATA2(20) => MUXB_OUT_20_port, 
                           DATA2(19) => MUXB_OUT_19_port, DATA2(18) => 
                           MUXB_OUT_18_port, DATA2(17) => MUXB_OUT_17_port, 
                           DATA2(16) => MUXB_OUT_16_port, DATA2(15) => 
                           MUXB_OUT_15_port, DATA2(14) => MUXB_OUT_14_port, 
                           DATA2(13) => MUXB_OUT_13_port, DATA2(12) => 
                           MUXB_OUT_12_port, DATA2(11) => MUXB_OUT_11_port, 
                           DATA2(10) => MUXB_OUT_10_port, DATA2(9) => 
                           MUXB_OUT_9_port, DATA2(8) => MUXB_OUT_8_port, 
                           DATA2(7) => MUXB_OUT_7_port, DATA2(6) => 
                           MUXB_OUT_6_port, DATA2(5) => MUXB_OUT_5_port, 
                           DATA2(4) => MUXB_OUT_4_port, DATA2(3) => 
                           MUXB_OUT_3_port, DATA2(2) => MUXB_OUT_2_port, 
                           DATA2(1) => MUXB_OUT_1_port, DATA2(0) => 
                           MUXB_OUT_0_port, FUNC(0) => ALU_OPCODE(0), FUNC(1) 
                           => ALU_OPCODE(1), FUNC(2) => ALU_OPCODE(2), FUNC(3) 
                           => ALU_OPCODE(3), FUNC(4) => ALU_OPCODE(4), 
                           OUTALU(31) => ALU_OUT_31_port, OUTALU(30) => 
                           ALU_OUT_30_port, OUTALU(29) => ALU_OUT_29_port, 
                           OUTALU(28) => ALU_OUT_28_port, OUTALU(27) => 
                           ALU_OUT_27_port, OUTALU(26) => ALU_OUT_26_port, 
                           OUTALU(25) => ALU_OUT_25_port, OUTALU(24) => 
                           ALU_OUT_24_port, OUTALU(23) => ALU_OUT_23_port, 
                           OUTALU(22) => ALU_OUT_22_port, OUTALU(21) => 
                           ALU_OUT_21_port, OUTALU(20) => ALU_OUT_20_port, 
                           OUTALU(19) => ALU_OUT_19_port, OUTALU(18) => 
                           ALU_OUT_18_port, OUTALU(17) => ALU_OUT_17_port, 
                           OUTALU(16) => ALU_OUT_16_port, OUTALU(15) => 
                           ALU_OUT_15_port, OUTALU(14) => ALU_OUT_14_port, 
                           OUTALU(13) => ALU_OUT_13_port, OUTALU(12) => 
                           ALU_OUT_12_port, OUTALU(11) => ALU_OUT_11_port, 
                           OUTALU(10) => ALU_OUT_10_port, OUTALU(9) => 
                           ALU_OUT_9_port, OUTALU(8) => ALU_OUT_8_port, 
                           OUTALU(7) => ALU_OUT_7_port, OUTALU(6) => 
                           ALU_OUT_6_port, OUTALU(5) => ALU_OUT_5_port, 
                           OUTALU(4) => ALU_OUT_4_port, OUTALU(3) => 
                           ALU_OUT_3_port, OUTALU(2) => ALU_OUT_2_port, 
                           OUTALU(1) => ALU_OUT_1_port, OUTALU(0) => 
                           ALU_OUT_0_port);
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   U3 : OAI221_X1 port map( B1 => net94215, B2 => n3, C1 => net92960, C2 => n5,
                           A => n6, ZN => MUX_FORWARDING_BRANCH_OUT_9_port);
   U4 : NAND2_X1 port map( A1 => RA_IN_9_port, A2 => n208, ZN => n6);
   U5 : OAI221_X1 port map( B1 => net94215, B2 => n8, C1 => net95433, C2 => n9,
                           A => n10, ZN => MUX_FORWARDING_BRANCH_OUT_8_port);
   U6 : NAND2_X1 port map( A1 => RA_IN_8_port, A2 => n209, ZN => n10);
   U7 : OAI221_X1 port map( B1 => net95422, B2 => n11, C1 => net95411, C2 => 
                           n12, A => n13, ZN => 
                           MUX_FORWARDING_BRANCH_OUT_7_port);
   U8 : NAND2_X1 port map( A1 => RA_IN_7_port, A2 => n208, ZN => n13);
   U9 : OAI221_X1 port map( B1 => net94217, B2 => n14, C1 => net95433, C2 => 
                           n15, A => n16, ZN => 
                           MUX_FORWARDING_BRANCH_OUT_6_port);
   U10 : NAND2_X1 port map( A1 => RA_IN_6_port, A2 => n208, ZN => n16);
   U12 : NAND2_X1 port map( A1 => RA_IN_5_port, A2 => n209, ZN => n19);
   U13 : OAI221_X1 port map( B1 => net95422, B2 => n20, C1 => net95411, C2 => 
                           n21, A => n22, ZN => 
                           MUX_FORWARDING_BRANCH_OUT_4_port);
   U14 : NAND2_X1 port map( A1 => RA_IN_4_port, A2 => n208, ZN => n22);
   U15 : OAI221_X1 port map( B1 => net95422, B2 => n23, C1 => net95411, C2 => 
                           n24, A => n25, ZN => 
                           MUX_FORWARDING_BRANCH_OUT_3_port);
   U16 : NAND2_X1 port map( A1 => RA_IN_3_port, A2 => n208, ZN => n25);
   U17 : OAI221_X1 port map( B1 => net94217, B2 => n26, C1 => net95434, C2 => 
                           n27, A => n28, ZN => 
                           MUX_FORWARDING_BRANCH_OUT_31_port);
   U18 : NAND2_X1 port map( A1 => RA_IN_31_port, A2 => n209, ZN => n28);
   U19 : OAI221_X1 port map( B1 => net95422, B2 => n29, C1 => net95434, C2 => 
                           n30, A => n31, ZN => 
                           MUX_FORWARDING_BRANCH_OUT_30_port);
   U20 : NAND2_X1 port map( A1 => RA_IN_30_port, A2 => n209, ZN => n31);
   U21 : OAI221_X1 port map( B1 => net94215, B2 => n32, C1 => net95434, C2 => 
                           n33, A => n34, ZN => 
                           MUX_FORWARDING_BRANCH_OUT_2_port);
   U22 : NAND2_X1 port map( A1 => RA_IN_2_port, A2 => n209, ZN => n34);
   U23 : OAI221_X1 port map( B1 => net94217, B2 => n35, C1 => net95433, C2 => 
                           n36, A => n37, ZN => 
                           MUX_FORWARDING_BRANCH_OUT_29_port);
   U24 : NAND2_X1 port map( A1 => RA_IN_29_port, A2 => n209, ZN => n37);
   U25 : OAI221_X1 port map( B1 => net94217, B2 => n38, C1 => net92959, C2 => 
                           n39, A => n40, ZN => 
                           MUX_FORWARDING_BRANCH_OUT_28_port);
   U26 : NAND2_X1 port map( A1 => RA_IN_28_port, A2 => n7, ZN => n40);
   U28 : NAND2_X1 port map( A1 => RA_IN_27_port, A2 => n208, ZN => n43);
   U29 : OAI221_X1 port map( B1 => net95422, B2 => n44, C1 => net95411, C2 => 
                           n45, A => n46, ZN => 
                           MUX_FORWARDING_BRANCH_OUT_26_port);
   U30 : NAND2_X1 port map( A1 => RA_IN_26_port, A2 => n7, ZN => n46);
   U31 : OAI221_X1 port map( B1 => net95422, B2 => n47, C1 => net95411, C2 => 
                           n48, A => n49, ZN => 
                           MUX_FORWARDING_BRANCH_OUT_25_port);
   U32 : NAND2_X1 port map( A1 => RA_IN_25_port, A2 => n7, ZN => n49);
   U33 : OAI221_X1 port map( B1 => net94215, B2 => n50, C1 => net95411, C2 => 
                           n51, A => n52, ZN => 
                           MUX_FORWARDING_BRANCH_OUT_24_port);
   U34 : NAND2_X1 port map( A1 => RA_IN_24_port, A2 => n7, ZN => n52);
   U35 : OAI221_X1 port map( B1 => net94215, B2 => n53, C1 => net95411, C2 => 
                           n54, A => n55, ZN => 
                           MUX_FORWARDING_BRANCH_OUT_23_port);
   U36 : NAND2_X1 port map( A1 => RA_IN_23_port, A2 => n208, ZN => n55);
   U37 : OAI221_X1 port map( B1 => net94215, B2 => n56, C1 => net95411, C2 => 
                           n57, A => n58, ZN => 
                           MUX_FORWARDING_BRANCH_OUT_22_port);
   U38 : NAND2_X1 port map( A1 => RA_IN_22_port, A2 => n7, ZN => n58);
   U39 : OAI221_X1 port map( B1 => net94217, B2 => n59, C1 => net92960, C2 => 
                           n60, A => n61, ZN => 
                           MUX_FORWARDING_BRANCH_OUT_21_port);
   U40 : NAND2_X1 port map( A1 => RA_IN_21_port, A2 => n7, ZN => n61);
   U41 : OAI221_X1 port map( B1 => net94217, B2 => n62, C1 => net92959, C2 => 
                           n63, A => n64, ZN => 
                           MUX_FORWARDING_BRANCH_OUT_20_port);
   U42 : NAND2_X1 port map( A1 => RA_IN_20_port, A2 => n209, ZN => n64);
   U44 : NAND2_X1 port map( A1 => RA_IN_1_port, A2 => n7, ZN => n67);
   U45 : OAI221_X1 port map( B1 => net95422, B2 => n68, C1 => net92960, C2 => 
                           n69, A => n70, ZN => 
                           MUX_FORWARDING_BRANCH_OUT_19_port);
   U46 : NAND2_X1 port map( A1 => RA_IN_19_port, A2 => n208, ZN => n70);
   U47 : OAI221_X1 port map( B1 => net94217, B2 => n71, C1 => net92960, C2 => 
                           n72, A => n73, ZN => 
                           MUX_FORWARDING_BRANCH_OUT_18_port);
   U48 : NAND2_X1 port map( A1 => RA_IN_18_port, A2 => n7, ZN => n73);
   U49 : OAI221_X1 port map( B1 => net94217, B2 => n74, C1 => net92959, C2 => 
                           n75, A => n76, ZN => 
                           MUX_FORWARDING_BRANCH_OUT_17_port);
   U50 : NAND2_X1 port map( A1 => RA_IN_17_port, A2 => n208, ZN => n76);
   U52 : NAND2_X1 port map( A1 => RA_IN_16_port, A2 => n7, ZN => n79);
   U53 : OAI221_X1 port map( B1 => net95422, B2 => n80, C1 => net95411, C2 => 
                           n81, A => n82, ZN => 
                           MUX_FORWARDING_BRANCH_OUT_15_port);
   U54 : NAND2_X1 port map( A1 => RA_IN_15_port, A2 => n209, ZN => n82);
   U55 : OAI221_X1 port map( B1 => net94217, B2 => n83, C1 => net95433, C2 => 
                           n84, A => n85, ZN => 
                           MUX_FORWARDING_BRANCH_OUT_14_port);
   U56 : NAND2_X1 port map( A1 => RA_IN_14_port, A2 => n208, ZN => n85);
   U57 : OAI221_X1 port map( B1 => net94217, B2 => n86, C1 => net92959, C2 => 
                           n87, A => n88, ZN => 
                           MUX_FORWARDING_BRANCH_OUT_13_port);
   U58 : NAND2_X1 port map( A1 => RA_IN_13_port, A2 => n7, ZN => n88);
   U60 : NAND2_X1 port map( A1 => RA_IN_12_port, A2 => n209, ZN => n91);
   U61 : OAI221_X1 port map( B1 => net95422, B2 => n92, C1 => net95411, C2 => 
                           n93, A => n94, ZN => 
                           MUX_FORWARDING_BRANCH_OUT_11_port);
   U62 : NAND2_X1 port map( A1 => RA_IN_11_port, A2 => n7, ZN => n94);
   U63 : OAI221_X1 port map( B1 => net95422, B2 => n95, C1 => net95434, C2 => 
                           n96, A => n97, ZN => 
                           MUX_FORWARDING_BRANCH_OUT_10_port);
   U64 : NAND2_X1 port map( A1 => RA_IN_10_port, A2 => n209, ZN => n97);
   U66 : NAND2_X1 port map( A1 => RA_IN_0_port, A2 => n209, ZN => n100);
   U68 : NAND2_X1 port map( A1 => n210, A2 => n101, ZN => n4);
   U70 : INV_X1 port map( A => ForwardD_1_port, ZN => n101);
   U71 : OAI221_X1 port map( B1 => n3, B2 => net95343, C1 => n5, C2 => net95310
                           , A => n104, ZN => ALU_inputB_9_port);
   U72 : NAND2_X1 port map( A1 => RB_OUT_9_port, A2 => n103, ZN => n104);
   U73 : OAI221_X1 port map( B1 => n8, B2 => n185, C1 => n9, C2 => net95310, A 
                           => n106, ZN => ALU_inputB_8_port);
   U74 : NAND2_X1 port map( A1 => RB_OUT_8_port, A2 => n103, ZN => n106);
   U75 : OAI221_X1 port map( B1 => n11, B2 => n184, C1 => n12, C2 => net95310, 
                           A => n107, ZN => ALU_inputB_7_port);
   U76 : NAND2_X1 port map( A1 => RB_OUT_7_port, A2 => n175, ZN => n107);
   U77 : OAI221_X1 port map( B1 => n14, B2 => n184, C1 => n15, C2 => net95310, 
                           A => n108, ZN => ALU_inputB_6_port);
   U78 : NAND2_X1 port map( A1 => RB_OUT_6_port, A2 => n176, ZN => n108);
   U79 : OAI221_X1 port map( B1 => n17, B2 => n184, C1 => n18, C2 => net95310, 
                           A => n109, ZN => ALU_inputB_5_port);
   U80 : NAND2_X1 port map( A1 => RB_OUT_5_port, A2 => n181, ZN => n109);
   U81 : OAI221_X1 port map( B1 => n20, B2 => net95343, C1 => n21, C2 => 
                           net95310, A => n110, ZN => ALU_inputB_4_port);
   U82 : NAND2_X1 port map( A1 => RB_OUT_4_port, A2 => n181, ZN => n110);
   U83 : OAI221_X1 port map( B1 => n23, B2 => n183, C1 => n24, C2 => net95311, 
                           A => n111, ZN => ALU_inputB_3_port);
   U84 : NAND2_X1 port map( A1 => RB_OUT_3_port, A2 => n102, ZN => n111);
   U85 : OAI221_X1 port map( B1 => n26, B2 => net95343, C1 => n27, C2 => 
                           net95310, A => n112, ZN => ALU_inputB_31_port);
   U86 : NAND2_X1 port map( A1 => RB_OUT_31_port, A2 => n178, ZN => n112);
   U87 : OAI221_X1 port map( B1 => n29, B2 => n184, C1 => n30, C2 => net95311, 
                           A => n113, ZN => ALU_inputB_30_port);
   U88 : NAND2_X1 port map( A1 => RB_OUT_30_port, A2 => n179, ZN => n113);
   U89 : OAI221_X1 port map( B1 => n32, B2 => net95343, C1 => n33, C2 => 
                           net95310, A => n114, ZN => ALU_inputB_2_port);
   U90 : NAND2_X1 port map( A1 => RB_OUT_2_port, A2 => n179, ZN => n114);
   U91 : OAI221_X1 port map( B1 => n35, B2 => n185, C1 => n36, C2 => net95311, 
                           A => n115, ZN => ALU_inputB_29_port);
   U92 : NAND2_X1 port map( A1 => RB_OUT_29_port, A2 => n177, ZN => n115);
   U93 : OAI221_X1 port map( B1 => n38, B2 => n184, C1 => n39, C2 => net95311, 
                           A => n116, ZN => ALU_inputB_28_port);
   U94 : NAND2_X1 port map( A1 => RB_OUT_28_port, A2 => n177, ZN => n116);
   U95 : OAI221_X1 port map( B1 => n41, B2 => net95343, C1 => n42, C2 => 
                           net95310, A => n117, ZN => ALU_inputB_27_port);
   U96 : NAND2_X1 port map( A1 => RB_OUT_27_port, A2 => n105, ZN => n117);
   U97 : OAI221_X1 port map( B1 => n44, B2 => net95343, C1 => n45, C2 => 
                           net95310, A => n118, ZN => ALU_inputB_26_port);
   U98 : NAND2_X1 port map( A1 => RB_OUT_26_port, A2 => n176, ZN => n118);
   U99 : OAI221_X1 port map( B1 => n47, B2 => n184, C1 => n48, C2 => net95311, 
                           A => n119, ZN => ALU_inputB_25_port);
   U100 : NAND2_X1 port map( A1 => RB_OUT_25_port, A2 => n175, ZN => n119);
   U101 : OAI221_X1 port map( B1 => n50, B2 => n185, C1 => n51, C2 => net95310,
                           A => n120, ZN => ALU_inputB_24_port);
   U102 : NAND2_X1 port map( A1 => RB_OUT_24_port, A2 => n177, ZN => n120);
   U103 : OAI221_X1 port map( B1 => n53, B2 => net95343, C1 => n54, C2 => 
                           net95311, A => n121, ZN => ALU_inputB_23_port);
   U104 : NAND2_X1 port map( A1 => RB_OUT_23_port, A2 => n180, ZN => n121);
   U105 : OAI221_X1 port map( B1 => n56, B2 => n184, C1 => n57, C2 => net95311,
                           A => n122, ZN => ALU_inputB_22_port);
   U106 : NAND2_X1 port map( A1 => RB_OUT_22_port, A2 => n180, ZN => n122);
   U107 : OAI221_X1 port map( B1 => n59, B2 => net95343, C1 => n60, C2 => 
                           net95310, A => n123, ZN => ALU_inputB_21_port);
   U108 : NAND2_X1 port map( A1 => RB_OUT_21_port, A2 => n174, ZN => n123);
   U109 : OAI221_X1 port map( B1 => n62, B2 => n184, C1 => n63, C2 => net95310,
                           A => n124, ZN => ALU_inputB_20_port);
   U110 : NAND2_X1 port map( A1 => RB_OUT_20_port, A2 => n103, ZN => n124);
   U111 : OAI221_X1 port map( B1 => n65, B2 => net95343, C1 => n66, C2 => 
                           net95311, A => n125, ZN => ALU_inputB_1_port);
   U112 : NAND2_X1 port map( A1 => RB_OUT_1_port, A2 => n175, ZN => n125);
   U113 : OAI221_X1 port map( B1 => n68, B2 => net95343, C1 => n69, C2 => 
                           net95310, A => n126, ZN => ALU_inputB_19_port);
   U114 : NAND2_X1 port map( A1 => RB_OUT_19_port, A2 => n102, ZN => n126);
   U115 : OAI221_X1 port map( B1 => n71, B2 => n185, C1 => n72, C2 => net95310,
                           A => n127, ZN => ALU_inputB_18_port);
   U116 : NAND2_X1 port map( A1 => RB_OUT_18_port, A2 => n174, ZN => n127);
   U117 : OAI221_X1 port map( B1 => n74, B2 => n185, C1 => n75, C2 => net95310,
                           A => n128, ZN => ALU_inputB_17_port);
   U118 : NAND2_X1 port map( A1 => RB_OUT_17_port, A2 => n105, ZN => n128);
   U119 : OAI221_X1 port map( B1 => n77, B2 => n185, C1 => n78, C2 => net95310,
                           A => n129, ZN => ALU_inputB_16_port);
   U120 : NAND2_X1 port map( A1 => RB_OUT_16_port, A2 => n176, ZN => n129);
   U121 : OAI221_X1 port map( B1 => n80, B2 => net95343, C1 => n81, C2 => 
                           net95310, A => n130, ZN => ALU_inputB_15_port);
   U122 : NAND2_X1 port map( A1 => RB_OUT_15_port, A2 => n102, ZN => n130);
   U123 : OAI221_X1 port map( B1 => n83, B2 => net95343, C1 => n84, C2 => 
                           net95310, A => n131, ZN => ALU_inputB_14_port);
   U124 : NAND2_X1 port map( A1 => RB_OUT_14_port, A2 => n179, ZN => n131);
   U125 : OAI221_X1 port map( B1 => n86, B2 => net95343, C1 => n87, C2 => 
                           net95311, A => n132, ZN => ALU_inputB_13_port);
   U126 : NAND2_X1 port map( A1 => RB_OUT_13_port, A2 => n174, ZN => n132);
   U127 : OAI221_X1 port map( B1 => n89, B2 => net95343, C1 => n90, C2 => 
                           net95310, A => n133, ZN => ALU_inputB_12_port);
   U128 : NAND2_X1 port map( A1 => RB_OUT_12_port, A2 => n105, ZN => n133);
   U129 : OAI221_X1 port map( B1 => n92, B2 => net95343, C1 => n93, C2 => 
                           net95310, A => n134, ZN => ALU_inputB_11_port);
   U130 : NAND2_X1 port map( A1 => RB_OUT_11_port, A2 => n178, ZN => n134);
   U131 : OAI221_X1 port map( B1 => n95, B2 => n185, C1 => n96, C2 => net95311,
                           A => n135, ZN => ALU_inputB_10_port);
   U132 : NAND2_X1 port map( A1 => RB_OUT_10_port, A2 => n178, ZN => n135);
   U140 : NAND2_X1 port map( A1 => RA_OUT_9_port, A2 => n141, ZN => n140);
   U141 : INV_X1 port map( A => MUXC_OUT_9_port, ZN => n5);
   U142 : INV_X1 port map( A => ADDR_DRAM_9_port, ZN => n3);
   U144 : NAND2_X1 port map( A1 => RA_OUT_8_port, A2 => n141, ZN => n142);
   U145 : INV_X1 port map( A => MUXC_OUT_8_port, ZN => n9);
   U146 : INV_X1 port map( A => ADDR_DRAM_8_port, ZN => n8);
   U148 : NAND2_X1 port map( A1 => RA_OUT_7_port, A2 => n141, ZN => n143);
   U149 : INV_X1 port map( A => MUXC_OUT_7_port, ZN => n12);
   U150 : INV_X1 port map( A => ADDR_DRAM_7_port, ZN => n11);
   U152 : NAND2_X1 port map( A1 => RA_OUT_6_port, A2 => n141, ZN => n144);
   U153 : INV_X1 port map( A => MUXC_OUT_6_port, ZN => n15);
   U154 : INV_X1 port map( A => ADDR_DRAM_6_port, ZN => n14);
   U156 : NAND2_X1 port map( A1 => RA_OUT_5_port, A2 => n141, ZN => n145);
   U157 : INV_X1 port map( A => MUXC_OUT_5_port, ZN => n18);
   U158 : INV_X1 port map( A => ADDR_DRAM_5_port, ZN => n17);
   U160 : NAND2_X1 port map( A1 => RA_OUT_4_port, A2 => n141, ZN => n146);
   U161 : INV_X1 port map( A => MUXC_OUT_4_port, ZN => n21);
   U162 : INV_X1 port map( A => ADDR_DRAM_4_port, ZN => n20);
   U164 : NAND2_X1 port map( A1 => RA_OUT_3_port, A2 => n141, ZN => n147);
   U165 : INV_X1 port map( A => MUXC_OUT_3_port, ZN => n24);
   U166 : INV_X1 port map( A => ADDR_DRAM_3_port, ZN => n23);
   U168 : NAND2_X1 port map( A1 => RA_OUT_31_port, A2 => n141, ZN => n148);
   U169 : INV_X1 port map( A => MUXC_OUT_31_port, ZN => n27);
   U170 : INV_X1 port map( A => ADDR_DRAM_31_port, ZN => n26);
   U171 : OAI221_X1 port map( B1 => n29, B2 => n138, C1 => n30, C2 => n139, A 
                           => n149, ZN => ALU_inputA_30_port);
   U172 : NAND2_X1 port map( A1 => RA_OUT_30_port, A2 => n141, ZN => n149);
   U173 : INV_X1 port map( A => MUXC_OUT_30_port, ZN => n30);
   U174 : INV_X1 port map( A => ADDR_DRAM_30_port, ZN => n29);
   U176 : NAND2_X1 port map( A1 => RA_OUT_2_port, A2 => n141, ZN => n150);
   U177 : INV_X1 port map( A => MUXC_OUT_2_port, ZN => n33);
   U178 : INV_X1 port map( A => ADDR_DRAM_2_port, ZN => n32);
   U180 : NAND2_X1 port map( A1 => RA_OUT_29_port, A2 => n141, ZN => n151);
   U181 : INV_X1 port map( A => MUXC_OUT_29_port, ZN => n36);
   U182 : INV_X1 port map( A => ADDR_DRAM_29_port, ZN => n35);
   U183 : OAI221_X1 port map( B1 => n38, B2 => n138, C1 => n39, C2 => n139, A 
                           => n152, ZN => ALU_inputA_28_port);
   U184 : NAND2_X1 port map( A1 => RA_OUT_28_port, A2 => n141, ZN => n152);
   U185 : INV_X1 port map( A => MUXC_OUT_28_port, ZN => n39);
   U186 : INV_X1 port map( A => ADDR_DRAM_28_port, ZN => n38);
   U187 : OAI221_X1 port map( B1 => n41, B2 => n138, C1 => n42, C2 => n139, A 
                           => n153, ZN => ALU_inputA_27_port);
   U188 : NAND2_X1 port map( A1 => RA_OUT_27_port, A2 => n141, ZN => n153);
   U189 : INV_X1 port map( A => MUXC_OUT_27_port, ZN => n42);
   U190 : INV_X1 port map( A => ADDR_DRAM_27_port, ZN => n41);
   U192 : NAND2_X1 port map( A1 => RA_OUT_26_port, A2 => n141, ZN => n154);
   U193 : INV_X1 port map( A => MUXC_OUT_26_port, ZN => n45);
   U194 : INV_X1 port map( A => ADDR_DRAM_26_port, ZN => n44);
   U196 : NAND2_X1 port map( A1 => RA_OUT_25_port, A2 => n141, ZN => n155);
   U197 : INV_X1 port map( A => MUXC_OUT_25_port, ZN => n48);
   U198 : INV_X1 port map( A => ADDR_DRAM_25_port, ZN => n47);
   U200 : NAND2_X1 port map( A1 => RA_OUT_24_port, A2 => n141, ZN => n156);
   U201 : INV_X1 port map( A => MUXC_OUT_24_port, ZN => n51);
   U202 : INV_X1 port map( A => ADDR_DRAM_24_port, ZN => n50);
   U204 : NAND2_X1 port map( A1 => RA_OUT_23_port, A2 => n141, ZN => n157);
   U205 : INV_X1 port map( A => MUXC_OUT_23_port, ZN => n54);
   U206 : INV_X1 port map( A => ADDR_DRAM_23_port, ZN => n53);
   U208 : NAND2_X1 port map( A1 => RA_OUT_22_port, A2 => n141, ZN => n158);
   U209 : INV_X1 port map( A => MUXC_OUT_22_port, ZN => n57);
   U210 : INV_X1 port map( A => ADDR_DRAM_22_port, ZN => n56);
   U212 : NAND2_X1 port map( A1 => RA_OUT_21_port, A2 => n141, ZN => n159);
   U213 : INV_X1 port map( A => MUXC_OUT_21_port, ZN => n60);
   U214 : INV_X1 port map( A => ADDR_DRAM_21_port, ZN => n59);
   U216 : NAND2_X1 port map( A1 => RA_OUT_20_port, A2 => n141, ZN => n160);
   U217 : INV_X1 port map( A => MUXC_OUT_20_port, ZN => n63);
   U218 : INV_X1 port map( A => ADDR_DRAM_20_port, ZN => n62);
   U220 : NAND2_X1 port map( A1 => RA_OUT_1_port, A2 => n141, ZN => n161);
   U221 : INV_X1 port map( A => MUXC_OUT_1_port, ZN => n66);
   U222 : INV_X1 port map( A => ADDR_DRAM_1_port, ZN => n65);
   U224 : NAND2_X1 port map( A1 => RA_OUT_19_port, A2 => n141, ZN => n162);
   U225 : INV_X1 port map( A => MUXC_OUT_19_port, ZN => n69);
   U226 : INV_X1 port map( A => ADDR_DRAM_19_port, ZN => n68);
   U228 : NAND2_X1 port map( A1 => RA_OUT_18_port, A2 => n141, ZN => n163);
   U229 : INV_X1 port map( A => MUXC_OUT_18_port, ZN => n72);
   U230 : INV_X1 port map( A => ADDR_DRAM_18_port, ZN => n71);
   U232 : NAND2_X1 port map( A1 => RA_OUT_17_port, A2 => n141, ZN => n164);
   U233 : INV_X1 port map( A => MUXC_OUT_17_port, ZN => n75);
   U234 : INV_X1 port map( A => ADDR_DRAM_17_port, ZN => n74);
   U236 : NAND2_X1 port map( A1 => RA_OUT_16_port, A2 => n141, ZN => n165);
   U237 : INV_X1 port map( A => MUXC_OUT_16_port, ZN => n78);
   U238 : INV_X1 port map( A => ADDR_DRAM_16_port, ZN => n77);
   U240 : NAND2_X1 port map( A1 => RA_OUT_15_port, A2 => n141, ZN => n166);
   U241 : INV_X1 port map( A => MUXC_OUT_15_port, ZN => n81);
   U242 : INV_X1 port map( A => ADDR_DRAM_15_port, ZN => n80);
   U244 : NAND2_X1 port map( A1 => RA_OUT_14_port, A2 => n141, ZN => n167);
   U245 : INV_X1 port map( A => MUXC_OUT_14_port, ZN => n84);
   U246 : INV_X1 port map( A => ADDR_DRAM_14_port, ZN => n83);
   U248 : NAND2_X1 port map( A1 => RA_OUT_13_port, A2 => n141, ZN => n168);
   U249 : INV_X1 port map( A => MUXC_OUT_13_port, ZN => n87);
   U250 : INV_X1 port map( A => ADDR_DRAM_13_port, ZN => n86);
   U252 : NAND2_X1 port map( A1 => RA_OUT_12_port, A2 => n141, ZN => n169);
   U253 : INV_X1 port map( A => MUXC_OUT_12_port, ZN => n90);
   U254 : INV_X1 port map( A => ADDR_DRAM_12_port, ZN => n89);
   U256 : NAND2_X1 port map( A1 => RA_OUT_11_port, A2 => n141, ZN => n170);
   U257 : INV_X1 port map( A => MUXC_OUT_11_port, ZN => n93);
   U258 : INV_X1 port map( A => ADDR_DRAM_11_port, ZN => n92);
   U260 : NAND2_X1 port map( A1 => RA_OUT_10_port, A2 => n141, ZN => n171);
   U261 : INV_X1 port map( A => MUXC_OUT_10_port, ZN => n96);
   U262 : INV_X1 port map( A => ADDR_DRAM_10_port, ZN => n95);
   U264 : NAND2_X1 port map( A1 => RA_OUT_0_port, A2 => n141, ZN => n172);
   U267 : INV_X1 port map( A => MUXC_OUT_0_port, ZN => n99);
   U269 : INV_X1 port map( A => ForwardA_1_port, ZN => n173);
   U65 : OAI221_X1 port map( B1 => net94217, B2 => n98, C1 => net95434, C2 => 
                           n99, A => n100, ZN => 
                           MUX_FORWARDING_BRANCH_OUT_0_port);
   U270 : INV_X1 port map( A => ADDR_DRAM_0_port, ZN => n98);
   U138 : INV_X1 port map( A => forwardB_1_port, ZN => n137);
   U11 : BUF_X1 port map( A => forwardB_1_port, Z => n1);
   U27 : INV_X1 port map( A => net95415, ZN => n102);
   U43 : INV_X1 port map( A => net95415, ZN => n103);
   U51 : INV_X1 port map( A => net95415, ZN => n105);
   U59 : INV_X1 port map( A => net95415, ZN => n174);
   U67 : INV_X1 port map( A => net95415, ZN => n175);
   U69 : INV_X1 port map( A => net95415, ZN => n176);
   U133 : INV_X1 port map( A => net95415, ZN => n177);
   U134 : INV_X1 port map( A => net95415, ZN => n178);
   U135 : BUF_X1 port map( A => net95551, Z => n179);
   U136 : BUF_X1 port map( A => net95252, Z => n180);
   U137 : BUF_X1 port map( A => net95253, Z => n181);
   U139 : INV_X1 port map( A => net95415, ZN => net95252);
   U143 : INV_X1 port map( A => net95342, ZN => n182);
   U147 : INV_X1 port map( A => n182, ZN => n183);
   U151 : INV_X1 port map( A => n182, ZN => n185);
   U155 : INV_X1 port map( A => n182, ZN => n184);
   U159 : CLKBUF_X1 port map( A => ALU_inputA_30_port, Z => n186);
   U163 : OAI221_X4 port map( B1 => n35, B2 => n138, C1 => n36, C2 => n139, A 
                           => n151, ZN => ALU_inputA_29_port);
   U167 : OAI221_X4 port map( B1 => n65, B2 => n138, C1 => n66, C2 => n139, A 
                           => n161, ZN => ALU_inputA_1_port);
   U175 : OAI221_X4 port map( B1 => n17, B2 => n138, C1 => n18, C2 => n139, A 
                           => n145, ZN => ALU_inputA_5_port);
   U179 : OAI221_X4 port map( B1 => n26, B2 => n138, C1 => n27, C2 => n139, A 
                           => n148, ZN => ALU_inputA_31_port);
   U203 : OAI221_X4 port map( B1 => n53, B2 => n138, C1 => n54, C2 => n139, A 
                           => n157, ZN => ALU_inputA_23_port);
   U207 : OAI221_X4 port map( B1 => n71, B2 => n138, C1 => n72, C2 => n139, A 
                           => n163, ZN => ALU_inputA_18_port);
   U211 : OAI221_X4 port map( B1 => n74, B2 => n138, C1 => n75, C2 => n139, A 
                           => n164, ZN => ALU_inputA_17_port);
   U215 : OAI221_X4 port map( B1 => n68, B2 => n138, C1 => n69, C2 => n139, A 
                           => n162, ZN => ALU_inputA_19_port);
   U219 : OAI221_X4 port map( B1 => n62, B2 => n138, C1 => n63, C2 => n139, A 
                           => n160, ZN => ALU_inputA_20_port);
   U223 : OAI221_X4 port map( B1 => n3, B2 => n138, C1 => n5, C2 => n139, A => 
                           n140, ZN => ALU_inputA_9_port);
   U227 : OAI221_X4 port map( B1 => n89, B2 => n138, C1 => n90, C2 => n139, A 
                           => n169, ZN => ALU_inputA_12_port);
   U231 : OAI221_X4 port map( B1 => n8, B2 => n138, C1 => n9, C2 => n139, A => 
                           n142, ZN => ALU_inputA_8_port);
   U235 : OAI221_X4 port map( B1 => n95, B2 => n138, C1 => n96, C2 => n139, A 
                           => n171, ZN => ALU_inputA_10_port);
   U239 : OAI221_X4 port map( B1 => n14, B2 => n138, C1 => n15, C2 => n139, A 
                           => n144, ZN => ALU_inputA_6_port);
   U243 : OAI221_X4 port map( B1 => n83, B2 => n138, C1 => n84, C2 => n139, A 
                           => n167, ZN => ALU_inputA_14_port);
   U247 : OAI221_X4 port map( B1 => n20, B2 => n138, C1 => n21, C2 => n139, A 
                           => n146, ZN => ALU_inputA_4_port);
   U251 : OAI221_X4 port map( B1 => n32, B2 => n138, C1 => n33, C2 => n139, A 
                           => n150, ZN => ALU_inputA_2_port);
   U255 : OAI221_X4 port map( B1 => n59, B2 => n138, C1 => n60, C2 => n139, A 
                           => n159, ZN => ALU_inputA_21_port);
   U259 : OAI221_X4 port map( B1 => n77, B2 => n138, C1 => n78, C2 => n139, A 
                           => n165, ZN => ALU_inputA_16_port);
   U263 : OAI221_X4 port map( B1 => n56, B2 => n138, C1 => n57, C2 => n139, A 
                           => n158, ZN => ALU_inputA_22_port);
   U265 : OAI221_X4 port map( B1 => n11, B2 => n138, C1 => n12, C2 => n139, A 
                           => n143, ZN => ALU_inputA_7_port);
   U266 : OAI221_X4 port map( B1 => n86, B2 => n138, C1 => n87, C2 => n139, A 
                           => n168, ZN => ALU_inputA_13_port);
   U268 : OR2_X2 port map( A1 => n1, A2 => forwardB_0_port, ZN => net95415);
   U271 : INV_X1 port map( A => net95521, ZN => n187);
   U272 : INV_X1 port map( A => n98, ZN => n188);
   U273 : NAND2_X1 port map( A1 => n187, A2 => n191, ZN => n189);
   U274 : NAND2_X1 port map( A1 => n193, A2 => n188, ZN => n190);
   U275 : AND2_X1 port map( A1 => forwardB_0_port, A2 => n137, ZN => n191);
   U276 : NAND2_X1 port map( A1 => n192, A2 => n189, ZN => ALU_inputB_0_port);
   U277 : AND2_X1 port map( A1 => n190, A2 => n136, ZN => n192);
   U278 : NOR2_X1 port map( A1 => n137, A2 => forwardB_0_port, ZN => n193);
   U279 : OR3_X1 port map( A1 => forwardB_0_port, A2 => n1, A3 => n194, ZN => 
                           n136);
   U280 : INV_X1 port map( A => RB_OUT_0_port, ZN => n194);
   U281 : INV_X1 port map( A => MUXC_OUT_0_port, ZN => net95521);
   U282 : OR2_X1 port map( A1 => n137, A2 => forwardB_0_port, ZN => net95342);
   U283 : OR2_X1 port map( A1 => n137, A2 => net95416, ZN => net95343);
   U284 : OAI221_X4 port map( B1 => n98, B2 => n138, C1 => n99, C2 => n139, A 
                           => n172, ZN => ALU_inputA_0_port);
   U285 : INV_X2 port map( A => n191, ZN => net95310);
   U286 : INV_X1 port map( A => n191, ZN => net95311);
   U287 : CLKBUF_X2 port map( A => n4, Z => net95411);
   U288 : OAI221_X4 port map( B1 => n23, B2 => n138, C1 => n24, C2 => n139, A 
                           => n147, ZN => ALU_inputA_3_port);
   U289 : OAI221_X4 port map( B1 => net94215, B2 => n17, C1 => net95433, C2 => 
                           n18, A => n19, ZN => 
                           MUX_FORWARDING_BRANCH_OUT_5_port);
   U290 : OAI221_X4 port map( B1 => n80, B2 => n138, C1 => n81, C2 => n139, A 
                           => n166, ZN => ALU_inputA_15_port);
   U291 : CLKBUF_X1 port map( A => MUX_IMM_OUT_16_port, Z => n195);
   U292 : INV_X1 port map( A => net95415, ZN => net95551);
   U293 : CLKBUF_X1 port map( A => RD2_OUT_4_port, Z => n196);
   U294 : CLKBUF_X1 port map( A => RD2_OUT_2_port, Z => n197);
   U295 : CLKBUF_X1 port map( A => RD2_OUT_1_port, Z => n198);
   U296 : CLKBUF_X1 port map( A => RD2_OUT_0_port, Z => n199);
   U297 : CLKBUF_X1 port map( A => RD3_OUT_4_port, Z => n200);
   U298 : CLKBUF_X1 port map( A => RD3_OUT_3_port, Z => n201);
   U299 : CLKBUF_X1 port map( A => RD3_OUT_0_port, Z => n202);
   U300 : CLKBUF_X1 port map( A => RD2_OUT_3_port, Z => n203);
   U301 : INV_X2 port map( A => net94214, ZN => net94215);
   U302 : INV_X1 port map( A => net92958, ZN => net95434);
   U303 : INV_X1 port map( A => net92958, ZN => net95433);
   U304 : INV_X1 port map( A => net92958, ZN => net92960);
   U305 : CLKBUF_X3 port map( A => n2, Z => net95422);
   U306 : CLKBUF_X1 port map( A => MUX_FORWARDING_BRANCH_OUT_10_port, Z => n204
                           );
   U307 : OAI221_X1 port map( B1 => net94215, B2 => n89, C1 => net95411, C2 => 
                           n90, A => n91, ZN => 
                           MUX_FORWARDING_BRANCH_OUT_12_port);
   U308 : OAI221_X1 port map( B1 => net95422, B2 => n41, C1 => net95411, C2 => 
                           n42, A => n43, ZN => 
                           MUX_FORWARDING_BRANCH_OUT_27_port);
   U309 : OAI221_X1 port map( B1 => net95422, B2 => n65, C1 => net95411, C2 => 
                           n66, A => n67, ZN => 
                           MUX_FORWARDING_BRANCH_OUT_1_port);
   U310 : CLKBUF_X1 port map( A => forwardB_0_port, Z => net95416);
   U311 : BUF_X4 port map( A => n214, Z => BRANCH_ALU_OUT(30));
   U312 : BUF_X4 port map( A => n215, Z => BRANCH_ALU_OUT(25));
   U313 : BUF_X1 port map( A => MUX_FORWARDING_BRANCH_OUT_3_port, Z => n205);
   U315 : OR2_X4 port map( A1 => n173, A2 => ForwardA_0_port, ZN => n138);
   U316 : OAI221_X4 port map( B1 => n92, B2 => n138, C1 => n93, C2 => n139, A 
                           => n170, ZN => ALU_inputA_11_port);
   U317 : NAND2_X4 port map( A1 => ForwardA_0_port, A2 => n173, ZN => n139);
   U318 : BUF_X2 port map( A => n216, Z => BRANCH_ALU_OUT(23));
   U319 : NOR2_X1 port map( A1 => ForwardD_0_port, A2 => n217, ZN => n208);
   U320 : NOR2_X1 port map( A1 => ForwardD_0_port, A2 => n217, ZN => n209);
   U321 : NOR2_X1 port map( A1 => ForwardD_0_port, A2 => ForwardD_1_port, ZN =>
                           n7);
   U322 : NOR2_X4 port map( A1 => ForwardA_0_port, A2 => ForwardA_1_port, ZN =>
                           n141);
   U323 : CLKBUF_X1 port map( A => ForwardD_0_port, Z => n210);
   U324 : OR2_X1 port map( A1 => n101, A2 => ForwardD_0_port, ZN => n2);
   U325 : INV_X1 port map( A => net95415, ZN => net95253);
   U326 : INV_X1 port map( A => n2, ZN => net94214);
   U327 : INV_X2 port map( A => net94214, ZN => net94217);
   U328 : OAI221_X1 port map( B1 => net95422, B2 => n77, C1 => net92960, C2 => 
                           n78, A => n79, ZN => 
                           MUX_FORWARDING_BRANCH_OUT_16_port);
   U329 : INV_X1 port map( A => n4, ZN => net92958);
   U330 : INV_X1 port map( A => net92958, ZN => net92959);
   reg_file_0 : register_file_NUMBIT32_BITADDR5 port map( CLK => CLK, RESET => 
                           RST, ENABLE => REGF_LATCH_EN, RD1 => RFR1_EN, RD2 =>
                           RFR2_EN, WR => RF_WE, ADD_WR(4) => 
                           MUX_WRaddr_OUT_4_port, ADD_WR(3) => 
                           MUX_WRaddr_OUT_3_port, ADD_WR(2) => 
                           MUX_WRaddr_OUT_2_port, ADD_WR(1) => 
                           MUX_WRaddr_OUT_1_port, ADD_WR(0) => 
                           MUX_WRaddr_OUT_0_port, ADD_RD1(4) => RS1(4), 
                           ADD_RD1(3) => RS1(3), ADD_RD1(2) => RS1(2), 
                           ADD_RD1(1) => RS1(1), ADD_RD1(0) => RS1(0), 
                           ADD_RD2(4) => RS2(4), ADD_RD2(3) => RS2(3), 
                           ADD_RD2(2) => RS2(2), ADD_RD2(1) => RS2(1), 
                           ADD_RD2(0) => RS2(0), DATAIN(31) => 
                           MUX_WRdata_OUT_31_port, DATAIN(30) => 
                           MUX_WRdata_OUT_30_port, DATAIN(29) => 
                           MUX_WRdata_OUT_29_port, DATAIN(28) => 
                           MUX_WRdata_OUT_28_port, DATAIN(27) => 
                           MUX_WRdata_OUT_27_port, DATAIN(26) => 
                           MUX_WRdata_OUT_26_port, DATAIN(25) => 
                           MUX_WRdata_OUT_25_port, DATAIN(24) => 
                           MUX_WRdata_OUT_24_port, DATAIN(23) => 
                           MUX_WRdata_OUT_23_port, DATAIN(22) => 
                           MUX_WRdata_OUT_22_port, DATAIN(21) => 
                           MUX_WRdata_OUT_21_port, DATAIN(20) => 
                           MUX_WRdata_OUT_20_port, DATAIN(19) => 
                           MUX_WRdata_OUT_19_port, DATAIN(18) => 
                           MUX_WRdata_OUT_18_port, DATAIN(17) => 
                           MUX_WRdata_OUT_17_port, DATAIN(16) => 
                           MUX_WRdata_OUT_16_port, DATAIN(15) => 
                           MUX_WRdata_OUT_15_port, DATAIN(14) => 
                           MUX_WRdata_OUT_14_port, DATAIN(13) => 
                           MUX_WRdata_OUT_13_port, DATAIN(12) => 
                           MUX_WRdata_OUT_12_port, DATAIN(11) => 
                           MUX_WRdata_OUT_11_port, DATAIN(10) => 
                           MUX_WRdata_OUT_10_port, DATAIN(9) => 
                           MUX_WRdata_OUT_9_port, DATAIN(8) => 
                           MUX_WRdata_OUT_8_port, DATAIN(7) => 
                           MUX_WRdata_OUT_7_port, DATAIN(6) => 
                           MUX_WRdata_OUT_6_port, DATAIN(5) => 
                           MUX_WRdata_OUT_5_port, DATAIN(4) => 
                           MUX_WRdata_OUT_4_port, DATAIN(3) => 
                           MUX_WRdata_OUT_3_port, DATAIN(2) => 
                           MUX_WRdata_OUT_2_port, DATAIN(1) => 
                           MUX_WRdata_OUT_1_port, DATAIN(0) => 
                           MUX_WRdata_OUT_0_port, OUT1(31) => RA_IN_31_port, 
                           OUT1(30) => RA_IN_30_port, OUT1(29) => RA_IN_29_port
                           , OUT1(28) => RA_IN_28_port, OUT1(27) => 
                           RA_IN_27_port, OUT1(26) => RA_IN_26_port, OUT1(25) 
                           => RA_IN_25_port, OUT1(24) => RA_IN_24_port, 
                           OUT1(23) => RA_IN_23_port, OUT1(22) => RA_IN_22_port
                           , OUT1(21) => RA_IN_21_port, OUT1(20) => 
                           RA_IN_20_port, OUT1(19) => RA_IN_19_port, OUT1(18) 
                           => RA_IN_18_port, OUT1(17) => RA_IN_17_port, 
                           OUT1(16) => RA_IN_16_port, OUT1(15) => RA_IN_15_port
                           , OUT1(14) => RA_IN_14_port, OUT1(13) => 
                           RA_IN_13_port, OUT1(12) => RA_IN_12_port, OUT1(11) 
                           => RA_IN_11_port, OUT1(10) => RA_IN_10_port, OUT1(9)
                           => RA_IN_9_port, OUT1(8) => RA_IN_8_port, OUT1(7) =>
                           RA_IN_7_port, OUT1(6) => RA_IN_6_port, OUT1(5) => 
                           RA_IN_5_port, OUT1(4) => RA_IN_4_port, OUT1(3) => 
                           RA_IN_3_port, OUT1(2) => RA_IN_2_port, OUT1(1) => 
                           RA_IN_1_port, OUT1(0) => RA_IN_0_port, OUT2(31) => 
                           RB_IN_31_port, OUT2(30) => RB_IN_30_port, OUT2(29) 
                           => RB_IN_29_port, OUT2(28) => RB_IN_28_port, 
                           OUT2(27) => RB_IN_27_port, OUT2(26) => RB_IN_26_port
                           , OUT2(25) => RB_IN_25_port, OUT2(24) => 
                           RB_IN_24_port, OUT2(23) => RB_IN_23_port, OUT2(22) 
                           => RB_IN_22_port, OUT2(21) => RB_IN_21_port, 
                           OUT2(20) => RB_IN_20_port, OUT2(19) => RB_IN_19_port
                           , OUT2(18) => RB_IN_18_port, OUT2(17) => 
                           RB_IN_17_port, OUT2(16) => RB_IN_16_port, OUT2(15) 
                           => RB_IN_15_port, OUT2(14) => RB_IN_14_port, 
                           OUT2(13) => RB_IN_13_port, OUT2(12) => RB_IN_12_port
                           , OUT2(11) => RB_IN_11_port, OUT2(10) => 
                           RB_IN_10_port, OUT2(9) => RB_IN_9_port, OUT2(8) => 
                           RB_IN_8_port, OUT2(7) => RB_IN_7_port, OUT2(6) => 
                           RB_IN_6_port, OUT2(5) => RB_IN_5_port, OUT2(4) => 
                           RB_IN_4_port, OUT2(3) => RB_IN_3_port, OUT2(2) => 
                           RB_IN_2_port, OUT2(1) => RB_IN_1_port, OUT2(0) => 
                           RB_IN_0_port);
   signExtend_0 : signExtend_NUMBIT_in16_NUMBIT_out32 port map( in_s(15) => 
                           INP2(15), in_s(14) => INP2(14), in_s(13) => INP2(13)
                           , in_s(12) => INP2(12), in_s(11) => INP2(11), 
                           in_s(10) => INP2(10), in_s(9) => INP2(9), in_s(8) =>
                           INP2(8), in_s(7) => INP2(7), in_s(6) => INP2(6), 
                           in_s(5) => INP2(5), in_s(4) => INP2(4), in_s(3) => 
                           INP2(3), in_s(2) => INP2(2), in_s(1) => INP2(1), 
                           in_s(0) => INP2(0), sign_unsign => SIGN_UNSIGN, 
                           out_s(31) => SIGNEXT_IMP2_31_port, out_s(30) => 
                           SIGNEXT_IMP2_30_port, out_s(29) => 
                           SIGNEXT_IMP2_29_port, out_s(28) => 
                           SIGNEXT_IMP2_28_port, out_s(27) => 
                           SIGNEXT_IMP2_27_port, out_s(26) => 
                           SIGNEXT_IMP2_26_port, out_s(25) => 
                           SIGNEXT_IMP2_25_port, out_s(24) => 
                           SIGNEXT_IMP2_24_port, out_s(23) => 
                           SIGNEXT_IMP2_23_port, out_s(22) => 
                           SIGNEXT_IMP2_22_port, out_s(21) => 
                           SIGNEXT_IMP2_21_port, out_s(20) => 
                           SIGNEXT_IMP2_20_port, out_s(19) => 
                           SIGNEXT_IMP2_19_port, out_s(18) => 
                           SIGNEXT_IMP2_18_port, out_s(17) => 
                           SIGNEXT_IMP2_17_port, out_s(16) => 
                           SIGNEXT_IMP2_16_port, out_s(15) => 
                           SIGNEXT_IMP2_15_port, out_s(14) => 
                           SIGNEXT_IMP2_14_port, out_s(13) => 
                           SIGNEXT_IMP2_13_port, out_s(12) => 
                           SIGNEXT_IMP2_12_port, out_s(11) => 
                           SIGNEXT_IMP2_11_port, out_s(10) => 
                           SIGNEXT_IMP2_10_port, out_s(9) => 
                           SIGNEXT_IMP2_9_port, out_s(8) => SIGNEXT_IMP2_8_port
                           , out_s(7) => SIGNEXT_IMP2_7_port, out_s(6) => 
                           SIGNEXT_IMP2_6_port, out_s(5) => SIGNEXT_IMP2_5_port
                           , out_s(4) => SIGNEXT_IMP2_4_port, out_s(3) => 
                           SIGNEXT_IMP2_3_port, out_s(2) => SIGNEXT_IMP2_2_port
                           , out_s(1) => SIGNEXT_IMP2_1_port, out_s(0) => 
                           SIGNEXT_IMP2_0_port);
   signExtend_1 : signExtend_NUMBIT_in26_NUMBIT_out32 port map( in_s(25) => 
                           IMM26(25), in_s(24) => IMM26(24), in_s(23) => 
                           IMM26(23), in_s(22) => IMM26(22), in_s(21) => 
                           IMM26(21), in_s(20) => IMM26(20), in_s(19) => 
                           IMM26(19), in_s(18) => IMM26(18), in_s(17) => 
                           IMM26(17), in_s(16) => IMM26(16), in_s(15) => 
                           IMM26(15), in_s(14) => IMM26(14), in_s(13) => 
                           IMM26(13), in_s(12) => IMM26(12), in_s(11) => 
                           IMM26(11), in_s(10) => IMM26(10), in_s(9) => 
                           IMM26(9), in_s(8) => IMM26(8), in_s(7) => IMM26(7), 
                           in_s(6) => IMM26(6), in_s(5) => IMM26(5), in_s(4) =>
                           IMM26(4), in_s(3) => IMM26(3), in_s(2) => IMM26(2), 
                           in_s(1) => IMM26(1), in_s(0) => IMM26(0), 
                           sign_unsign => X_Logic1_port, out_s(31) => 
                           SIGNEXT_IMM26_31_port, out_s(30) => 
                           SIGNEXT_IMM26_30_port, out_s(29) => 
                           SIGNEXT_IMM26_29_port, out_s(28) => 
                           SIGNEXT_IMM26_28_port, out_s(27) => 
                           SIGNEXT_IMM26_27_port, out_s(26) => 
                           SIGNEXT_IMM26_26_port, out_s(25) => 
                           SIGNEXT_IMM26_25_port, out_s(24) => 
                           SIGNEXT_IMM26_24_port, out_s(23) => 
                           SIGNEXT_IMM26_23_port, out_s(22) => 
                           SIGNEXT_IMM26_22_port, out_s(21) => 
                           SIGNEXT_IMM26_21_port, out_s(20) => 
                           SIGNEXT_IMM26_20_port, out_s(19) => 
                           SIGNEXT_IMM26_19_port, out_s(18) => 
                           SIGNEXT_IMM26_18_port, out_s(17) => 
                           SIGNEXT_IMM26_17_port, out_s(16) => 
                           SIGNEXT_IMM26_16_port, out_s(15) => 
                           SIGNEXT_IMM26_15_port, out_s(14) => 
                           SIGNEXT_IMM26_14_port, out_s(13) => 
                           SIGNEXT_IMM26_13_port, out_s(12) => 
                           SIGNEXT_IMM26_12_port, out_s(11) => 
                           SIGNEXT_IMM26_11_port, out_s(10) => 
                           SIGNEXT_IMM26_10_port, out_s(9) => 
                           SIGNEXT_IMM26_9_port, out_s(8) => 
                           SIGNEXT_IMM26_8_port, out_s(7) => 
                           SIGNEXT_IMM26_7_port, out_s(6) => 
                           SIGNEXT_IMM26_6_port, out_s(5) => 
                           SIGNEXT_IMM26_5_port, out_s(4) => 
                           SIGNEXT_IMM26_4_port, out_s(3) => 
                           SIGNEXT_IMM26_3_port, out_s(2) => 
                           SIGNEXT_IMM26_2_port, out_s(1) => 
                           SIGNEXT_IMM26_1_port, out_s(0) => 
                           SIGNEXT_IMM26_0_port);
   mux_IMM : MUX21_GENERIC_N32_0 port map( A(31) => SIGNEXT_IMP2_31_port, A(30)
                           => SIGNEXT_IMP2_30_port, A(29) => 
                           SIGNEXT_IMP2_29_port, A(28) => SIGNEXT_IMP2_28_port,
                           A(27) => SIGNEXT_IMP2_27_port, A(26) => 
                           SIGNEXT_IMP2_26_port, A(25) => SIGNEXT_IMP2_25_port,
                           A(24) => SIGNEXT_IMP2_24_port, A(23) => 
                           SIGNEXT_IMP2_23_port, A(22) => SIGNEXT_IMP2_22_port,
                           A(21) => SIGNEXT_IMP2_21_port, A(20) => 
                           SIGNEXT_IMP2_20_port, A(19) => SIGNEXT_IMP2_19_port,
                           A(18) => SIGNEXT_IMP2_18_port, A(17) => 
                           SIGNEXT_IMP2_17_port, A(16) => SIGNEXT_IMP2_16_port,
                           A(15) => SIGNEXT_IMP2_15_port, A(14) => 
                           SIGNEXT_IMP2_14_port, A(13) => SIGNEXT_IMP2_13_port,
                           A(12) => SIGNEXT_IMP2_12_port, A(11) => 
                           SIGNEXT_IMP2_11_port, A(10) => SIGNEXT_IMP2_10_port,
                           A(9) => SIGNEXT_IMP2_9_port, A(8) => 
                           SIGNEXT_IMP2_8_port, A(7) => SIGNEXT_IMP2_7_port, 
                           A(6) => SIGNEXT_IMP2_6_port, A(5) => 
                           SIGNEXT_IMP2_5_port, A(4) => SIGNEXT_IMP2_4_port, 
                           A(3) => SIGNEXT_IMP2_3_port, A(2) => 
                           SIGNEXT_IMP2_2_port, A(1) => SIGNEXT_IMP2_1_port, 
                           A(0) => SIGNEXT_IMP2_0_port, B(31) => 
                           SIGNEXT_IMM26_31_port, B(30) => 
                           SIGNEXT_IMM26_30_port, B(29) => 
                           SIGNEXT_IMM26_29_port, B(28) => 
                           SIGNEXT_IMM26_28_port, B(27) => 
                           SIGNEXT_IMM26_27_port, B(26) => 
                           SIGNEXT_IMM26_26_port, B(25) => 
                           SIGNEXT_IMM26_25_port, B(24) => 
                           SIGNEXT_IMM26_24_port, B(23) => 
                           SIGNEXT_IMM26_23_port, B(22) => 
                           SIGNEXT_IMM26_22_port, B(21) => 
                           SIGNEXT_IMM26_21_port, B(20) => 
                           SIGNEXT_IMM26_20_port, B(19) => 
                           SIGNEXT_IMM26_19_port, B(18) => 
                           SIGNEXT_IMM26_18_port, B(17) => 
                           SIGNEXT_IMM26_17_port, B(16) => 
                           SIGNEXT_IMM26_16_port, B(15) => 
                           SIGNEXT_IMM26_15_port, B(14) => 
                           SIGNEXT_IMM26_14_port, B(13) => 
                           SIGNEXT_IMM26_13_port, B(12) => 
                           SIGNEXT_IMM26_12_port, B(11) => 
                           SIGNEXT_IMM26_11_port, B(10) => 
                           SIGNEXT_IMM26_10_port, B(9) => SIGNEXT_IMM26_9_port,
                           B(8) => SIGNEXT_IMM26_8_port, B(7) => 
                           SIGNEXT_IMM26_7_port, B(6) => SIGNEXT_IMM26_6_port, 
                           B(5) => SIGNEXT_IMM26_5_port, B(4) => 
                           SIGNEXT_IMM26_4_port, B(3) => SIGNEXT_IMM26_3_port, 
                           B(2) => SIGNEXT_IMM26_2_port, B(1) => 
                           SIGNEXT_IMM26_1_port, B(0) => SIGNEXT_IMM26_0_port, 
                           SEL => MUX_IMM_SEL, Y(31) => MUX_IMM_OUT_31_port, 
                           Y(30) => MUX_IMM_OUT_30_port, Y(29) => 
                           MUX_IMM_OUT_29_port, Y(28) => MUX_IMM_OUT_28_port, 
                           Y(27) => MUX_IMM_OUT_27_port, Y(26) => 
                           MUX_IMM_OUT_26_port, Y(25) => MUX_IMM_OUT_25_port, 
                           Y(24) => MUX_IMM_OUT_24_port, Y(23) => 
                           MUX_IMM_OUT_23_port, Y(22) => MUX_IMM_OUT_22_port, 
                           Y(21) => MUX_IMM_OUT_21_port, Y(20) => 
                           MUX_IMM_OUT_20_port, Y(19) => MUX_IMM_OUT_19_port, 
                           Y(18) => MUX_IMM_OUT_18_port, Y(17) => 
                           MUX_IMM_OUT_17_port, Y(16) => MUX_IMM_OUT_16_port, 
                           Y(15) => MUX_IMM_OUT_15_port, Y(14) => 
                           MUX_IMM_OUT_14_port, Y(13) => MUX_IMM_OUT_13_port, 
                           Y(12) => MUX_IMM_OUT_12_port, Y(11) => 
                           MUX_IMM_OUT_11_port, Y(10) => MUX_IMM_OUT_10_port, 
                           Y(9) => MUX_IMM_OUT_9_port, Y(8) => 
                           MUX_IMM_OUT_8_port, Y(7) => MUX_IMM_OUT_7_port, Y(6)
                           => MUX_IMM_OUT_6_port, Y(5) => MUX_IMM_OUT_5_port, 
                           Y(4) => MUX_IMM_OUT_4_port, Y(3) => 
                           MUX_IMM_OUT_3_port, Y(2) => MUX_IMM_OUT_2_port, Y(1)
                           => MUX_IMM_OUT_1_port, Y(0) => MUX_IMM_OUT_0_port);
   reg_in1 : reg_NUMBIT32_0 port map( clk => CLK, en => RegIMM_LATCH_EN, rst =>
                           RST, d(31) => INP1(31), d(30) => INP1(30), d(29) => 
                           INP1(29), d(28) => INP1(28), d(27) => INP1(27), 
                           d(26) => INP1(26), d(25) => INP1(25), d(24) => 
                           INP1(24), d(23) => INP1(23), d(22) => INP1(22), 
                           d(21) => INP1(21), d(20) => INP1(20), d(19) => 
                           INP1(19), d(18) => INP1(18), d(17) => INP1(17), 
                           d(16) => INP1(16), d(15) => INP1(15), d(14) => 
                           INP1(14), d(13) => INP1(13), d(12) => INP1(12), 
                           d(11) => INP1(11), d(10) => INP1(10), d(9) => 
                           INP1(9), d(8) => INP1(8), d(7) => INP1(7), d(6) => 
                           INP1(6), d(5) => INP1(5), d(4) => INP1(4), d(3) => 
                           INP1(3), d(2) => INP1(2), d(1) => INP1(1), d(0) => 
                           INP1(0), q(31) => RIMM1_OUT_31_port, q(30) => 
                           RIMM1_OUT_30_port, q(29) => RIMM1_OUT_29_port, q(28)
                           => RIMM1_OUT_28_port, q(27) => RIMM1_OUT_27_port, 
                           q(26) => RIMM1_OUT_26_port, q(25) => 
                           RIMM1_OUT_25_port, q(24) => RIMM1_OUT_24_port, q(23)
                           => RIMM1_OUT_23_port, q(22) => RIMM1_OUT_22_port, 
                           q(21) => RIMM1_OUT_21_port, q(20) => 
                           RIMM1_OUT_20_port, q(19) => RIMM1_OUT_19_port, q(18)
                           => RIMM1_OUT_18_port, q(17) => RIMM1_OUT_17_port, 
                           q(16) => RIMM1_OUT_16_port, q(15) => 
                           RIMM1_OUT_15_port, q(14) => RIMM1_OUT_14_port, q(13)
                           => RIMM1_OUT_13_port, q(12) => RIMM1_OUT_12_port, 
                           q(11) => RIMM1_OUT_11_port, q(10) => 
                           RIMM1_OUT_10_port, q(9) => RIMM1_OUT_9_port, q(8) =>
                           RIMM1_OUT_8_port, q(7) => RIMM1_OUT_7_port, q(6) => 
                           RIMM1_OUT_6_port, q(5) => RIMM1_OUT_5_port, q(4) => 
                           RIMM1_OUT_4_port, q(3) => RIMM1_OUT_3_port, q(2) => 
                           RIMM1_OUT_2_port, q(1) => RIMM1_OUT_1_port, q(0) => 
                           RIMM1_OUT_0_port);
   reg_A : reg_NUMBIT32_9 port map( clk => CLK, en => RegA_LATCH_EN, rst => RST
                           , d(31) => RA_IN_31_port, d(30) => RA_IN_30_port, 
                           d(29) => RA_IN_29_port, d(28) => RA_IN_28_port, 
                           d(27) => RA_IN_27_port, d(26) => RA_IN_26_port, 
                           d(25) => RA_IN_25_port, d(24) => RA_IN_24_port, 
                           d(23) => RA_IN_23_port, d(22) => RA_IN_22_port, 
                           d(21) => RA_IN_21_port, d(20) => RA_IN_20_port, 
                           d(19) => RA_IN_19_port, d(18) => RA_IN_18_port, 
                           d(17) => RA_IN_17_port, d(16) => RA_IN_16_port, 
                           d(15) => RA_IN_15_port, d(14) => RA_IN_14_port, 
                           d(13) => RA_IN_13_port, d(12) => RA_IN_12_port, 
                           d(11) => RA_IN_11_port, d(10) => RA_IN_10_port, d(9)
                           => RA_IN_9_port, d(8) => RA_IN_8_port, d(7) => 
                           RA_IN_7_port, d(6) => RA_IN_6_port, d(5) => 
                           RA_IN_5_port, d(4) => RA_IN_4_port, d(3) => 
                           RA_IN_3_port, d(2) => RA_IN_2_port, d(1) => 
                           RA_IN_1_port, d(0) => RA_IN_0_port, q(31) => 
                           RA_OUT_31_port, q(30) => RA_OUT_30_port, q(29) => 
                           RA_OUT_29_port, q(28) => RA_OUT_28_port, q(27) => 
                           RA_OUT_27_port, q(26) => RA_OUT_26_port, q(25) => 
                           RA_OUT_25_port, q(24) => RA_OUT_24_port, q(23) => 
                           RA_OUT_23_port, q(22) => RA_OUT_22_port, q(21) => 
                           RA_OUT_21_port, q(20) => RA_OUT_20_port, q(19) => 
                           RA_OUT_19_port, q(18) => RA_OUT_18_port, q(17) => 
                           RA_OUT_17_port, q(16) => RA_OUT_16_port, q(15) => 
                           RA_OUT_15_port, q(14) => RA_OUT_14_port, q(13) => 
                           RA_OUT_13_port, q(12) => RA_OUT_12_port, q(11) => 
                           RA_OUT_11_port, q(10) => RA_OUT_10_port, q(9) => 
                           RA_OUT_9_port, q(8) => RA_OUT_8_port, q(7) => 
                           RA_OUT_7_port, q(6) => RA_OUT_6_port, q(5) => 
                           RA_OUT_5_port, q(4) => RA_OUT_4_port, q(3) => 
                           RA_OUT_3_port, q(2) => RA_OUT_2_port, q(1) => 
                           RA_OUT_1_port, q(0) => RA_OUT_0_port);
   reg_B : reg_NUMBIT32_8 port map( clk => CLK, en => RegB_LATCH_EN, rst => RST
                           , d(31) => RB_IN_31_port, d(30) => RB_IN_30_port, 
                           d(29) => RB_IN_29_port, d(28) => RB_IN_28_port, 
                           d(27) => RB_IN_27_port, d(26) => RB_IN_26_port, 
                           d(25) => RB_IN_25_port, d(24) => RB_IN_24_port, 
                           d(23) => RB_IN_23_port, d(22) => RB_IN_22_port, 
                           d(21) => RB_IN_21_port, d(20) => RB_IN_20_port, 
                           d(19) => RB_IN_19_port, d(18) => RB_IN_18_port, 
                           d(17) => RB_IN_17_port, d(16) => RB_IN_16_port, 
                           d(15) => RB_IN_15_port, d(14) => RB_IN_14_port, 
                           d(13) => RB_IN_13_port, d(12) => RB_IN_12_port, 
                           d(11) => RB_IN_11_port, d(10) => RB_IN_10_port, d(9)
                           => RB_IN_9_port, d(8) => RB_IN_8_port, d(7) => 
                           RB_IN_7_port, d(6) => RB_IN_6_port, d(5) => 
                           RB_IN_5_port, d(4) => RB_IN_4_port, d(3) => 
                           RB_IN_3_port, d(2) => RB_IN_2_port, d(1) => 
                           RB_IN_1_port, d(0) => RB_IN_0_port, q(31) => 
                           RB_OUT_31_port, q(30) => RB_OUT_30_port, q(29) => 
                           RB_OUT_29_port, q(28) => RB_OUT_28_port, q(27) => 
                           RB_OUT_27_port, q(26) => RB_OUT_26_port, q(25) => 
                           RB_OUT_25_port, q(24) => RB_OUT_24_port, q(23) => 
                           RB_OUT_23_port, q(22) => RB_OUT_22_port, q(21) => 
                           RB_OUT_21_port, q(20) => RB_OUT_20_port, q(19) => 
                           RB_OUT_19_port, q(18) => RB_OUT_18_port, q(17) => 
                           RB_OUT_17_port, q(16) => RB_OUT_16_port, q(15) => 
                           RB_OUT_15_port, q(14) => RB_OUT_14_port, q(13) => 
                           RB_OUT_13_port, q(12) => RB_OUT_12_port, q(11) => 
                           RB_OUT_11_port, q(10) => RB_OUT_10_port, q(9) => 
                           RB_OUT_9_port, q(8) => RB_OUT_8_port, q(7) => 
                           RB_OUT_7_port, q(6) => RB_OUT_6_port, q(5) => 
                           RB_OUT_5_port, q(4) => RB_OUT_4_port, q(3) => 
                           RB_OUT_3_port, q(2) => RB_OUT_2_port, q(1) => 
                           RB_OUT_1_port, q(0) => RB_OUT_0_port);
   reg_in2 : reg_NUMBIT32_7 port map( clk => CLK, en => RegIMM_LATCH_EN, rst =>
                           RST, d(31) => MUX_IMM_OUT_31_port, d(30) => 
                           MUX_IMM_OUT_30_port, d(29) => MUX_IMM_OUT_29_port, 
                           d(28) => MUX_IMM_OUT_28_port, d(27) => 
                           MUX_IMM_OUT_27_port, d(26) => MUX_IMM_OUT_26_port, 
                           d(25) => MUX_IMM_OUT_25_port, d(24) => 
                           MUX_IMM_OUT_24_port, d(23) => MUX_IMM_OUT_23_port, 
                           d(22) => MUX_IMM_OUT_22_port, d(21) => 
                           MUX_IMM_OUT_21_port, d(20) => MUX_IMM_OUT_20_port, 
                           d(19) => MUX_IMM_OUT_19_port, d(18) => 
                           MUX_IMM_OUT_18_port, d(17) => MUX_IMM_OUT_17_port, 
                           d(16) => n195, d(15) => MUX_IMM_OUT_15_port, d(14) 
                           => MUX_IMM_OUT_14_port, d(13) => MUX_IMM_OUT_13_port
                           , d(12) => MUX_IMM_OUT_12_port, d(11) => 
                           MUX_IMM_OUT_11_port, d(10) => MUX_IMM_OUT_10_port, 
                           d(9) => MUX_IMM_OUT_9_port, d(8) => 
                           MUX_IMM_OUT_8_port, d(7) => MUX_IMM_OUT_7_port, d(6)
                           => MUX_IMM_OUT_6_port, d(5) => MUX_IMM_OUT_5_port, 
                           d(4) => MUX_IMM_OUT_4_port, d(3) => 
                           MUX_IMM_OUT_3_port, d(2) => MUX_IMM_OUT_2_port, d(1)
                           => MUX_IMM_OUT_1_port, d(0) => MUX_IMM_OUT_0_port, 
                           q(31) => RIMM2_OUT_31_port, q(30) => 
                           RIMM2_OUT_30_port, q(29) => RIMM2_OUT_29_port, q(28)
                           => RIMM2_OUT_28_port, q(27) => RIMM2_OUT_27_port, 
                           q(26) => RIMM2_OUT_26_port, q(25) => 
                           RIMM2_OUT_25_port, q(24) => RIMM2_OUT_24_port, q(23)
                           => RIMM2_OUT_23_port, q(22) => RIMM2_OUT_22_port, 
                           q(21) => RIMM2_OUT_21_port, q(20) => 
                           RIMM2_OUT_20_port, q(19) => RIMM2_OUT_19_port, q(18)
                           => RIMM2_OUT_18_port, q(17) => RIMM2_OUT_17_port, 
                           q(16) => RIMM2_OUT_16_port, q(15) => 
                           RIMM2_OUT_15_port, q(14) => RIMM2_OUT_14_port, q(13)
                           => RIMM2_OUT_13_port, q(12) => RIMM2_OUT_12_port, 
                           q(11) => RIMM2_OUT_11_port, q(10) => 
                           RIMM2_OUT_10_port, q(9) => RIMM2_OUT_9_port, q(8) =>
                           RIMM2_OUT_8_port, q(7) => RIMM2_OUT_7_port, q(6) => 
                           RIMM2_OUT_6_port, q(5) => RIMM2_OUT_5_port, q(4) => 
                           RIMM2_OUT_4_port, q(3) => RIMM2_OUT_3_port, q(2) => 
                           RIMM2_OUT_2_port, q(1) => RIMM2_OUT_1_port, q(0) => 
                           RIMM2_OUT_0_port);
   reg_RD1 : reg_NUMBIT5_0 port map( clk => CLK, en => RegRD1_LATCH_EN, rst => 
                           RST, d(4) => RD(4), d(3) => RD(3), d(2) => RD(2), 
                           d(1) => RD(1), d(0) => RD(0), q(4) => RD1_OUT_4_port
                           , q(3) => RD1_OUT_3_port, q(2) => RD1_OUT_2_port, 
                           q(1) => RD1_OUT_1_port, q(0) => RD1_OUT_0_port);
   BranchMgmt_0 : BranchMgmt_NUMBIT32 port map( Rin(31) => 
                           MUX_FORWARDING_BRANCH_OUT_31_port, Rin(30) => 
                           MUX_FORWARDING_BRANCH_OUT_30_port, Rin(29) => 
                           MUX_FORWARDING_BRANCH_OUT_29_port, Rin(28) => 
                           MUX_FORWARDING_BRANCH_OUT_28_port, Rin(27) => 
                           MUX_FORWARDING_BRANCH_OUT_27_port, Rin(26) => 
                           MUX_FORWARDING_BRANCH_OUT_26_port, Rin(25) => 
                           MUX_FORWARDING_BRANCH_OUT_25_port, Rin(24) => 
                           MUX_FORWARDING_BRANCH_OUT_24_port, Rin(23) => 
                           MUX_FORWARDING_BRANCH_OUT_23_port, Rin(22) => 
                           MUX_FORWARDING_BRANCH_OUT_22_port, Rin(21) => 
                           MUX_FORWARDING_BRANCH_OUT_21_port, Rin(20) => 
                           MUX_FORWARDING_BRANCH_OUT_20_port, Rin(19) => 
                           MUX_FORWARDING_BRANCH_OUT_19_port, Rin(18) => 
                           MUX_FORWARDING_BRANCH_OUT_18_port, Rin(17) => 
                           MUX_FORWARDING_BRANCH_OUT_17_port, Rin(16) => 
                           MUX_FORWARDING_BRANCH_OUT_16_port, Rin(15) => 
                           MUX_FORWARDING_BRANCH_OUT_15_port, Rin(14) => 
                           MUX_FORWARDING_BRANCH_OUT_14_port, Rin(13) => 
                           MUX_FORWARDING_BRANCH_OUT_13_port, Rin(12) => 
                           MUX_FORWARDING_BRANCH_OUT_12_port, Rin(11) => 
                           MUX_FORWARDING_BRANCH_OUT_11_port, Rin(10) => 
                           MUX_FORWARDING_BRANCH_OUT_10_port, Rin(9) => 
                           MUX_FORWARDING_BRANCH_OUT_9_port, Rin(8) => 
                           MUX_FORWARDING_BRANCH_OUT_8_port, Rin(7) => 
                           MUX_FORWARDING_BRANCH_OUT_7_port, Rin(6) => 
                           MUX_FORWARDING_BRANCH_OUT_6_port, Rin(5) => 
                           MUX_FORWARDING_BRANCH_OUT_5_port, Rin(4) => 
                           MUX_FORWARDING_BRANCH_OUT_4_port, Rin(3) => 
                           MUX_FORWARDING_BRANCH_OUT_3_port, Rin(2) => 
                           MUX_FORWARDING_BRANCH_OUT_2_port, Rin(1) => 
                           MUX_FORWARDING_BRANCH_OUT_1_port, Rin(0) => 
                           MUX_FORWARDING_BRANCH_OUT_0_port, Cond => EQ_COND, 
                           Jump => JUMP, Branch => BRANCH_T_NT);
   mux_BRANCH : MUX21 port map( A => BRANCH_T_NT, B => X_Logic0_port, SEL => 
                           JUMP_EN, Y => BRANCH_CTRL_SIG);
   mux_A : MUX21_GENERIC_N32_5 port map( A(31) => INP1(31), A(30) => INP1(30), 
                           A(29) => INP1(29), A(28) => INP1(28), A(27) => 
                           INP1(27), A(26) => INP1(26), A(25) => INP1(25), 
                           A(24) => INP1(24), A(23) => INP1(23), A(22) => 
                           INP1(22), A(21) => INP1(21), A(20) => INP1(20), 
                           A(19) => INP1(19), A(18) => INP1(18), A(17) => 
                           INP1(17), A(16) => INP1(16), A(15) => INP1(15), 
                           A(14) => INP1(14), A(13) => INP1(13), A(12) => 
                           INP1(12), A(11) => INP1(11), A(10) => INP1(10), A(9)
                           => INP1(9), A(8) => INP1(8), A(7) => INP1(7), A(6) 
                           => INP1(6), A(5) => INP1(5), A(4) => INP1(4), A(3) 
                           => INP1(3), A(2) => INP1(2), A(1) => INP1(1), A(0) 
                           => INP1(0), B(31) => 
                           MUX_FORWARDING_BRANCH_OUT_31_port, B(30) => 
                           MUX_FORWARDING_BRANCH_OUT_30_port, B(29) => 
                           MUX_FORWARDING_BRANCH_OUT_29_port, B(28) => 
                           MUX_FORWARDING_BRANCH_OUT_28_port, B(27) => 
                           MUX_FORWARDING_BRANCH_OUT_27_port, B(26) => 
                           MUX_FORWARDING_BRANCH_OUT_26_port, B(25) => 
                           MUX_FORWARDING_BRANCH_OUT_25_port, B(24) => 
                           MUX_FORWARDING_BRANCH_OUT_24_port, B(23) => 
                           MUX_FORWARDING_BRANCH_OUT_23_port, B(22) => 
                           MUX_FORWARDING_BRANCH_OUT_22_port, B(21) => 
                           MUX_FORWARDING_BRANCH_OUT_21_port, B(20) => 
                           MUX_FORWARDING_BRANCH_OUT_20_port, B(19) => 
                           MUX_FORWARDING_BRANCH_OUT_19_port, B(18) => 
                           MUX_FORWARDING_BRANCH_OUT_18_port, B(17) => 
                           MUX_FORWARDING_BRANCH_OUT_17_port, B(16) => 
                           MUX_FORWARDING_BRANCH_OUT_16_port, B(15) => 
                           MUX_FORWARDING_BRANCH_OUT_15_port, B(14) => 
                           MUX_FORWARDING_BRANCH_OUT_14_port, B(13) => 
                           MUX_FORWARDING_BRANCH_OUT_13_port, B(12) => 
                           MUX_FORWARDING_BRANCH_OUT_12_port, B(11) => 
                           MUX_FORWARDING_BRANCH_OUT_11_port, B(10) => n204, 
                           B(9) => MUX_FORWARDING_BRANCH_OUT_9_port, B(8) => 
                           MUX_FORWARDING_BRANCH_OUT_8_port, B(7) => 
                           MUX_FORWARDING_BRANCH_OUT_7_port, B(6) => 
                           MUX_FORWARDING_BRANCH_OUT_6_port, B(5) => 
                           MUX_FORWARDING_BRANCH_OUT_5_port, B(4) => 
                           MUX_FORWARDING_BRANCH_OUT_4_port, B(3) => n205, B(2)
                           => MUX_FORWARDING_BRANCH_OUT_2_port, B(1) => 
                           MUX_FORWARDING_BRANCH_OUT_1_port, B(0) => 
                           MUX_FORWARDING_BRANCH_OUT_0_port, SEL => MUXA_SEL, 
                           Y(31) => MUXA_OUT_31_port, Y(30) => MUXA_OUT_30_port
                           , Y(29) => MUXA_OUT_29_port, Y(28) => 
                           MUXA_OUT_28_port, Y(27) => MUXA_OUT_27_port, Y(26) 
                           => MUXA_OUT_26_port, Y(25) => MUXA_OUT_25_port, 
                           Y(24) => MUXA_OUT_24_port, Y(23) => MUXA_OUT_23_port
                           , Y(22) => MUXA_OUT_22_port, Y(21) => 
                           MUXA_OUT_21_port, Y(20) => MUXA_OUT_20_port, Y(19) 
                           => MUXA_OUT_19_port, Y(18) => MUXA_OUT_18_port, 
                           Y(17) => MUXA_OUT_17_port, Y(16) => MUXA_OUT_16_port
                           , Y(15) => MUXA_OUT_15_port, Y(14) => 
                           MUXA_OUT_14_port, Y(13) => MUXA_OUT_13_port, Y(12) 
                           => MUXA_OUT_12_port, Y(11) => MUXA_OUT_11_port, 
                           Y(10) => MUXA_OUT_10_port, Y(9) => MUXA_OUT_9_port, 
                           Y(8) => MUXA_OUT_8_port, Y(7) => MUXA_OUT_7_port, 
                           Y(6) => MUXA_OUT_6_port, Y(5) => MUXA_OUT_5_port, 
                           Y(4) => MUXA_OUT_4_port, Y(3) => MUXA_OUT_3_port, 
                           Y(2) => MUXA_OUT_2_port, Y(1) => MUXA_OUT_1_port, 
                           Y(0) => MUXA_OUT_0_port);
   mux_B : MUX21_GENERIC_N32_4 port map( A(31) => ALU_inputB_31_port, A(30) => 
                           ALU_inputB_30_port, A(29) => ALU_inputB_29_port, 
                           A(28) => ALU_inputB_28_port, A(27) => 
                           ALU_inputB_27_port, A(26) => ALU_inputB_26_port, 
                           A(25) => ALU_inputB_25_port, A(24) => 
                           ALU_inputB_24_port, A(23) => ALU_inputB_23_port, 
                           A(22) => ALU_inputB_22_port, A(21) => 
                           ALU_inputB_21_port, A(20) => ALU_inputB_20_port, 
                           A(19) => ALU_inputB_19_port, A(18) => 
                           ALU_inputB_18_port, A(17) => ALU_inputB_17_port, 
                           A(16) => ALU_inputB_16_port, A(15) => 
                           ALU_inputB_15_port, A(14) => ALU_inputB_14_port, 
                           A(13) => ALU_inputB_13_port, A(12) => 
                           ALU_inputB_12_port, A(11) => ALU_inputB_11_port, 
                           A(10) => ALU_inputB_10_port, A(9) => 
                           ALU_inputB_9_port, A(8) => ALU_inputB_8_port, A(7) 
                           => ALU_inputB_7_port, A(6) => ALU_inputB_6_port, 
                           A(5) => ALU_inputB_5_port, A(4) => ALU_inputB_4_port
                           , A(3) => ALU_inputB_3_port, A(2) => 
                           ALU_inputB_2_port, A(1) => ALU_inputB_1_port, A(0) 
                           => ALU_inputB_0_port, B(31) => RIMM2_OUT_31_port, 
                           B(30) => RIMM2_OUT_30_port, B(29) => 
                           RIMM2_OUT_29_port, B(28) => RIMM2_OUT_28_port, B(27)
                           => RIMM2_OUT_27_port, B(26) => RIMM2_OUT_26_port, 
                           B(25) => RIMM2_OUT_25_port, B(24) => 
                           RIMM2_OUT_24_port, B(23) => RIMM2_OUT_23_port, B(22)
                           => RIMM2_OUT_22_port, B(21) => RIMM2_OUT_21_port, 
                           B(20) => RIMM2_OUT_20_port, B(19) => 
                           RIMM2_OUT_19_port, B(18) => RIMM2_OUT_18_port, B(17)
                           => RIMM2_OUT_17_port, B(16) => RIMM2_OUT_16_port, 
                           B(15) => RIMM2_OUT_15_port, B(14) => 
                           RIMM2_OUT_14_port, B(13) => RIMM2_OUT_13_port, B(12)
                           => RIMM2_OUT_12_port, B(11) => RIMM2_OUT_11_port, 
                           B(10) => RIMM2_OUT_10_port, B(9) => RIMM2_OUT_9_port
                           , B(8) => RIMM2_OUT_8_port, B(7) => RIMM2_OUT_7_port
                           , B(6) => RIMM2_OUT_6_port, B(5) => RIMM2_OUT_5_port
                           , B(4) => RIMM2_OUT_4_port, B(3) => RIMM2_OUT_3_port
                           , B(2) => RIMM2_OUT_2_port, B(1) => RIMM2_OUT_1_port
                           , B(0) => RIMM2_OUT_0_port, SEL => MUXB_SEL, Y(31) 
                           => MUXB_OUT_31_port, Y(30) => MUXB_OUT_30_port, 
                           Y(29) => MUXB_OUT_29_port, Y(28) => MUXB_OUT_28_port
                           , Y(27) => MUXB_OUT_27_port, Y(26) => 
                           MUXB_OUT_26_port, Y(25) => MUXB_OUT_25_port, Y(24) 
                           => MUXB_OUT_24_port, Y(23) => MUXB_OUT_23_port, 
                           Y(22) => MUXB_OUT_22_port, Y(21) => MUXB_OUT_21_port
                           , Y(20) => MUXB_OUT_20_port, Y(19) => 
                           MUXB_OUT_19_port, Y(18) => MUXB_OUT_18_port, Y(17) 
                           => MUXB_OUT_17_port, Y(16) => MUXB_OUT_16_port, 
                           Y(15) => MUXB_OUT_15_port, Y(14) => MUXB_OUT_14_port
                           , Y(13) => MUXB_OUT_13_port, Y(12) => 
                           MUXB_OUT_12_port, Y(11) => MUXB_OUT_11_port, Y(10) 
                           => MUXB_OUT_10_port, Y(9) => MUXB_OUT_9_port, Y(8) 
                           => MUXB_OUT_8_port, Y(7) => MUXB_OUT_7_port, Y(6) =>
                           MUXB_OUT_6_port, Y(5) => MUXB_OUT_5_port, Y(4) => 
                           MUXB_OUT_4_port, Y(3) => MUXB_OUT_3_port, Y(2) => 
                           MUXB_OUT_2_port, Y(1) => MUXB_OUT_1_port, Y(0) => 
                           MUXB_OUT_0_port);
   reg_ALUOUT : reg_NUMBIT32_6 port map( clk => CLK, en => RALUOUT_LATCH_EN, 
                           rst => RST, d(31) => ALU_OUT_31_port, d(30) => 
                           ALU_OUT_30_port, d(29) => ALU_OUT_29_port, d(28) => 
                           ALU_OUT_28_port, d(27) => ALU_OUT_27_port, d(26) => 
                           ALU_OUT_26_port, d(25) => ALU_OUT_25_port, d(24) => 
                           ALU_OUT_24_port, d(23) => ALU_OUT_23_port, d(22) => 
                           ALU_OUT_22_port, d(21) => ALU_OUT_21_port, d(20) => 
                           ALU_OUT_20_port, d(19) => ALU_OUT_19_port, d(18) => 
                           ALU_OUT_18_port, d(17) => ALU_OUT_17_port, d(16) => 
                           ALU_OUT_16_port, d(15) => ALU_OUT_15_port, d(14) => 
                           ALU_OUT_14_port, d(13) => ALU_OUT_13_port, d(12) => 
                           ALU_OUT_12_port, d(11) => ALU_OUT_11_port, d(10) => 
                           ALU_OUT_10_port, d(9) => ALU_OUT_9_port, d(8) => 
                           ALU_OUT_8_port, d(7) => ALU_OUT_7_port, d(6) => 
                           ALU_OUT_6_port, d(5) => ALU_OUT_5_port, d(4) => 
                           ALU_OUT_4_port, d(3) => ALU_OUT_3_port, d(2) => 
                           ALU_OUT_2_port, d(1) => ALU_OUT_1_port, d(0) => 
                           ALU_OUT_0_port, q(31) => ADDR_DRAM_31_port, q(30) =>
                           ADDR_DRAM_30_port, q(29) => ADDR_DRAM_29_port, q(28)
                           => ADDR_DRAM_28_port, q(27) => ADDR_DRAM_27_port, 
                           q(26) => ADDR_DRAM_26_port, q(25) => 
                           ADDR_DRAM_25_port, q(24) => ADDR_DRAM_24_port, q(23)
                           => ADDR_DRAM_23_port, q(22) => ADDR_DRAM_22_port, 
                           q(21) => ADDR_DRAM_21_port, q(20) => 
                           ADDR_DRAM_20_port, q(19) => ADDR_DRAM_19_port, q(18)
                           => ADDR_DRAM_18_port, q(17) => ADDR_DRAM_17_port, 
                           q(16) => ADDR_DRAM_16_port, q(15) => 
                           ADDR_DRAM_15_port, q(14) => ADDR_DRAM_14_port, q(13)
                           => ADDR_DRAM_13_port, q(12) => ADDR_DRAM_12_port, 
                           q(11) => ADDR_DRAM_11_port, q(10) => 
                           ADDR_DRAM_10_port, q(9) => ADDR_DRAM_9_port, q(8) =>
                           ADDR_DRAM_8_port, q(7) => ADDR_DRAM_7_port, q(6) => 
                           ADDR_DRAM_6_port, q(5) => ADDR_DRAM_5_port, q(4) => 
                           ADDR_DRAM_4_port, q(3) => ADDR_DRAM_3_port, q(2) => 
                           ADDR_DRAM_2_port, q(1) => ADDR_DRAM_1_port, q(0) => 
                           ADDR_DRAM_0_port);
   reg_ME : reg_NUMBIT32_5 port map( clk => CLK, en => REGME_LATCH_EN, rst => 
                           RST, d(31) => RB_OUT_31_port, d(30) => 
                           RB_OUT_30_port, d(29) => RB_OUT_29_port, d(28) => 
                           RB_OUT_28_port, d(27) => RB_OUT_27_port, d(26) => 
                           RB_OUT_26_port, d(25) => RB_OUT_25_port, d(24) => 
                           RB_OUT_24_port, d(23) => RB_OUT_23_port, d(22) => 
                           RB_OUT_22_port, d(21) => RB_OUT_21_port, d(20) => 
                           RB_OUT_20_port, d(19) => RB_OUT_19_port, d(18) => 
                           RB_OUT_18_port, d(17) => RB_OUT_17_port, d(16) => 
                           RB_OUT_16_port, d(15) => RB_OUT_15_port, d(14) => 
                           RB_OUT_14_port, d(13) => RB_OUT_13_port, d(12) => 
                           RB_OUT_12_port, d(11) => RB_OUT_11_port, d(10) => 
                           RB_OUT_10_port, d(9) => RB_OUT_9_port, d(8) => 
                           RB_OUT_8_port, d(7) => RB_OUT_7_port, d(6) => 
                           RB_OUT_6_port, d(5) => RB_OUT_5_port, d(4) => 
                           RB_OUT_4_port, d(3) => RB_OUT_3_port, d(2) => 
                           RB_OUT_2_port, d(1) => RB_OUT_1_port, d(0) => 
                           RB_OUT_0_port, q(31) => RME_OUT_31_port, q(30) => 
                           RME_OUT_30_port, q(29) => RME_OUT_29_port, q(28) => 
                           RME_OUT_28_port, q(27) => RME_OUT_27_port, q(26) => 
                           RME_OUT_26_port, q(25) => RME_OUT_25_port, q(24) => 
                           RME_OUT_24_port, q(23) => RME_OUT_23_port, q(22) => 
                           RME_OUT_22_port, q(21) => RME_OUT_21_port, q(20) => 
                           RME_OUT_20_port, q(19) => RME_OUT_19_port, q(18) => 
                           RME_OUT_18_port, q(17) => RME_OUT_17_port, q(16) => 
                           RME_OUT_16_port, q(15) => RME_OUT_15_port, q(14) => 
                           RME_OUT_14_port, q(13) => RME_OUT_13_port, q(12) => 
                           RME_OUT_12_port, q(11) => RME_OUT_11_port, q(10) => 
                           RME_OUT_10_port, q(9) => RME_OUT_9_port, q(8) => 
                           RME_OUT_8_port, q(7) => RME_OUT_7_port, q(6) => 
                           RME_OUT_6_port, q(5) => RME_OUT_5_port, q(4) => 
                           RME_OUT_4_port, q(3) => RME_OUT_3_port, q(2) => 
                           RME_OUT_2_port, q(1) => RME_OUT_1_port, q(0) => 
                           RME_OUT_0_port);
   reg_RD2 : reg_NUMBIT5_2 port map( clk => CLK, en => RegRD2_LATCH_EN, rst => 
                           RST, d(4) => RD1_OUT_4_port, d(3) => RD1_OUT_3_port,
                           d(2) => RD1_OUT_2_port, d(1) => RD1_OUT_1_port, d(0)
                           => RD1_OUT_0_port, q(4) => RD2_OUT_4_port, q(3) => 
                           RD2_OUT_3_port, q(2) => RD2_OUT_2_port, q(1) => 
                           RD2_OUT_1_port, q(0) => RD2_OUT_0_port);
   reg_LMD : reg_NUMBIT32_4 port map( clk => CLK, en => LMD_LATCH_EN, rst => 
                           RST, d(31) => DATAOUT_DRAM(31), d(30) => 
                           DATAOUT_DRAM(30), d(29) => DATAOUT_DRAM(29), d(28) 
                           => DATAOUT_DRAM(28), d(27) => DATAOUT_DRAM(27), 
                           d(26) => DATAOUT_DRAM(26), d(25) => DATAOUT_DRAM(25)
                           , d(24) => DATAOUT_DRAM(24), d(23) => 
                           DATAOUT_DRAM(23), d(22) => DATAOUT_DRAM(22), d(21) 
                           => DATAOUT_DRAM(21), d(20) => DATAOUT_DRAM(20), 
                           d(19) => DATAOUT_DRAM(19), d(18) => DATAOUT_DRAM(18)
                           , d(17) => DATAOUT_DRAM(17), d(16) => 
                           DATAOUT_DRAM(16), d(15) => DATAOUT_DRAM(15), d(14) 
                           => DATAOUT_DRAM(14), d(13) => DATAOUT_DRAM(13), 
                           d(12) => DATAOUT_DRAM(12), d(11) => DATAOUT_DRAM(11)
                           , d(10) => DATAOUT_DRAM(10), d(9) => DATAOUT_DRAM(9)
                           , d(8) => DATAOUT_DRAM(8), d(7) => DATAOUT_DRAM(7), 
                           d(6) => DATAOUT_DRAM(6), d(5) => DATAOUT_DRAM(5), 
                           d(4) => DATAOUT_DRAM(4), d(3) => DATAOUT_DRAM(3), 
                           d(2) => DATAOUT_DRAM(2), d(1) => DATAOUT_DRAM(1), 
                           d(0) => DATAOUT_DRAM(0), q(31) => LMD_OUT_31_port, 
                           q(30) => LMD_OUT_30_port, q(29) => LMD_OUT_29_port, 
                           q(28) => LMD_OUT_28_port, q(27) => LMD_OUT_27_port, 
                           q(26) => LMD_OUT_26_port, q(25) => LMD_OUT_25_port, 
                           q(24) => LMD_OUT_24_port, q(23) => LMD_OUT_23_port, 
                           q(22) => LMD_OUT_22_port, q(21) => LMD_OUT_21_port, 
                           q(20) => LMD_OUT_20_port, q(19) => LMD_OUT_19_port, 
                           q(18) => LMD_OUT_18_port, q(17) => LMD_OUT_17_port, 
                           q(16) => LMD_OUT_16_port, q(15) => LMD_OUT_15_port, 
                           q(14) => LMD_OUT_14_port, q(13) => LMD_OUT_13_port, 
                           q(12) => LMD_OUT_12_port, q(11) => LMD_OUT_11_port, 
                           q(10) => LMD_OUT_10_port, q(9) => LMD_OUT_9_port, 
                           q(8) => LMD_OUT_8_port, q(7) => LMD_OUT_7_port, q(6)
                           => LMD_OUT_6_port, q(5) => LMD_OUT_5_port, q(4) => 
                           LMD_OUT_4_port, q(3) => LMD_OUT_3_port, q(2) => 
                           LMD_OUT_2_port, q(1) => LMD_OUT_1_port, q(0) => 
                           LMD_OUT_0_port);
   reg_ALUOUT2 : reg_NUMBIT32_3 port map( clk => CLK, en => RALUOUT2_LATCH_EN, 
                           rst => RST, d(31) => ADDR_DRAM_31_port, d(30) => 
                           ADDR_DRAM_30_port, d(29) => ADDR_DRAM_29_port, d(28)
                           => ADDR_DRAM_28_port, d(27) => ADDR_DRAM_27_port, 
                           d(26) => ADDR_DRAM_26_port, d(25) => 
                           ADDR_DRAM_25_port, d(24) => ADDR_DRAM_24_port, d(23)
                           => ADDR_DRAM_23_port, d(22) => ADDR_DRAM_22_port, 
                           d(21) => ADDR_DRAM_21_port, d(20) => 
                           ADDR_DRAM_20_port, d(19) => ADDR_DRAM_19_port, d(18)
                           => ADDR_DRAM_18_port, d(17) => ADDR_DRAM_17_port, 
                           d(16) => ADDR_DRAM_16_port, d(15) => 
                           ADDR_DRAM_15_port, d(14) => ADDR_DRAM_14_port, d(13)
                           => ADDR_DRAM_13_port, d(12) => ADDR_DRAM_12_port, 
                           d(11) => ADDR_DRAM_11_port, d(10) => 
                           ADDR_DRAM_10_port, d(9) => ADDR_DRAM_9_port, d(8) =>
                           ADDR_DRAM_8_port, d(7) => ADDR_DRAM_7_port, d(6) => 
                           ADDR_DRAM_6_port, d(5) => ADDR_DRAM_5_port, d(4) => 
                           ADDR_DRAM_4_port, d(3) => ADDR_DRAM_3_port, d(2) => 
                           ADDR_DRAM_2_port, d(1) => ADDR_DRAM_1_port, d(0) => 
                           ADDR_DRAM_0_port, q(31) => RALUOUT2_OUT_31_port, 
                           q(30) => RALUOUT2_OUT_30_port, q(29) => 
                           RALUOUT2_OUT_29_port, q(28) => RALUOUT2_OUT_28_port,
                           q(27) => RALUOUT2_OUT_27_port, q(26) => 
                           RALUOUT2_OUT_26_port, q(25) => RALUOUT2_OUT_25_port,
                           q(24) => RALUOUT2_OUT_24_port, q(23) => 
                           RALUOUT2_OUT_23_port, q(22) => RALUOUT2_OUT_22_port,
                           q(21) => RALUOUT2_OUT_21_port, q(20) => 
                           RALUOUT2_OUT_20_port, q(19) => RALUOUT2_OUT_19_port,
                           q(18) => RALUOUT2_OUT_18_port, q(17) => 
                           RALUOUT2_OUT_17_port, q(16) => RALUOUT2_OUT_16_port,
                           q(15) => RALUOUT2_OUT_15_port, q(14) => 
                           RALUOUT2_OUT_14_port, q(13) => RALUOUT2_OUT_13_port,
                           q(12) => RALUOUT2_OUT_12_port, q(11) => 
                           RALUOUT2_OUT_11_port, q(10) => RALUOUT2_OUT_10_port,
                           q(9) => RALUOUT2_OUT_9_port, q(8) => 
                           RALUOUT2_OUT_8_port, q(7) => RALUOUT2_OUT_7_port, 
                           q(6) => RALUOUT2_OUT_6_port, q(5) => 
                           RALUOUT2_OUT_5_port, q(4) => RALUOUT2_OUT_4_port, 
                           q(3) => RALUOUT2_OUT_3_port, q(2) => 
                           RALUOUT2_OUT_2_port, q(1) => RALUOUT2_OUT_1_port, 
                           q(0) => RALUOUT2_OUT_0_port);
   reg_RD3 : reg_NUMBIT5_1 port map( clk => CLK, en => RegRD3_LATCH_EN, rst => 
                           RST, d(4) => n196, d(3) => n203, d(2) => n197, d(1) 
                           => n198, d(0) => n199, q(4) => RD3_OUT_4_port, q(3) 
                           => RD3_OUT_3_port, q(2) => RD3_OUT_2_port, q(1) => 
                           RD3_OUT_1_port, q(0) => RD3_OUT_0_port);
   PCplus8 : reg_NUMBIT32_2 port map( clk => CLK, en => RPCplus8_LATCH_EN, rst 
                           => RST, d(31) => RIMM1_OUT_31_port, d(30) => 
                           RIMM1_OUT_30_port, d(29) => RIMM1_OUT_29_port, d(28)
                           => RIMM1_OUT_28_port, d(27) => RIMM1_OUT_27_port, 
                           d(26) => RIMM1_OUT_26_port, d(25) => 
                           RIMM1_OUT_25_port, d(24) => RIMM1_OUT_24_port, d(23)
                           => RIMM1_OUT_23_port, d(22) => RIMM1_OUT_22_port, 
                           d(21) => RIMM1_OUT_21_port, d(20) => 
                           RIMM1_OUT_20_port, d(19) => RIMM1_OUT_19_port, d(18)
                           => RIMM1_OUT_18_port, d(17) => RIMM1_OUT_17_port, 
                           d(16) => RIMM1_OUT_16_port, d(15) => 
                           RIMM1_OUT_15_port, d(14) => RIMM1_OUT_14_port, d(13)
                           => RIMM1_OUT_13_port, d(12) => RIMM1_OUT_12_port, 
                           d(11) => RIMM1_OUT_11_port, d(10) => 
                           RIMM1_OUT_10_port, d(9) => RIMM1_OUT_9_port, d(8) =>
                           RIMM1_OUT_8_port, d(7) => RIMM1_OUT_7_port, d(6) => 
                           RIMM1_OUT_6_port, d(5) => RIMM1_OUT_5_port, d(4) => 
                           RIMM1_OUT_4_port, d(3) => RIMM1_OUT_3_port, d(2) => 
                           RIMM1_OUT_2_port, d(1) => RIMM1_OUT_1_port, d(0) => 
                           RIMM1_OUT_0_port, q(31) => RPCplus8_OUT_31_port, 
                           q(30) => RPCplus8_OUT_30_port, q(29) => 
                           RPCplus8_OUT_29_port, q(28) => RPCplus8_OUT_28_port,
                           q(27) => RPCplus8_OUT_27_port, q(26) => 
                           RPCplus8_OUT_26_port, q(25) => RPCplus8_OUT_25_port,
                           q(24) => RPCplus8_OUT_24_port, q(23) => 
                           RPCplus8_OUT_23_port, q(22) => RPCplus8_OUT_22_port,
                           q(21) => RPCplus8_OUT_21_port, q(20) => 
                           RPCplus8_OUT_20_port, q(19) => RPCplus8_OUT_19_port,
                           q(18) => RPCplus8_OUT_18_port, q(17) => 
                           RPCplus8_OUT_17_port, q(16) => RPCplus8_OUT_16_port,
                           q(15) => RPCplus8_OUT_15_port, q(14) => 
                           RPCplus8_OUT_14_port, q(13) => RPCplus8_OUT_13_port,
                           q(12) => RPCplus8_OUT_12_port, q(11) => 
                           RPCplus8_OUT_11_port, q(10) => RPCplus8_OUT_10_port,
                           q(9) => RPCplus8_OUT_9_port, q(8) => 
                           RPCplus8_OUT_8_port, q(7) => RPCplus8_OUT_7_port, 
                           q(6) => RPCplus8_OUT_6_port, q(5) => 
                           RPCplus8_OUT_5_port, q(4) => RPCplus8_OUT_4_port, 
                           q(3) => RPCplus8_OUT_3_port, q(2) => 
                           RPCplus8_OUT_2_port, q(1) => RPCplus8_OUT_1_port, 
                           q(0) => RPCplus8_OUT_0_port);
   MUX_FORWARD_MEM : MUX21_GENERIC_N32_3 port map( A(31) => MUXC_OUT_31_port, 
                           A(30) => MUXC_OUT_30_port, A(29) => MUXC_OUT_29_port
                           , A(28) => MUXC_OUT_28_port, A(27) => 
                           MUXC_OUT_27_port, A(26) => MUXC_OUT_26_port, A(25) 
                           => MUXC_OUT_25_port, A(24) => MUXC_OUT_24_port, 
                           A(23) => MUXC_OUT_23_port, A(22) => MUXC_OUT_22_port
                           , A(21) => MUXC_OUT_21_port, A(20) => 
                           MUXC_OUT_20_port, A(19) => MUXC_OUT_19_port, A(18) 
                           => MUXC_OUT_18_port, A(17) => MUXC_OUT_17_port, 
                           A(16) => MUXC_OUT_16_port, A(15) => MUXC_OUT_15_port
                           , A(14) => MUXC_OUT_14_port, A(13) => 
                           MUXC_OUT_13_port, A(12) => MUXC_OUT_12_port, A(11) 
                           => MUXC_OUT_11_port, A(10) => MUXC_OUT_10_port, A(9)
                           => MUXC_OUT_9_port, A(8) => MUXC_OUT_8_port, A(7) =>
                           MUXC_OUT_7_port, A(6) => MUXC_OUT_6_port, A(5) => 
                           MUXC_OUT_5_port, A(4) => MUXC_OUT_4_port, A(3) => 
                           MUXC_OUT_3_port, A(2) => MUXC_OUT_2_port, A(1) => 
                           MUXC_OUT_1_port, A(0) => MUXC_OUT_0_port, B(31) => 
                           RME_OUT_31_port, B(30) => RME_OUT_30_port, B(29) => 
                           RME_OUT_29_port, B(28) => RME_OUT_28_port, B(27) => 
                           RME_OUT_27_port, B(26) => RME_OUT_26_port, B(25) => 
                           RME_OUT_25_port, B(24) => RME_OUT_24_port, B(23) => 
                           RME_OUT_23_port, B(22) => RME_OUT_22_port, B(21) => 
                           RME_OUT_21_port, B(20) => RME_OUT_20_port, B(19) => 
                           RME_OUT_19_port, B(18) => RME_OUT_18_port, B(17) => 
                           RME_OUT_17_port, B(16) => RME_OUT_16_port, B(15) => 
                           RME_OUT_15_port, B(14) => RME_OUT_14_port, B(13) => 
                           RME_OUT_13_port, B(12) => RME_OUT_12_port, B(11) => 
                           RME_OUT_11_port, B(10) => RME_OUT_10_port, B(9) => 
                           RME_OUT_9_port, B(8) => RME_OUT_8_port, B(7) => 
                           RME_OUT_7_port, B(6) => RME_OUT_6_port, B(5) => 
                           RME_OUT_5_port, B(4) => RME_OUT_4_port, B(3) => 
                           RME_OUT_3_port, B(2) => RME_OUT_2_port, B(1) => 
                           RME_OUT_1_port, B(0) => RME_OUT_0_port, SEL => 
                           ForwardC, Y(31) => DATAIN_DRAM(31), Y(30) => 
                           DATAIN_DRAM(30), Y(29) => DATAIN_DRAM(29), Y(28) => 
                           DATAIN_DRAM(28), Y(27) => DATAIN_DRAM(27), Y(26) => 
                           DATAIN_DRAM(26), Y(25) => DATAIN_DRAM(25), Y(24) => 
                           DATAIN_DRAM(24), Y(23) => DATAIN_DRAM(23), Y(22) => 
                           DATAIN_DRAM(22), Y(21) => DATAIN_DRAM(21), Y(20) => 
                           DATAIN_DRAM(20), Y(19) => DATAIN_DRAM(19), Y(18) => 
                           DATAIN_DRAM(18), Y(17) => DATAIN_DRAM(17), Y(16) => 
                           DATAIN_DRAM(16), Y(15) => DATAIN_DRAM(15), Y(14) => 
                           DATAIN_DRAM(14), Y(13) => DATAIN_DRAM(13), Y(12) => 
                           DATAIN_DRAM(12), Y(11) => DATAIN_DRAM(11), Y(10) => 
                           DATAIN_DRAM(10), Y(9) => DATAIN_DRAM(9), Y(8) => 
                           DATAIN_DRAM(8), Y(7) => DATAIN_DRAM(7), Y(6) => 
                           DATAIN_DRAM(6), Y(5) => DATAIN_DRAM(5), Y(4) => 
                           DATAIN_DRAM(4), Y(3) => DATAIN_DRAM(3), Y(2) => 
                           DATAIN_DRAM(2), Y(1) => DATAIN_DRAM(1), Y(0) => 
                           DATAIN_DRAM(0));
   mux_C : MUX21_GENERIC_N32_2 port map( A(31) => LMD_OUT_31_port, A(30) => 
                           LMD_OUT_30_port, A(29) => LMD_OUT_29_port, A(28) => 
                           LMD_OUT_28_port, A(27) => LMD_OUT_27_port, A(26) => 
                           LMD_OUT_26_port, A(25) => LMD_OUT_25_port, A(24) => 
                           LMD_OUT_24_port, A(23) => LMD_OUT_23_port, A(22) => 
                           LMD_OUT_22_port, A(21) => LMD_OUT_21_port, A(20) => 
                           LMD_OUT_20_port, A(19) => LMD_OUT_19_port, A(18) => 
                           LMD_OUT_18_port, A(17) => LMD_OUT_17_port, A(16) => 
                           LMD_OUT_16_port, A(15) => LMD_OUT_15_port, A(14) => 
                           LMD_OUT_14_port, A(13) => LMD_OUT_13_port, A(12) => 
                           LMD_OUT_12_port, A(11) => LMD_OUT_11_port, A(10) => 
                           LMD_OUT_10_port, A(9) => LMD_OUT_9_port, A(8) => 
                           LMD_OUT_8_port, A(7) => LMD_OUT_7_port, A(6) => 
                           LMD_OUT_6_port, A(5) => LMD_OUT_5_port, A(4) => 
                           LMD_OUT_4_port, A(3) => LMD_OUT_3_port, A(2) => 
                           LMD_OUT_2_port, A(1) => LMD_OUT_1_port, A(0) => 
                           LMD_OUT_0_port, B(31) => RALUOUT2_OUT_31_port, B(30)
                           => RALUOUT2_OUT_30_port, B(29) => 
                           RALUOUT2_OUT_29_port, B(28) => RALUOUT2_OUT_28_port,
                           B(27) => RALUOUT2_OUT_27_port, B(26) => 
                           RALUOUT2_OUT_26_port, B(25) => RALUOUT2_OUT_25_port,
                           B(24) => RALUOUT2_OUT_24_port, B(23) => 
                           RALUOUT2_OUT_23_port, B(22) => RALUOUT2_OUT_22_port,
                           B(21) => RALUOUT2_OUT_21_port, B(20) => 
                           RALUOUT2_OUT_20_port, B(19) => RALUOUT2_OUT_19_port,
                           B(18) => RALUOUT2_OUT_18_port, B(17) => 
                           RALUOUT2_OUT_17_port, B(16) => RALUOUT2_OUT_16_port,
                           B(15) => RALUOUT2_OUT_15_port, B(14) => 
                           RALUOUT2_OUT_14_port, B(13) => RALUOUT2_OUT_13_port,
                           B(12) => RALUOUT2_OUT_12_port, B(11) => 
                           RALUOUT2_OUT_11_port, B(10) => RALUOUT2_OUT_10_port,
                           B(9) => RALUOUT2_OUT_9_port, B(8) => 
                           RALUOUT2_OUT_8_port, B(7) => RALUOUT2_OUT_7_port, 
                           B(6) => RALUOUT2_OUT_6_port, B(5) => 
                           RALUOUT2_OUT_5_port, B(4) => RALUOUT2_OUT_4_port, 
                           B(3) => RALUOUT2_OUT_3_port, B(2) => 
                           RALUOUT2_OUT_2_port, B(1) => RALUOUT2_OUT_1_port, 
                           B(0) => RALUOUT2_OUT_0_port, SEL => WB_MUX_SEL, 
                           Y(31) => MUXC_OUT_31_port, Y(30) => MUXC_OUT_30_port
                           , Y(29) => MUXC_OUT_29_port, Y(28) => 
                           MUXC_OUT_28_port, Y(27) => MUXC_OUT_27_port, Y(26) 
                           => MUXC_OUT_26_port, Y(25) => MUXC_OUT_25_port, 
                           Y(24) => MUXC_OUT_24_port, Y(23) => MUXC_OUT_23_port
                           , Y(22) => MUXC_OUT_22_port, Y(21) => 
                           MUXC_OUT_21_port, Y(20) => MUXC_OUT_20_port, Y(19) 
                           => MUXC_OUT_19_port, Y(18) => MUXC_OUT_18_port, 
                           Y(17) => MUXC_OUT_17_port, Y(16) => MUXC_OUT_16_port
                           , Y(15) => MUXC_OUT_15_port, Y(14) => 
                           MUXC_OUT_14_port, Y(13) => MUXC_OUT_13_port, Y(12) 
                           => MUXC_OUT_12_port, Y(11) => MUXC_OUT_11_port, 
                           Y(10) => MUXC_OUT_10_port, Y(9) => MUXC_OUT_9_port, 
                           Y(8) => MUXC_OUT_8_port, Y(7) => MUXC_OUT_7_port, 
                           Y(6) => MUXC_OUT_6_port, Y(5) => MUXC_OUT_5_port, 
                           Y(4) => MUXC_OUT_4_port, Y(3) => MUXC_OUT_3_port, 
                           Y(2) => MUXC_OUT_2_port, Y(1) => MUXC_OUT_1_port, 
                           Y(0) => MUXC_OUT_0_port);
   reg_OUT : reg_NUMBIT32_1 port map( clk => CLK, en => ROUT_LATCH_EN, rst => 
                           RST, d(31) => MUXC_OUT_31_port, d(30) => 
                           MUXC_OUT_30_port, d(29) => MUXC_OUT_29_port, d(28) 
                           => MUXC_OUT_28_port, d(27) => MUXC_OUT_27_port, 
                           d(26) => MUXC_OUT_26_port, d(25) => MUXC_OUT_25_port
                           , d(24) => MUXC_OUT_24_port, d(23) => 
                           MUXC_OUT_23_port, d(22) => MUXC_OUT_22_port, d(21) 
                           => MUXC_OUT_21_port, d(20) => MUXC_OUT_20_port, 
                           d(19) => MUXC_OUT_19_port, d(18) => MUXC_OUT_18_port
                           , d(17) => MUXC_OUT_17_port, d(16) => 
                           MUXC_OUT_16_port, d(15) => MUXC_OUT_15_port, d(14) 
                           => MUXC_OUT_14_port, d(13) => MUXC_OUT_13_port, 
                           d(12) => MUXC_OUT_12_port, d(11) => MUXC_OUT_11_port
                           , d(10) => MUXC_OUT_10_port, d(9) => MUXC_OUT_9_port
                           , d(8) => MUXC_OUT_8_port, d(7) => MUXC_OUT_7_port, 
                           d(6) => MUXC_OUT_6_port, d(5) => MUXC_OUT_5_port, 
                           d(4) => MUXC_OUT_4_port, d(3) => MUXC_OUT_3_port, 
                           d(2) => MUXC_OUT_2_port, d(1) => MUXC_OUT_1_port, 
                           d(0) => MUXC_OUT_0_port, q(31) => Data_out(31), 
                           q(30) => Data_out(30), q(29) => Data_out(29), q(28) 
                           => Data_out(28), q(27) => Data_out(27), q(26) => 
                           Data_out(26), q(25) => Data_out(25), q(24) => 
                           Data_out(24), q(23) => Data_out(23), q(22) => 
                           Data_out(22), q(21) => Data_out(21), q(20) => 
                           Data_out(20), q(19) => Data_out(19), q(18) => 
                           Data_out(18), q(17) => Data_out(17), q(16) => 
                           Data_out(16), q(15) => Data_out(15), q(14) => 
                           Data_out(14), q(13) => Data_out(13), q(12) => 
                           Data_out(12), q(11) => Data_out(11), q(10) => 
                           Data_out(10), q(9) => Data_out(9), q(8) => 
                           Data_out(8), q(7) => Data_out(7), q(6) => 
                           Data_out(6), q(5) => Data_out(5), q(4) => 
                           Data_out(4), q(3) => Data_out(3), q(2) => 
                           Data_out(2), q(1) => Data_out(1), q(0) => 
                           Data_out(0));
   mux_WRaddr : MUX21_GENERIC_N5 port map( A(4) => X_Logic1_port, A(3) => 
                           X_Logic1_port, A(2) => X_Logic1_port, A(1) => 
                           X_Logic1_port, A(0) => X_Logic1_port, B(4) => n200, 
                           B(3) => n201, B(2) => RD3_OUT_2_port, B(1) => 
                           RD3_OUT_1_port, B(0) => n202, SEL => JandL, Y(4) => 
                           MUX_WRaddr_OUT_4_port, Y(3) => MUX_WRaddr_OUT_3_port
                           , Y(2) => MUX_WRaddr_OUT_2_port, Y(1) => 
                           MUX_WRaddr_OUT_1_port, Y(0) => MUX_WRaddr_OUT_0_port
                           );
   mux_WRdata : MUX21_GENERIC_N32_1 port map( A(31) => RPCplus8_OUT_31_port, 
                           A(30) => RPCplus8_OUT_30_port, A(29) => 
                           RPCplus8_OUT_29_port, A(28) => RPCplus8_OUT_28_port,
                           A(27) => RPCplus8_OUT_27_port, A(26) => 
                           RPCplus8_OUT_26_port, A(25) => RPCplus8_OUT_25_port,
                           A(24) => RPCplus8_OUT_24_port, A(23) => 
                           RPCplus8_OUT_23_port, A(22) => RPCplus8_OUT_22_port,
                           A(21) => RPCplus8_OUT_21_port, A(20) => 
                           RPCplus8_OUT_20_port, A(19) => RPCplus8_OUT_19_port,
                           A(18) => RPCplus8_OUT_18_port, A(17) => 
                           RPCplus8_OUT_17_port, A(16) => RPCplus8_OUT_16_port,
                           A(15) => RPCplus8_OUT_15_port, A(14) => 
                           RPCplus8_OUT_14_port, A(13) => RPCplus8_OUT_13_port,
                           A(12) => RPCplus8_OUT_12_port, A(11) => 
                           RPCplus8_OUT_11_port, A(10) => RPCplus8_OUT_10_port,
                           A(9) => RPCplus8_OUT_9_port, A(8) => 
                           RPCplus8_OUT_8_port, A(7) => RPCplus8_OUT_7_port, 
                           A(6) => RPCplus8_OUT_6_port, A(5) => 
                           RPCplus8_OUT_5_port, A(4) => RPCplus8_OUT_4_port, 
                           A(3) => RPCplus8_OUT_3_port, A(2) => 
                           RPCplus8_OUT_2_port, A(1) => RPCplus8_OUT_1_port, 
                           A(0) => RPCplus8_OUT_0_port, B(31) => 
                           MUXC_OUT_31_port, B(30) => MUXC_OUT_30_port, B(29) 
                           => MUXC_OUT_29_port, B(28) => MUXC_OUT_28_port, 
                           B(27) => MUXC_OUT_27_port, B(26) => MUXC_OUT_26_port
                           , B(25) => MUXC_OUT_25_port, B(24) => 
                           MUXC_OUT_24_port, B(23) => MUXC_OUT_23_port, B(22) 
                           => MUXC_OUT_22_port, B(21) => MUXC_OUT_21_port, 
                           B(20) => MUXC_OUT_20_port, B(19) => MUXC_OUT_19_port
                           , B(18) => MUXC_OUT_18_port, B(17) => 
                           MUXC_OUT_17_port, B(16) => MUXC_OUT_16_port, B(15) 
                           => MUXC_OUT_15_port, B(14) => MUXC_OUT_14_port, 
                           B(13) => MUXC_OUT_13_port, B(12) => MUXC_OUT_12_port
                           , B(11) => MUXC_OUT_11_port, B(10) => 
                           MUXC_OUT_10_port, B(9) => MUXC_OUT_9_port, B(8) => 
                           MUXC_OUT_8_port, B(7) => MUXC_OUT_7_port, B(6) => 
                           MUXC_OUT_6_port, B(5) => MUXC_OUT_5_port, B(4) => 
                           MUXC_OUT_4_port, B(3) => MUXC_OUT_3_port, B(2) => 
                           MUXC_OUT_2_port, B(1) => MUXC_OUT_1_port, B(0) => 
                           MUXC_OUT_0_port, SEL => JandL, Y(31) => 
                           MUX_WRdata_OUT_31_port, Y(30) => 
                           MUX_WRdata_OUT_30_port, Y(29) => 
                           MUX_WRdata_OUT_29_port, Y(28) => 
                           MUX_WRdata_OUT_28_port, Y(27) => 
                           MUX_WRdata_OUT_27_port, Y(26) => 
                           MUX_WRdata_OUT_26_port, Y(25) => 
                           MUX_WRdata_OUT_25_port, Y(24) => 
                           MUX_WRdata_OUT_24_port, Y(23) => 
                           MUX_WRdata_OUT_23_port, Y(22) => 
                           MUX_WRdata_OUT_22_port, Y(21) => 
                           MUX_WRdata_OUT_21_port, Y(20) => 
                           MUX_WRdata_OUT_20_port, Y(19) => 
                           MUX_WRdata_OUT_19_port, Y(18) => 
                           MUX_WRdata_OUT_18_port, Y(17) => 
                           MUX_WRdata_OUT_17_port, Y(16) => 
                           MUX_WRdata_OUT_16_port, Y(15) => 
                           MUX_WRdata_OUT_15_port, Y(14) => 
                           MUX_WRdata_OUT_14_port, Y(13) => 
                           MUX_WRdata_OUT_13_port, Y(12) => 
                           MUX_WRdata_OUT_12_port, Y(11) => 
                           MUX_WRdata_OUT_11_port, Y(10) => 
                           MUX_WRdata_OUT_10_port, Y(9) => 
                           MUX_WRdata_OUT_9_port, Y(8) => MUX_WRdata_OUT_8_port
                           , Y(7) => MUX_WRdata_OUT_7_port, Y(6) => 
                           MUX_WRdata_OUT_6_port, Y(5) => MUX_WRdata_OUT_5_port
                           , Y(4) => MUX_WRdata_OUT_4_port, Y(3) => 
                           MUX_WRdata_OUT_3_port, Y(2) => MUX_WRdata_OUT_2_port
                           , Y(1) => MUX_WRdata_OUT_1_port, Y(0) => 
                           MUX_WRdata_OUT_0_port);
   FORWARDING_UNIT_0 : ForwardingUnit_NUMBIT32_ADDRESS_WIDTH_RF5 port map( CLK 
                           => CLK, RST => RST, RS1(4) => RS1(4), RS1(3) => 
                           RS1(3), RS1(2) => RS1(2), RS1(1) => RS1(1), RS1(0) 
                           => RS1(0), RS2(4) => RS2(4), RS2(3) => RS2(3), 
                           RS2(2) => RS2(2), RS2(1) => RS2(1), RS2(0) => RS2(0)
                           , RD_XM(4) => RD2_OUT_4_port, RD_XM(3) => 
                           RD2_OUT_3_port, RD_XM(2) => RD2_OUT_2_port, RD_XM(1)
                           => RD2_OUT_1_port, RD_XM(0) => RD2_OUT_0_port, 
                           RD_MW(4) => RD3_OUT_4_port, RD_MW(3) => 
                           RD3_OUT_3_port, RD_MW(2) => RD3_OUT_2_port, RD_MW(1)
                           => RD3_OUT_1_port, RD_MW(0) => RD3_OUT_0_port, 
                           REGWRITE_XM => REGWRITE_XM, REGWRITE_MW => 
                           REGWRITE_MW, ForwardA(1) => ForwardA_1_port, 
                           ForwardA(0) => ForwardA_0_port, forwardB(1) => 
                           forwardB_1_port, forwardB(0) => forwardB_0_port, 
                           ForwardC => ForwardC, ForwardD(1) => ForwardD_1_port
                           , ForwardD(0) => ForwardD_0_port);
   U191 : OAI221_X2 port map( B1 => n50, B2 => n138, C1 => n51, C2 => n139, A 
                           => n156, ZN => ALU_inputA_24_port);
   U195 : OAI221_X2 port map( B1 => n47, B2 => n138, C1 => n48, C2 => n139, A 
                           => n155, ZN => ALU_inputA_25_port);
   U199 : OAI221_X2 port map( B1 => n44, B2 => n138, C1 => n45, C2 => n139, A 
                           => n154, ZN => ALU_inputA_26_port);
   U314 : INV_X1 port map( A => n101, ZN => n217);

end SYN_Struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity dlx_cu_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE29 is

   port( Clk, Rst, Flush_BTB, STALL : in std_logic;  IR_IN : in 
         std_logic_vector (31 downto 0);  IR_LATCH_EN, NPC_LATCH_EN, I_R_type, 
         REGF_LATCH_EN, RegA_LATCH_EN, RegB_LATCH_EN, RegIMM_LATCH_EN, 
         RegRD1_LATCH_EN, SIGN_UNSIGN, RFR1_EN, RFR2_EN, MUX_IMM_SEL, JUMP, 
         JUMP_EN, EQ_COND, MUXA_SEL, MUXB_SEL, ALU_OUTREG_EN, REGME_LATCH_EN, 
         RegRD2_LATCH_EN : out std_logic;  ALU_OPCODE : out std_logic_vector (0
         to 4);  DRAM_EN, DRAM_RE, DRAM_WE, LMD_LATCH_EN, RALUOUT2_LATCH_EN, 
         RegRD3_LATCH_EN, PC_LATCH_EN, RPCplus8_LATCH_EN, WB_MUX_SEL, RF_WE, 
         ROUT_LATCH_EN, JandL, REGWRITE_DX, REGWRITE_XM, REGWRITE_MW, 
         MEMREAD_DX : out std_logic);

end dlx_cu_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE29;

architecture SYN_dlx_cu_hw of 
   dlx_cu_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE29 is

   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component AND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X4
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal NPC_LATCH_EN_port, n205, RFR2_EN_port, MUXA_SEL_port, n206, 
      REGWRITE_MW_port, REGWRITE_DX_port, REGWRITE_XM_port, MEMREAD_DX_port, 
      cw_15_port, cw_14_port, cw_13_port, cw_8_port, cw_6_port, cw_5_port, cw_3
      , cw_2, cw_0, cw3_11, cw3_10, cw3_8_port, cw3_7_port, cw3_6_port, 
      cw3_5_port, cw3_3, cw3_0, cw4_3, cw4_0_port, aluOpcode_i_4_port, 
      aluOpcode_i_3_port, aluOpcode_i_2_port, aluOpcode_i_1_port, 
      aluOpcode_i_0_port, n30, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42
      , n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
      n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71
      , n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, 
      n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, 
      n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, 
      n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, 
      n124, n125, n126, n127, n128, n129, n131, n132, n133, n134, n135, n136, 
      n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, 
      n150, n151, n152, n153, n155, n156, n157, n158, n159, n160, n161, n162, 
      n163, n164, n165, n166, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n178, n179, n180, n1, n2, n130, n149, n154, n167, n177, n181, n182,
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, RegA_LATCH_EN_port, MUX_IMM_SEL_port, n207, n208, n209, n210,
      n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, 
      n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, 
      n235, n236, n238, n239 : std_logic;

begin
   IR_LATCH_EN <= NPC_LATCH_EN_port;
   NPC_LATCH_EN <= NPC_LATCH_EN_port;
   RegA_LATCH_EN <= RegA_LATCH_EN_port;
   RegB_LATCH_EN <= RFR2_EN_port;
   RegRD1_LATCH_EN <= cw_5_port;
   RFR2_EN <= RFR2_EN_port;
   MUX_IMM_SEL <= MUX_IMM_SEL_port;
   MUXA_SEL <= MUXA_SEL_port;
   RF_WE <= REGWRITE_MW_port;
   REGWRITE_DX <= REGWRITE_DX_port;
   REGWRITE_XM <= REGWRITE_XM_port;
   REGWRITE_MW <= REGWRITE_MW_port;
   MEMREAD_DX <= MEMREAD_DX_port;
   
   aluOpcode3_reg_4_inst : DFFS_X1 port map( D => aluOpcode_i_4_port, CK => Clk
                           , SN => n238, Q => ALU_OPCODE(0), QN => n33);
   aluOpcode3_reg_1_inst : DFFS_X1 port map( D => aluOpcode_i_1_port, CK => Clk
                           , SN => n238, Q => ALU_OPCODE(3), QN => n30);
   ROUT_LATCH_EN <= '0';
   U4 : AND2_X1 port map( A1 => n34, A2 => n35, ZN => cw_2);
   U5 : NOR2_X1 port map( A1 => n36, A2 => n192, ZN => cw_6_port);
   U6 : NOR2_X1 port map( A1 => n38, A2 => n192, ZN => cw_13_port);
   U7 : OR2_X1 port map( A1 => cw_3, A2 => cw_8_port, ZN => cw_14_port);
   U8 : NOR2_X1 port map( A1 => n192, A2 => n39, ZN => cw_3);
   U9 : OAI211_X1 port map( C1 => n185, C2 => n40, A => n41, B => n42, ZN => 
                           aluOpcode_i_4_port);
   U10 : OAI21_X1 port map( B1 => n43, B2 => n44, A => n183, ZN => n41);
   U11 : NAND4_X1 port map( A1 => n46, A2 => n47, A3 => n48, A4 => n49, ZN => 
                           aluOpcode_i_3_port);
   U12 : OAI211_X1 port map( C1 => n50, C2 => n181, A => n154, B => IR_IN(29), 
                           ZN => n48);
   U13 : AND2_X1 port map( A1 => n194, A2 => n53, ZN => n50);
   U14 : OAI21_X1 port map( B1 => n54, B2 => n55, A => n56, ZN => n47);
   U15 : INV_X1 port map( A => n57, ZN => n55);
   U16 : NOR4_X1 port map( A1 => IR_IN(4), A2 => IR_IN(2), A3 => n58, A4 => n59
                           , ZN => n54);
   U17 : INV_X1 port map( A => n60, ZN => n46);
   U18 : NAND4_X1 port map( A1 => n61, A2 => n62, A3 => n63, A4 => n64, ZN => 
                           aluOpcode_i_2_port);
   U19 : AOI21_X1 port map( B1 => n56, B2 => n65, A => n60, ZN => n64);
   U20 : OAI211_X1 port map( C1 => n66, C2 => n67, A => n68, B => n69, ZN => 
                           n60);
   U21 : NAND3_X1 port map( A1 => n70, A2 => n71, A3 => n57, ZN => n65);
   U22 : AOI22_X1 port map( A1 => IR_IN(5), A2 => n72, B1 => IR_IN(2), B2 => 
                           n73, ZN => n57);
   U23 : NAND4_X1 port map( A1 => n74, A2 => IR_IN(2), A3 => n75, A4 => n76, ZN
                           => n70);
   U24 : OAI211_X1 port map( C1 => n77, C2 => n181, A => IR_IN(28), B => n78, 
                           ZN => n63);
   U25 : NOR2_X1 port map( A1 => IR_IN(31), A2 => IR_IN(29), ZN => n77);
   U26 : NAND4_X1 port map( A1 => n42, A2 => n79, A3 => n80, A4 => n81, ZN => 
                           aluOpcode_i_1_port);
   U28 : NOR3_X1 port map( A1 => n86, A2 => n154, A3 => n194, ZN => n85);
   U29 : NOR2_X1 port map( A1 => IR_IN(28), A2 => n181, ZN => n82);
   U30 : OAI21_X1 port map( B1 => n44, B2 => n87, A => n183, ZN => n79);
   U31 : NAND2_X1 port map( A1 => n88, A2 => n89, ZN => n87);
   U32 : OAI211_X1 port map( C1 => n90, C2 => n91, A => IR_IN(2), B => n74, ZN 
                           => n88);
   U33 : NOR2_X1 port map( A1 => IR_IN(5), A2 => n92, ZN => n90);
   U34 : OAI211_X1 port map( C1 => IR_IN(5), C2 => n93, A => n94, B => n95, ZN 
                           => n44);
   U35 : AOI211_X1 port map( C1 => n96, C2 => IR_IN(2), A => n97, B => n98, ZN 
                           => n95);
   U36 : NOR3_X1 port map( A1 => n99, A2 => IR_IN(2), A3 => IR_IN(1), ZN => n97
                           );
   U37 : NOR2_X1 port map( A1 => n100, A2 => n92, ZN => n96);
   U38 : AOI21_X1 port map( B1 => IR_IN(5), B2 => IR_IN(0), A => IR_IN(3), ZN 
                           => n100);
   U39 : AOI211_X1 port map( C1 => IR_IN(0), C2 => n92, A => n101, B => 
                           IR_IN(3), ZN => n93);
   U40 : INV_X1 port map( A => n102, ZN => n42);
   U41 : OAI222_X1 port map( A1 => n154, A2 => n103, B1 => n190, B2 => n105, C1
                           => n106, C2 => n40, ZN => n102);
   U43 : AOI21_X1 port map( B1 => n154, B2 => IR_IN(28), A => IR_IN(27), ZN => 
                           n110);
   U44 : AOI22_X1 port map( A1 => n111, A2 => n2, B1 => n112, B2 => n185, ZN =>
                           n105);
   U45 : NAND2_X1 port map( A1 => n113, A2 => IR_IN(28), ZN => n111);
   U46 : AOI21_X1 port map( B1 => n114, B2 => n2, A => n115, ZN => n103);
   U47 : NOR3_X1 port map( A1 => n184, A2 => n194, A3 => n53, ZN => n115);
   U48 : NOR2_X1 port map( A1 => IR_IN(31), A2 => IR_IN(26), ZN => n53);
   U49 : NAND3_X1 port map( A1 => n117, A2 => n113, A3 => n194, ZN => n114);
   U50 : INV_X1 port map( A => n118, ZN => n113);
   U51 : OAI211_X1 port map( C1 => n119, C2 => n2, A => n80, B => n120, ZN => 
                           aluOpcode_i_0_port);
   U52 : AOI21_X1 port map( B1 => n56, B2 => n121, A => n122, ZN => n120);
   U53 : NAND4_X1 port map( A1 => n71, A2 => n123, A3 => n124, A4 => n125, ZN 
                           => n121);
   U54 : AOI22_X1 port map( A1 => IR_IN(2), A2 => n126, B1 => n73, B2 => 
                           IR_IN(0), ZN => n125);
   U55 : NOR3_X1 port map( A1 => n59, A2 => IR_IN(4), A3 => n75, ZN => n73);
   U56 : OAI33_X1 port map( A1 => n75, A2 => n98, A3 => n76, B1 => n127, B2 => 
                           IR_IN(0), B3 => n128, ZN => n126);
   U57 : NAND2_X1 port map( A1 => n92, A2 => n58, ZN => n127);
   U58 : INV_X1 port map( A => IR_IN(1), ZN => n92);
   U59 : NOR2_X1 port map( A1 => n99, A2 => IR_IN(3), ZN => n98);
   U60 : INV_X1 port map( A => n91, ZN => n75);
   U61 : NOR2_X1 port map( A1 => n58, A2 => IR_IN(1), ZN => n91);
   U62 : NAND4_X1 port map( A1 => n74, A2 => IR_IN(1), A3 => IR_IN(5), A4 => 
                           n101, ZN => n124);
   U63 : OR3_X1 port map( A1 => n58, A2 => n76, A3 => n89, ZN => n123);
   U64 : NAND4_X1 port map( A1 => n129, A2 => IR_IN(2), A3 => IR_IN(1), A4 => 
                           n58, ZN => n71);
   U65 : INV_X1 port map( A => IR_IN(5), ZN => n58);
   U66 : AND2_X1 port map( A1 => n94, A2 => n183, ZN => n56);
   U67 : AND3_X1 port map( A1 => n62, A2 => n49, A3 => n69, ZN => n80);
   U68 : AOI221_X1 port map( B1 => n167, B2 => n189, C1 => n118, C2 => n131, A 
                           => n132, ZN => n119);
   U69 : NOR3_X1 port map( A1 => n194, A2 => n185, A3 => n66, ZN => n132);
   U70 : NOR2_X1 port map( A1 => n133, A2 => n109, ZN => n118);
   U71 : AOI21_X1 port map( B1 => n134, B2 => n135, A => n187, ZN => 
                           SIGN_UNSIGN);
   U73 : INV_X1 port map( A => n139, ZN => n138);
   U74 : OAI22_X1 port map( A1 => n140, A2 => n141, B1 => IR_IN(26), B2 => n86,
                           ZN => n137);
   U75 : NAND3_X1 port map( A1 => IR_IN(5), A2 => n142, A3 => n94, ZN => n136);
   U76 : NOR3_X1 port map( A1 => IR_IN(6), A2 => IR_IN(10), A3 => n143, ZN => 
                           n94);
   U77 : OR3_X1 port map( A1 => IR_IN(9), A2 => IR_IN(8), A3 => IR_IN(7), ZN =>
                           n143);
   U78 : INV_X1 port map( A => n144, ZN => n142);
   U79 : AOI211_X1 port map( C1 => n101, C2 => n129, A => n72, B => n43, ZN => 
                           n144);
   U80 : NOR4_X1 port map( A1 => n59, A2 => n101, A3 => n99, A4 => IR_IN(1), ZN
                           => n43);
   U81 : INV_X1 port map( A => IR_IN(3), ZN => n59);
   U82 : NOR2_X1 port map( A1 => n89, A2 => n99, ZN => n72);
   U83 : INV_X1 port map( A => IR_IN(4), ZN => n99);
   U84 : NAND3_X1 port map( A1 => IR_IN(1), A2 => n101, A3 => IR_IN(3), ZN => 
                           n89);
   U85 : NOR2_X1 port map( A1 => n128, A2 => n76, ZN => n129);
   U86 : INV_X1 port map( A => IR_IN(0), ZN => n76);
   U87 : INV_X1 port map( A => n74, ZN => n128);
   U88 : NOR2_X1 port map( A1 => IR_IN(3), A2 => IR_IN(4), ZN => n74);
   U89 : INV_X1 port map( A => IR_IN(2), ZN => n101);
   U90 : NOR3_X1 port map( A1 => n145, A2 => n146, A3 => n196, ZN => n134);
   U91 : AOI21_X1 port map( B1 => n39, B2 => n36, A => n192, ZN => cw_5_port);
   U92 : AND2_X1 port map( A1 => n148, A2 => n177, ZN => n36);
   U93 : NOR2_X1 port map( A1 => n150, A2 => n192, ZN => RegIMM_LATCH_EN);
   U94 : OR2_X1 port map( A1 => cw_8_port, A2 => cw_15_port, ZN => RFR2_EN_port
                           );
   U95 : AND2_X1 port map( A1 => n183, A2 => n35, ZN => cw_15_port);
   U96 : NOR2_X1 port map( A1 => n139, A2 => n192, ZN => cw_8_port);
   U97 : OR2_X1 port map( A1 => n151, A2 => n239, ZN => n206);
   U98 : AOI21_X1 port map( B1 => n152, B2 => n150, A => STALL, ZN => n151);
   U99 : NOR2_X1 port map( A1 => n34, A2 => n153, ZN => n150);
   U100 : NAND3_X1 port map( A1 => n188, A2 => n155, A3 => n148, ZN => n34);
   U104 : NOR2_X1 port map( A1 => n159, A2 => n183, ZN => n148);
   U105 : NOR4_X1 port map( A1 => n133, A2 => n131, A3 => IR_IN(26), A4 => 
                           IR_IN(29), ZN => n45);
   U106 : OR2_X1 port map( A1 => n160, A2 => MUXA_SEL_port, ZN => JUMP_EN);
   U108 : NAND3_X1 port map( A1 => n161, A2 => n155, A3 => n156, ZN => n145);
   U109 : NAND4_X1 port map( A1 => n181, A2 => IR_IN(28), A3 => n2, A4 => n190,
                           ZN => n156);
   U110 : INV_X1 port map( A => n186, ZN => n35);
   U111 : AOI21_X1 port map( B1 => n162, B2 => n157, A => n186, ZN => n160);
   U112 : OAI21_X1 port map( B1 => n163, B2 => n187, A => n164, ZN => JUMP);
   U113 : INV_X1 port map( A => cw_0, ZN => n164);
   U114 : AOI21_X1 port map( B1 => n162, B2 => n155, A => n187, ZN => cw_0);
   U115 : NOR2_X1 port map( A1 => n165, A2 => n192, ZN => I_R_type);
   U116 : NOR4_X1 port map( A1 => n166, A2 => n159, A3 => n158, A4 => n153, ZN 
                           => n165);
   U117 : OAI211_X1 port map( C1 => n133, C2 => n193, A => n139, B => n163, ZN 
                           => n153);
   U118 : AND2_X1 port map( A1 => n161, A2 => n157, ZN => n163);
   U119 : NAND2_X1 port map( A1 => n78, A2 => n168, ZN => n157);
   U120 : NAND2_X1 port map( A1 => n169, A2 => n168, ZN => n161);
   U121 : NAND2_X1 port map( A1 => n170, A2 => n171, ZN => n139);
   U123 : INV_X1 port map( A => n147, ZN => n172);
   U124 : OAI211_X1 port map( C1 => n140, C2 => n173, A => n49, B => n39, ZN =>
                           n147);
   U125 : NAND4_X1 port map( A1 => IR_IN(31), A2 => IR_IN(27), A3 => n171, A4 
                           => n2, ZN => n39);
   U126 : NOR2_X1 port map( A1 => n109, A2 => n131, ZN => n171);
   U127 : INV_X1 port map( A => n108, ZN => n131);
   U128 : NOR2_X1 port map( A1 => IR_IN(30), A2 => IR_IN(28), ZN => n108);
   U130 : NAND2_X1 port map( A1 => n168, A2 => n174, ZN => n162);
   U132 : NAND4_X1 port map( A1 => n191, A2 => n62, A3 => n68, A4 => n69, ZN =>
                           n176);
   U133 : NAND3_X1 port map( A1 => n174, A2 => n194, A3 => n170, ZN => n69);
   U134 : NAND3_X1 port map( A1 => n78, A2 => n194, A3 => n170, ZN => n68);
   U136 : INV_X1 port map( A => IR_IN(31), ZN => n40);
   U137 : NAND3_X1 port map( A1 => n195, A2 => n174, A3 => n83, ZN => n62);
   U140 : OAI211_X1 port map( C1 => n66, C2 => n86, A => n61, B => n67, ZN => 
                           n146);
   U141 : NAND2_X1 port map( A1 => n112, A2 => n181, ZN => n67);
   U142 : NAND3_X1 port map( A1 => n112, A2 => n195, A3 => n169, ZN => n61);
   U143 : OAI22_X1 port map( A1 => n173, A2 => n178, B1 => n179, B2 => n66, ZN 
                           => n175);
   U144 : INV_X1 port map( A => n174, ZN => n66);
   U146 : INV_X1 port map( A => IR_IN(26), ZN => n109);
   U147 : AOI21_X1 port map( B1 => n195, B2 => n83, A => n180, ZN => n178);
   U148 : INV_X1 port map( A => n179, ZN => n180);
   U149 : NAND2_X1 port map( A1 => n112, A2 => n184, ZN => n179);
   U152 : INV_X1 port map( A => n78, ZN => n173);
   U154 : NAND2_X1 port map( A1 => n140, A2 => n86, ZN => n159);
   U155 : NAND2_X1 port map( A1 => IR_IN(29), A2 => n51, ZN => n86);
   U156 : NAND2_X1 port map( A1 => IR_IN(29), A2 => n167, ZN => n140);
   U158 : INV_X1 port map( A => n155, ZN => n166);
   U159 : NAND3_X1 port map( A1 => IR_IN(26), A2 => n104, A3 => n168, ZN => 
                           n155);
   U160 : NOR2_X1 port map( A1 => n117, A2 => IR_IN(29), ZN => n168);
   U163 : INV_X1 port map( A => IR_IN(27), ZN => n116);
   U164 : INV_X1 port map( A => IR_IN(30), ZN => n104);
   U165 : NOR4_X1 port map( A1 => n186, A2 => n133, A3 => n193, A4 => n141, ZN 
                           => EQ_COND);
   U166 : INV_X1 port map( A => n169, ZN => n141);
   U167 : NOR2_X1 port map( A1 => IR_IN(30), A2 => IR_IN(26), ZN => n169);
   U169 : NOR2_X1 port map( A1 => n194, A2 => IR_IN(29), ZN => n83);
   U170 : INV_X1 port map( A => IR_IN(28), ZN => n52);
   U171 : INV_X1 port map( A => n51, ZN => n133);
   U172 : NOR2_X1 port map( A1 => IR_IN(31), A2 => IR_IN(27), ZN => n51);
   U174 : INV_X1 port map( A => Flush_BTB, ZN => n152);
   U27 : INV_X1 port map( A => n107, ZN => n1);
   U42 : INV_X1 port map( A => n1, ZN => n2);
   U72 : AOI221_X1 port map( B1 => n154, B2 => n2, C1 => n108, C2 => n109, A =>
                           n110, ZN => n106);
   U101 : CLKBUF_X3 port map( A => n206, Z => PC_LATCH_EN);
   U102 : INV_X1 port map( A => IR_IN(29), ZN => n107);
   U103 : AND2_X1 port map( A1 => IR_IN(30), A2 => n130, ZN => n78);
   U107 : INV_X1 port map( A => IR_IN(26), ZN => n130);
   U122 : NOR3_X2 port map( A1 => n40, A2 => n184, A3 => n107, ZN => n170);
   U129 : NOR2_X2 port map( A1 => n109, A2 => n189, ZN => n174);
   U131 : INV_X1 port map( A => IR_IN(30), ZN => n149);
   U135 : INV_X1 port map( A => n149, ZN => n154);
   U138 : AND2_X2 port map( A1 => n84, A2 => n52, ZN => n167);
   U139 : INV_X4 port map( A => n167, ZN => n117);
   U145 : AOI221_X1 port map( B1 => n82, B2 => n78, C1 => n83, C2 => n195, A =>
                           n85, ZN => n81);
   U150 : NOR3_X1 port map( A1 => n175, A2 => n146, A3 => n176, ZN => n177);
   U151 : BUF_X1 port map( A => n51, Z => n181);
   U153 : INV_X1 port map( A => n45, ZN => n182);
   U157 : INV_X1 port map( A => n182, ZN => n183);
   U161 : AOI211_X4 port map( C1 => n183, C2 => n136, A => n137, B => n138, ZN 
                           => n135);
   U162 : INV_X1 port map( A => IR_IN(27), ZN => n184);
   U168 : INV_X1 port map( A => n184, ZN => n185);
   U173 : NAND2_X1 port map( A1 => NPC_LATCH_EN_port, A2 => n152, ZN => n187);
   U175 : NAND2_X1 port map( A1 => NPC_LATCH_EN_port, A2 => n152, ZN => n186);
   U176 : NOR2_X4 port map( A1 => n239, A2 => STALL, ZN => NPC_LATCH_EN_port);
   U177 : NAND2_X1 port map( A1 => NPC_LATCH_EN_port, A2 => n152, ZN => n37);
   U178 : AND3_X2 port map( A1 => n177, A2 => n162, A3 => n172, ZN => n188);
   U179 : INV_X4 port map( A => n188, ZN => n158);
   U180 : INV_X1 port map( A => n154, ZN => n190);
   U181 : INV_X1 port map( A => IR_IN(30), ZN => n189);
   U182 : AND2_X1 port map( A1 => IR_IN(29), A2 => IR_IN(28), ZN => n112);
   U183 : OR3_X2 port map( A1 => n173, A2 => n133, A3 => n193, ZN => n191);
   U184 : INV_X4 port map( A => n191, ZN => n122);
   U185 : CLKBUF_X1 port map( A => n186, Z => n192);
   U186 : OR2_X1 port map( A1 => n52, A2 => IR_IN(29), ZN => n193);
   U187 : INV_X1 port map( A => IR_IN(28), ZN => n194);
   U188 : BUF_X1 port map( A => n84, Z => n195);
   U189 : NOR2_X1 port map( A1 => n116, A2 => IR_IN(31), ZN => n84);
   U190 : CLKBUF_X1 port map( A => n147, Z => n196);
   U191 : CLKBUF_X1 port map( A => MUX_IMM_SEL_port, Z => RegA_LATCH_EN_port);
   U192 : OR2_X2 port map( A1 => n66, A2 => n140, ZN => n49);
   U193 : CLKBUF_X1 port map( A => RegA_LATCH_EN_port, Z => RFR1_EN);
   U194 : BUF_X4 port map( A => n205, Z => MUX_IMM_SEL_port);
   U195 : AOI21_X1 port map( B1 => n156, B2 => n38, A => n37, ZN => n205);
   U196 : AND4_X2 port map( A1 => n148, A2 => n188, A3 => n157, A4 => n139, ZN 
                           => n38);
   U197 : AND2_X4 port map( A1 => n35, A2 => n145, ZN => MUXA_SEL_port);
   cw5_reg_0_inst : DFFR_X1 port map( D => cw4_0_port, CK => Clk, RN => Rst, Q 
                           => JandL, QN => n236);
   cw5_reg_3_inst : DFFR_X1 port map( D => cw4_3, CK => Clk, RN => Rst, Q => 
                           WB_MUX_SEL, QN => n235);
   cw4_reg_11_inst : DFFR_X1 port map( D => cw3_11, CK => Clk, RN => Rst, Q => 
                           RPCplus8_LATCH_EN, QN => n234);
   cw4_reg_10_inst : DFFR_X1 port map( D => cw3_10, CK => Clk, RN => Rst, Q => 
                           DRAM_EN, QN => n233);
   cw4_reg_8_inst : DFFR_X1 port map( D => cw3_8_port, CK => Clk, RN => Rst, Q 
                           => DRAM_WE, QN => n232);
   cw4_reg_7_inst : DFFR_X1 port map( D => cw3_7_port, CK => Clk, RN => Rst, Q 
                           => LMD_LATCH_EN, QN => n231);
   cw4_reg_6_inst : DFFR_X1 port map( D => cw3_6_port, CK => Clk, RN => Rst, Q 
                           => RALUOUT2_LATCH_EN, QN => n230);
   cw4_reg_5_inst : DFFR_X1 port map( D => cw3_5_port, CK => Clk, RN => Rst, Q 
                           => RegRD3_LATCH_EN, QN => n229);
   cw4_reg_3_inst : DFFR_X1 port map( D => cw3_3, CK => Clk, RN => Rst, Q => 
                           cw4_3, QN => n228);
   cw4_reg_0_inst : DFFR_X1 port map( D => cw3_0, CK => Clk, RN => Rst, Q => 
                           cw4_0_port, QN => n227);
   cw4_reg_2_inst : DFFR_X1 port map( D => REGWRITE_DX_port, CK => Clk, RN => 
                           Rst, Q => REGWRITE_XM_port, QN => n226);
   cw4_reg_9_inst : DFFR_X1 port map( D => MEMREAD_DX_port, CK => Clk, RN => 
                           Rst, Q => DRAM_RE, QN => n225);
   cw5_reg_2_inst : DFFR_X1 port map( D => REGWRITE_XM_port, CK => Clk, RN => 
                           Rst, Q => REGWRITE_MW_port, QN => n224);
   aluOpcode3_reg_3_inst : DFFR_X1 port map( D => aluOpcode_i_3_port, CK => Clk
                           , RN => Rst, Q => ALU_OPCODE(1), QN => n223);
   aluOpcode3_reg_0_inst : DFFR_X1 port map( D => aluOpcode_i_0_port, CK => Clk
                           , RN => Rst, Q => ALU_OPCODE(4), QN => n222);
   aluOpcode3_reg_2_inst : DFFR_X1 port map( D => aluOpcode_i_2_port, CK => Clk
                           , RN => Rst, Q => ALU_OPCODE(2), QN => n221);
   cw3_reg_11_inst : DFFR_X1 port map( D => cw_0, CK => Clk, RN => Rst, Q => 
                           cw3_11, QN => n220);
   cw3_reg_0_inst : DFFR_X1 port map( D => cw_0, CK => Clk, RN => Rst, Q => 
                           cw3_0, QN => n219);
   cw3_reg_2_inst : DFFR_X1 port map( D => cw_2, CK => Clk, RN => Rst, Q => 
                           REGWRITE_DX_port, QN => n218);
   cw3_reg_15_inst : DFFR_X1 port map( D => cw_15_port, CK => Clk, RN => Rst, Q
                           => MUXB_SEL, QN => n217);
   cw3_reg_13_inst : DFFR_X1 port map( D => cw_13_port, CK => Clk, RN => Rst, Q
                           => ALU_OUTREG_EN, QN => n216);
   cw3_reg_6_inst : DFFR_X1 port map( D => cw_6_port, CK => Clk, RN => Rst, Q 
                           => cw3_6_port, QN => n215);
   cw3_reg_8_inst : DFFR_X1 port map( D => cw_8_port, CK => Clk, RN => Rst, Q 
                           => cw3_8_port, QN => n214);
   cw3_reg_12_inst : DFFR_X1 port map( D => cw_5_port, CK => Clk, RN => Rst, Q 
                           => RegRD2_LATCH_EN, QN => n213);
   cw3_reg_5_inst : DFFR_X1 port map( D => cw_5_port, CK => Clk, RN => Rst, Q 
                           => cw3_5_port, QN => n212);
   cw3_reg_9_inst : DFFR_X1 port map( D => cw_3, CK => Clk, RN => Rst, Q => 
                           MEMREAD_DX_port, QN => n211);
   cw3_reg_7_inst : DFFR_X1 port map( D => cw_3, CK => Clk, RN => Rst, Q => 
                           cw3_7_port, QN => n210);
   cw3_reg_3_inst : DFFR_X1 port map( D => cw_3, CK => Clk, RN => Rst, Q => 
                           cw3_3, QN => n209);
   cw3_reg_14_inst : DFFR_X1 port map( D => cw_14_port, CK => Clk, RN => Rst, Q
                           => REGME_LATCH_EN, QN => n208);
   cw3_reg_10_inst : DFFR_X1 port map( D => cw_14_port, CK => Clk, RN => Rst, Q
                           => cw3_10, QN => n207);
   U198 : INV_X1 port map( A => n239, ZN => REGF_LATCH_EN);
   U199 : INV_X1 port map( A => n239, ZN => n238);
   U200 : INV_X2 port map( A => Rst, ZN => n239);

end SYN_dlx_cu_hw;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity NPC_logic_PC_SIZE32 is

   port( Flush_BTB, BRANCH_CTRL_SIG, OUTT_NT_i : in std_logic;  PC_next, 
         BRANCH_ALU_OUT, OUT_PC_target_i, NPC : in std_logic_vector (31 downto 
         0);  PC_BUS : out std_logic_vector (31 downto 0));

end NPC_logic_PC_SIZE32;

architecture SYN_arch of NPC_logic_PC_SIZE32 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17, n18, n19, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32
      , n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, 
      n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61
      , n62, n63, n64, n65, n66, n67, n68, n69, n70, n20, n1, n71, n72, n73 : 
      std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => PC_BUS(9));
   U2 : AOI22_X1 port map( A1 => NPC(9), A2 => n73, B1 => BRANCH_ALU_OUT(9), B2
                           => n71, ZN => n3);
   U3 : AOI22_X1 port map( A1 => PC_next(9), A2 => n6, B1 => OUT_PC_target_i(9)
                           , B2 => n7, ZN => n2);
   U4 : NAND2_X1 port map( A1 => n8, A2 => n9, ZN => PC_BUS(8));
   U5 : AOI22_X1 port map( A1 => NPC(8), A2 => n73, B1 => BRANCH_ALU_OUT(8), B2
                           => n71, ZN => n9);
   U6 : AOI22_X1 port map( A1 => PC_next(8), A2 => n6, B1 => OUT_PC_target_i(8)
                           , B2 => n7, ZN => n8);
   U7 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => PC_BUS(7));
   U8 : AOI22_X1 port map( A1 => NPC(7), A2 => n73, B1 => BRANCH_ALU_OUT(7), B2
                           => n71, ZN => n11);
   U9 : AOI22_X1 port map( A1 => PC_next(7), A2 => n6, B1 => OUT_PC_target_i(7)
                           , B2 => n7, ZN => n10);
   U10 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => PC_BUS(6));
   U11 : AOI22_X1 port map( A1 => NPC(6), A2 => n73, B1 => BRANCH_ALU_OUT(6), 
                           B2 => n71, ZN => n13);
   U12 : AOI22_X1 port map( A1 => PC_next(6), A2 => n6, B1 => 
                           OUT_PC_target_i(6), B2 => n7, ZN => n12);
   U13 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => PC_BUS(5));
   U14 : AOI22_X1 port map( A1 => NPC(5), A2 => n73, B1 => BRANCH_ALU_OUT(5), 
                           B2 => n71, ZN => n15);
   U15 : AOI22_X1 port map( A1 => PC_next(5), A2 => n6, B1 => 
                           OUT_PC_target_i(5), B2 => n7, ZN => n14);
   U16 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => PC_BUS(4));
   U17 : AOI22_X1 port map( A1 => NPC(4), A2 => n73, B1 => BRANCH_ALU_OUT(4), 
                           B2 => n71, ZN => n17);
   U18 : AOI22_X1 port map( A1 => PC_next(4), A2 => n6, B1 => 
                           OUT_PC_target_i(4), B2 => n7, ZN => n16);
   U19 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => PC_BUS(3));
   U20 : AOI22_X1 port map( A1 => NPC(3), A2 => n73, B1 => BRANCH_ALU_OUT(3), 
                           B2 => n71, ZN => n19);
   U21 : AOI22_X1 port map( A1 => PC_next(3), A2 => n6, B1 => 
                           OUT_PC_target_i(3), B2 => n7, ZN => n18);
   U23 : AOI22_X1 port map( A1 => NPC(31), A2 => n73, B1 => BRANCH_ALU_OUT(31),
                           B2 => n71, ZN => n21);
   U25 : NAND2_X1 port map( A1 => n23, A2 => n22, ZN => PC_BUS(30));
   U26 : AOI22_X1 port map( A1 => NPC(30), A2 => n73, B1 => BRANCH_ALU_OUT(30),
                           B2 => n71, ZN => n23);
   U27 : AOI22_X1 port map( A1 => PC_next(30), A2 => n6, B1 => 
                           OUT_PC_target_i(30), B2 => n7, ZN => n22);
   U28 : NAND2_X1 port map( A1 => n24, A2 => n25, ZN => PC_BUS(2));
   U29 : AOI22_X1 port map( A1 => NPC(2), A2 => n73, B1 => BRANCH_ALU_OUT(2), 
                           B2 => n71, ZN => n25);
   U30 : AOI22_X1 port map( A1 => PC_next(2), A2 => n6, B1 => 
                           OUT_PC_target_i(2), B2 => n7, ZN => n24);
   U31 : NAND2_X1 port map( A1 => n26, A2 => n27, ZN => PC_BUS(29));
   U32 : AOI22_X1 port map( A1 => NPC(29), A2 => n73, B1 => BRANCH_ALU_OUT(29),
                           B2 => n71, ZN => n27);
   U33 : AOI22_X1 port map( A1 => PC_next(29), A2 => n6, B1 => 
                           OUT_PC_target_i(29), B2 => n7, ZN => n26);
   U34 : NAND2_X1 port map( A1 => n28, A2 => n29, ZN => PC_BUS(28));
   U35 : AOI22_X1 port map( A1 => NPC(28), A2 => n73, B1 => BRANCH_ALU_OUT(28),
                           B2 => n71, ZN => n29);
   U36 : AOI22_X1 port map( A1 => PC_next(28), A2 => n6, B1 => 
                           OUT_PC_target_i(28), B2 => n7, ZN => n28);
   U37 : NAND2_X1 port map( A1 => n30, A2 => n31, ZN => PC_BUS(27));
   U38 : AOI22_X1 port map( A1 => NPC(27), A2 => n73, B1 => BRANCH_ALU_OUT(27),
                           B2 => n71, ZN => n31);
   U39 : AOI22_X1 port map( A1 => PC_next(27), A2 => n6, B1 => 
                           OUT_PC_target_i(27), B2 => n7, ZN => n30);
   U40 : NAND2_X1 port map( A1 => n32, A2 => n33, ZN => PC_BUS(26));
   U41 : AOI22_X1 port map( A1 => NPC(26), A2 => n73, B1 => BRANCH_ALU_OUT(26),
                           B2 => n71, ZN => n33);
   U42 : AOI22_X1 port map( A1 => PC_next(26), A2 => n6, B1 => 
                           OUT_PC_target_i(26), B2 => n7, ZN => n32);
   U43 : NAND2_X1 port map( A1 => n34, A2 => n35, ZN => PC_BUS(25));
   U44 : AOI22_X1 port map( A1 => NPC(25), A2 => n73, B1 => BRANCH_ALU_OUT(25),
                           B2 => n71, ZN => n35);
   U45 : AOI22_X1 port map( A1 => PC_next(25), A2 => n6, B1 => 
                           OUT_PC_target_i(25), B2 => n7, ZN => n34);
   U46 : NAND2_X1 port map( A1 => n36, A2 => n37, ZN => PC_BUS(24));
   U47 : AOI22_X1 port map( A1 => NPC(24), A2 => n73, B1 => BRANCH_ALU_OUT(24),
                           B2 => n71, ZN => n37);
   U48 : AOI22_X1 port map( A1 => PC_next(24), A2 => n6, B1 => 
                           OUT_PC_target_i(24), B2 => n7, ZN => n36);
   U49 : NAND2_X1 port map( A1 => n38, A2 => n39, ZN => PC_BUS(23));
   U50 : AOI22_X1 port map( A1 => NPC(23), A2 => n73, B1 => BRANCH_ALU_OUT(23),
                           B2 => n71, ZN => n39);
   U51 : AOI22_X1 port map( A1 => PC_next(23), A2 => n6, B1 => 
                           OUT_PC_target_i(23), B2 => n7, ZN => n38);
   U52 : NAND2_X1 port map( A1 => n40, A2 => n41, ZN => PC_BUS(22));
   U53 : AOI22_X1 port map( A1 => NPC(22), A2 => n73, B1 => BRANCH_ALU_OUT(22),
                           B2 => n71, ZN => n41);
   U54 : AOI22_X1 port map( A1 => PC_next(22), A2 => n6, B1 => 
                           OUT_PC_target_i(22), B2 => n7, ZN => n40);
   U55 : NAND2_X1 port map( A1 => n42, A2 => n43, ZN => PC_BUS(21));
   U56 : AOI22_X1 port map( A1 => NPC(21), A2 => n73, B1 => BRANCH_ALU_OUT(21),
                           B2 => n71, ZN => n43);
   U57 : AOI22_X1 port map( A1 => PC_next(21), A2 => n6, B1 => 
                           OUT_PC_target_i(21), B2 => n7, ZN => n42);
   U58 : NAND2_X1 port map( A1 => n44, A2 => n45, ZN => PC_BUS(20));
   U59 : AOI22_X1 port map( A1 => NPC(20), A2 => n73, B1 => BRANCH_ALU_OUT(20),
                           B2 => n71, ZN => n45);
   U60 : AOI22_X1 port map( A1 => PC_next(20), A2 => n6, B1 => 
                           OUT_PC_target_i(20), B2 => n7, ZN => n44);
   U61 : NAND2_X1 port map( A1 => n46, A2 => n47, ZN => PC_BUS(1));
   U62 : AOI22_X1 port map( A1 => NPC(1), A2 => n73, B1 => BRANCH_ALU_OUT(1), 
                           B2 => n71, ZN => n47);
   U63 : AOI22_X1 port map( A1 => PC_next(1), A2 => n6, B1 => 
                           OUT_PC_target_i(1), B2 => n7, ZN => n46);
   U64 : NAND2_X1 port map( A1 => n49, A2 => n48, ZN => PC_BUS(19));
   U65 : AOI22_X1 port map( A1 => NPC(19), A2 => n73, B1 => BRANCH_ALU_OUT(19),
                           B2 => n71, ZN => n49);
   U66 : AOI22_X1 port map( A1 => PC_next(19), A2 => n6, B1 => 
                           OUT_PC_target_i(19), B2 => n7, ZN => n48);
   U67 : NAND2_X1 port map( A1 => n50, A2 => n51, ZN => PC_BUS(18));
   U68 : AOI22_X1 port map( A1 => NPC(18), A2 => n73, B1 => BRANCH_ALU_OUT(18),
                           B2 => n71, ZN => n51);
   U69 : AOI22_X1 port map( A1 => PC_next(18), A2 => n6, B1 => 
                           OUT_PC_target_i(18), B2 => n7, ZN => n50);
   U70 : NAND2_X1 port map( A1 => n52, A2 => n53, ZN => PC_BUS(17));
   U71 : AOI22_X1 port map( A1 => NPC(17), A2 => n73, B1 => BRANCH_ALU_OUT(17),
                           B2 => n71, ZN => n53);
   U72 : AOI22_X1 port map( A1 => PC_next(17), A2 => n6, B1 => 
                           OUT_PC_target_i(17), B2 => n7, ZN => n52);
   U73 : NAND2_X1 port map( A1 => n54, A2 => n55, ZN => PC_BUS(16));
   U74 : AOI22_X1 port map( A1 => NPC(16), A2 => n73, B1 => BRANCH_ALU_OUT(16),
                           B2 => n71, ZN => n55);
   U75 : AOI22_X1 port map( A1 => PC_next(16), A2 => n6, B1 => 
                           OUT_PC_target_i(16), B2 => n7, ZN => n54);
   U76 : NAND2_X1 port map( A1 => n56, A2 => n57, ZN => PC_BUS(15));
   U77 : AOI22_X1 port map( A1 => NPC(15), A2 => n73, B1 => BRANCH_ALU_OUT(15),
                           B2 => n71, ZN => n57);
   U78 : AOI22_X1 port map( A1 => PC_next(15), A2 => n6, B1 => 
                           OUT_PC_target_i(15), B2 => n7, ZN => n56);
   U79 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => PC_BUS(14));
   U80 : AOI22_X1 port map( A1 => NPC(14), A2 => n73, B1 => BRANCH_ALU_OUT(14),
                           B2 => n71, ZN => n59);
   U81 : AOI22_X1 port map( A1 => PC_next(14), A2 => n6, B1 => 
                           OUT_PC_target_i(14), B2 => n7, ZN => n58);
   U82 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => PC_BUS(13));
   U83 : AOI22_X1 port map( A1 => NPC(13), A2 => n73, B1 => BRANCH_ALU_OUT(13),
                           B2 => n71, ZN => n61);
   U84 : AOI22_X1 port map( A1 => PC_next(13), A2 => n6, B1 => 
                           OUT_PC_target_i(13), B2 => n7, ZN => n60);
   U85 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => PC_BUS(12));
   U86 : AOI22_X1 port map( A1 => NPC(12), A2 => n73, B1 => BRANCH_ALU_OUT(12),
                           B2 => n71, ZN => n63);
   U87 : AOI22_X1 port map( A1 => PC_next(12), A2 => n6, B1 => 
                           OUT_PC_target_i(12), B2 => n7, ZN => n62);
   U88 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => PC_BUS(11));
   U89 : AOI22_X1 port map( A1 => NPC(11), A2 => n73, B1 => BRANCH_ALU_OUT(11),
                           B2 => n71, ZN => n65);
   U90 : AOI22_X1 port map( A1 => PC_next(11), A2 => n6, B1 => 
                           OUT_PC_target_i(11), B2 => n7, ZN => n64);
   U91 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => PC_BUS(10));
   U92 : AOI22_X1 port map( A1 => NPC(10), A2 => n73, B1 => BRANCH_ALU_OUT(10),
                           B2 => n71, ZN => n67);
   U93 : AOI22_X1 port map( A1 => PC_next(10), A2 => n6, B1 => 
                           OUT_PC_target_i(10), B2 => n7, ZN => n66);
   U94 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => PC_BUS(0));
   U95 : AOI22_X1 port map( A1 => NPC(0), A2 => n73, B1 => BRANCH_ALU_OUT(0), 
                           B2 => n71, ZN => n69);
   U98 : AOI22_X1 port map( A1 => PC_next(0), A2 => n6, B1 => 
                           OUT_PC_target_i(0), B2 => n7, ZN => n68);
   U96 : AND2_X1 port map( A1 => BRANCH_CTRL_SIG, A2 => Flush_BTB, ZN => n5);
   U100 : INV_X1 port map( A => Flush_BTB, ZN => n70);
   U22 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => PC_BUS(31));
   U24 : AOI22_X1 port map( A1 => PC_next(31), A2 => n6, B1 => 
                           OUT_PC_target_i(31), B2 => n7, ZN => n20);
   U97 : INV_X1 port map( A => n5, ZN => n1);
   U99 : INV_X2 port map( A => n1, ZN => n71);
   U101 : NOR2_X4 port map( A1 => Flush_BTB, A2 => OUTT_NT_i, ZN => n6);
   U102 : AND2_X4 port map( A1 => OUTT_NT_i, A2 => n70, ZN => n7);
   U103 : INV_X1 port map( A => n4, ZN => n72);
   U104 : INV_X2 port map( A => n72, ZN => n73);
   U105 : NOR2_X1 port map( A1 => n70, A2 => BRANCH_CTRL_SIG, ZN => n4);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity DLX_IR_SIZE32_PC_SIZE32 is

   port( Clk, Rst : in std_logic;  Iaddr : out std_logic_vector (31 downto 0); 
         Idata : in std_logic_vector (31 downto 0);  Denable, Drd, Dwd : out 
         std_logic;  Daddr, Ddatain : out std_logic_vector (31 downto 0);  
         Ddataout : in std_logic_vector (31 downto 0);  DataOut : out 
         std_logic_vector (31 downto 0));

end DLX_IR_SIZE32_PC_SIZE32;

architecture SYN_dlx_rtl of DLX_IR_SIZE32_PC_SIZE32 is

   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X8
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLX_IR_SIZE32_PC_SIZE32_DW01_inc_1
      port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component HazardUnit_NUMBIT32_ADDRESS_WIDTH_RF5_OP_CODE_SIZE6
      port( CLK, RST : in std_logic;  RS1, RS2 : in std_logic_vector (4 downto 
            0);  REGWRITE_DX, MEMREAD_DX : in std_logic;  RD : in 
            std_logic_vector (4 downto 0);  OPCODE : in std_logic_vector (5 
            downto 0);  STALL : out std_logic);
   end component;
   
   component BTB_PC_SIZE32_BTBSIZE5
      port( Reset, Clk, Enable : in std_logic;  PC_read : in std_logic_vector 
            (31 downto 0);  WR : in std_logic;  PC_write : in std_logic_vector 
            (31 downto 0);  SetT_NT : in std_logic;  Set_target : in 
            std_logic_vector (31 downto 0);  OUT_PC_target : out 
            std_logic_vector (31 downto 0);  OUTT_NT, prevT_NT : out std_logic
            );
   end component;
   
   component datapath_NUMBIT32_ADDRESS_WIDTH_RF5_ADDRESS_WIDTH_DM32
      port( CLK, RST : in std_logic;  INP1 : in std_logic_vector (31 downto 0);
            INP2 : in std_logic_vector (15 downto 0);  IMM26 : in 
            std_logic_vector (25 downto 0);  RS1, RS2, RD : in std_logic_vector
            (4 downto 0);  REGF_LATCH_EN, RegA_LATCH_EN, RegB_LATCH_EN, 
            RegIMM_LATCH_EN, RegRD1_LATCH_EN, SIGN_UNSIGN, RFR1_EN, RFR2_EN, 
            MUX_IMM_SEL, JUMP, JUMP_EN, EQ_COND, MUXA_SEL, MUXB_SEL, 
            RALUOUT_LATCH_EN, REGME_LATCH_EN, RegRD2_LATCH_EN : in std_logic;  
            ALU_OPCODE : in std_logic_vector (0 to 4);  ADDR_DRAM, DATAIN_DRAM 
            : out std_logic_vector (31 downto 0);  DATAOUT_DRAM : in 
            std_logic_vector (31 downto 0);  LMD_LATCH_EN, RALUOUT2_LATCH_EN, 
            RegRD3_LATCH_EN, RPCplus8_LATCH_EN, WB_MUX_SEL, RF_WE, 
            ROUT_LATCH_EN, JandL : in std_logic;  BRANCH_CTRL_SIG : out 
            std_logic;  BRANCH_ALU_OUT, Data_out : out std_logic_vector (31 
            downto 0);  REGWRITE_XM, REGWRITE_MW : in std_logic);
   end component;
   
   component dlx_cu_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE29
      port( Clk, Rst, Flush_BTB, STALL : in std_logic;  IR_IN : in 
            std_logic_vector (31 downto 0);  IR_LATCH_EN, NPC_LATCH_EN, 
            I_R_type, REGF_LATCH_EN, RegA_LATCH_EN, RegB_LATCH_EN, 
            RegIMM_LATCH_EN, RegRD1_LATCH_EN, SIGN_UNSIGN, RFR1_EN, RFR2_EN, 
            MUX_IMM_SEL, JUMP, JUMP_EN, EQ_COND, MUXA_SEL, MUXB_SEL, 
            ALU_OUTREG_EN, REGME_LATCH_EN, RegRD2_LATCH_EN : out std_logic;  
            ALU_OPCODE : out std_logic_vector (0 to 4);  DRAM_EN, DRAM_RE, 
            DRAM_WE, LMD_LATCH_EN, RALUOUT2_LATCH_EN, RegRD3_LATCH_EN, 
            PC_LATCH_EN, RPCplus8_LATCH_EN, WB_MUX_SEL, RF_WE, ROUT_LATCH_EN, 
            JandL, REGWRITE_DX, REGWRITE_XM, REGWRITE_MW, MEMREAD_DX : out 
            std_logic);
   end component;
   
   component NPC_logic_PC_SIZE32
      port( Flush_BTB, BRANCH_CTRL_SIG, OUTT_NT_i : in std_logic;  PC_next, 
            BRANCH_ALU_OUT, OUT_PC_target_i, NPC : in std_logic_vector (31 
            downto 0);  PC_BUS : out std_logic_vector (31 downto 0));
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic1_port, Iaddr_31_port, Iaddr_30_port, Iaddr_29_port, 
      Iaddr_28_port, Iaddr_27_port, Iaddr_26_port, Iaddr_25_port, Iaddr_24_port
      , Iaddr_23_port, Iaddr_22_port, Iaddr_21_port, Iaddr_20_port, 
      Iaddr_19_port, Iaddr_18_port, Iaddr_17_port, Iaddr_16_port, Iaddr_15_port
      , Iaddr_14_port, Iaddr_13_port, Iaddr_12_port, Iaddr_11_port, 
      Iaddr_10_port, Iaddr_9_port, Iaddr_8_port, Iaddr_7_port, Iaddr_6_port, 
      Iaddr_5_port, Iaddr_4_port, Iaddr_3_port, Iaddr_2_port, Iaddr_1_port, 
      n314, INP2_15_port, INP2_14_port, INP2_13_port, INP2_12_port, 
      INP2_11_port, INP2_10_port, INP2_9_port, INP2_8_port, INP2_7_port, 
      INP2_6_port, INP2_5_port, INP2_4_port, INP2_3_port, INP2_2_port, 
      INP2_1_port, INP2_0_port, IR_31_port, IR_30_port, IR_29_port, IR_28_port,
      IR_27_port, IR_26_port, IMM26_25_port, IMM26_24_port, IMM26_23_port, 
      IMM26_22_port, IMM26_21_port, IMM26_20_port, IMM26_19_port, IMM26_18_port
      , IMM26_17_port, IMM26_16_port, I_R_TYPE_i, N2, RD_4_port, RD_3_port, 
      RD_2_port, RD_1_port, RD_0_port, prevT_NT_i, Flush_BTB_i, BRANCH_CTRL_SIG
      , Flush_BTB, IR_LATCH_EN_i, PC_LATCH_EN_i, PC_BUS_31_port, PC_BUS_30_port
      , PC_BUS_29_port, PC_BUS_28_port, PC_BUS_27_port, PC_BUS_26_port, 
      PC_BUS_25_port, PC_BUS_24_port, PC_BUS_23_port, PC_BUS_22_port, 
      PC_BUS_21_port, PC_BUS_20_port, PC_BUS_19_port, PC_BUS_18_port, 
      PC_BUS_17_port, PC_BUS_16_port, PC_BUS_15_port, PC_BUS_14_port, 
      PC_BUS_13_port, PC_BUS_12_port, PC_BUS_11_port, PC_BUS_10_port, 
      PC_BUS_9_port, PC_BUS_8_port, PC_BUS_7_port, PC_BUS_6_port, PC_BUS_5_port
      , PC_BUS_4_port, PC_BUS_3_port, PC_BUS_2_port, PC_BUS_1_port, 
      PC_BUS_0_port, NPC_31_port, NPC_30_port, NPC_29_port, NPC_28_port, 
      NPC_27_port, NPC_26_port, NPC_25_port, NPC_24_port, NPC_23_port, 
      NPC_22_port, NPC_21_port, NPC_20_port, NPC_19_port, NPC_18_port, 
      NPC_17_port, NPC_16_port, NPC_15_port, NPC_14_port, NPC_13_port, 
      NPC_12_port, NPC_11_port, NPC_10_port, NPC_9_port, NPC_8_port, NPC_7_port
      , NPC_6_port, NPC_5_port, NPC_4_port, NPC_3_port, NPC_2_port, NPC_1_port,
      NPC_0_port, NPC_LATCH_EN_i, PC_next_31_port, PC_next_30_port, 
      PC_next_29_port, PC_next_28_port, PC_next_27_port, PC_next_26_port, 
      PC_next_25_port, PC_next_24_port, PC_next_23_port, PC_next_22_port, 
      PC_next_21_port, PC_next_20_port, PC_next_19_port, PC_next_18_port, 
      PC_next_17_port, PC_next_16_port, PC_next_15_port, PC_next_14_port, 
      PC_next_13_port, PC_next_12_port, PC_next_11_port, PC_next_10_port, 
      PC_next_9_port, PC_next_8_port, PC_next_7_port, PC_next_6_port, 
      PC_next_5_port, PC_next_4_port, PC_next_3_port, PC_next_2_port, 
      PC_next_1_port, PC_next_0_port, OUTT_NT_i, BRANCH_ALU_OUT_31_port, 
      BRANCH_ALU_OUT_30_port, BRANCH_ALU_OUT_29_port, BRANCH_ALU_OUT_28_port, 
      BRANCH_ALU_OUT_27_port, BRANCH_ALU_OUT_26_port, BRANCH_ALU_OUT_25_port, 
      BRANCH_ALU_OUT_24_port, BRANCH_ALU_OUT_23_port, BRANCH_ALU_OUT_22_port, 
      BRANCH_ALU_OUT_21_port, BRANCH_ALU_OUT_20_port, BRANCH_ALU_OUT_19_port, 
      BRANCH_ALU_OUT_18_port, BRANCH_ALU_OUT_17_port, BRANCH_ALU_OUT_16_port, 
      BRANCH_ALU_OUT_15_port, BRANCH_ALU_OUT_14_port, BRANCH_ALU_OUT_13_port, 
      BRANCH_ALU_OUT_12_port, BRANCH_ALU_OUT_11_port, BRANCH_ALU_OUT_10_port, 
      BRANCH_ALU_OUT_9_port, BRANCH_ALU_OUT_8_port, BRANCH_ALU_OUT_7_port, 
      BRANCH_ALU_OUT_6_port, BRANCH_ALU_OUT_5_port, BRANCH_ALU_OUT_4_port, 
      BRANCH_ALU_OUT_3_port, BRANCH_ALU_OUT_2_port, BRANCH_ALU_OUT_1_port, 
      BRANCH_ALU_OUT_0_port, OUT_PC_target_i_31_port, OUT_PC_target_i_30_port, 
      OUT_PC_target_i_29_port, OUT_PC_target_i_28_port, OUT_PC_target_i_27_port
      , OUT_PC_target_i_26_port, OUT_PC_target_i_25_port, 
      OUT_PC_target_i_24_port, OUT_PC_target_i_23_port, OUT_PC_target_i_22_port
      , OUT_PC_target_i_21_port, OUT_PC_target_i_20_port, 
      OUT_PC_target_i_19_port, OUT_PC_target_i_18_port, OUT_PC_target_i_17_port
      , OUT_PC_target_i_16_port, OUT_PC_target_i_15_port, 
      OUT_PC_target_i_14_port, OUT_PC_target_i_13_port, OUT_PC_target_i_12_port
      , OUT_PC_target_i_11_port, OUT_PC_target_i_10_port, 
      OUT_PC_target_i_9_port, OUT_PC_target_i_8_port, OUT_PC_target_i_7_port, 
      OUT_PC_target_i_6_port, OUT_PC_target_i_5_port, OUT_PC_target_i_4_port, 
      OUT_PC_target_i_3_port, OUT_PC_target_i_2_port, OUT_PC_target_i_1_port, 
      OUT_PC_target_i_0_port, STALL_i, RegRF_LATCH_EN_i, RegA_LATCH_EN_i, 
      RegB_LATCH_EN_i, RegIMM_LATCH_EN_i, RegRD1_LATCH_EN_i, SIGN_UNSIGN_i, 
      RFR1_EN_i, RFR2_EN_i, MUX_IMM_SEL_i, JUMP_i, JUMP_EN_i, EQ_COND_i, 
      MUXA_SEL_i, MUXB_SEL_i, ALU_OUTREG_EN_i, REGME_LATCH_EN_i, 
      RegRD2_LATCH_EN_i, ALU_OPCODE_i_4_port, ALU_OPCODE_i_3_port, 
      ALU_OPCODE_i_2_port, ALU_OPCODE_i_1_port, ALU_OPCODE_i_0_port, 
      LMD_LATCH_EN_i, RALUOUT2_LATCH_EN_i, RegRD3_LATCH_EN_i, 
      RPCplus8_LATCH_EN_i, WB_MUX_SEL_i, RF_WE_i, ROUT_LATCH_EN_i, JandL_i, 
      REGWRITE_DX_i, REGWRITE_XM_i, REGWRITE_MW_i, MEMREAD_DX_i, N4, N5, 
      n2_port, n3, n4_port, n5_port, n6, n7, n8, n9, n10, n11, n12, n13, n14, 
      n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29
      , n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, 
      n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58
      , n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, 
      n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
      n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, 
      n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, 
      n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, 
      n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, 
      n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, 
      n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, 
      n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, 
      n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, 
      n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, 
      n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, 
      n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, 
      n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, 
      n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, 
      n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, 
      n294, n295, n296, Iaddr_0_port, n298, n299, n300, n301, n302, n303, n304,
      n305, n306, n307, n308, n309, n310, n311, n312, n313, n_1117 : std_logic;

begin
   Iaddr <= ( Iaddr_31_port, Iaddr_30_port, Iaddr_29_port, Iaddr_28_port, 
      Iaddr_27_port, Iaddr_26_port, Iaddr_25_port, Iaddr_24_port, Iaddr_23_port
      , Iaddr_22_port, Iaddr_21_port, Iaddr_20_port, Iaddr_19_port, 
      Iaddr_18_port, Iaddr_17_port, Iaddr_16_port, Iaddr_15_port, Iaddr_14_port
      , Iaddr_13_port, Iaddr_12_port, Iaddr_11_port, Iaddr_10_port, 
      Iaddr_9_port, Iaddr_8_port, Iaddr_7_port, Iaddr_6_port, Iaddr_5_port, 
      Iaddr_4_port, Iaddr_3_port, Iaddr_2_port, Iaddr_1_port, Iaddr_0_port );
   
   X_Logic1_port <= '1';
   C628 : AND2_X2 port map( A1 => prevT_NT_i, A2 => N4, ZN => N5);
   C627 : XOR2_X1 port map( A => N5, B => BRANCH_CTRL_SIG, Z => Flush_BTB);
   I_1 : INV_X2 port map( A => I_R_TYPE_i, ZN => N2);
   NPC_reg_0_inst : DFFR_X1 port map( D => n289, CK => Clk, RN => n311, Q => 
                           NPC_0_port, QN => n193);
   Flush_BTB_i_reg : DFFR_X1 port map( D => Flush_BTB, CK => Clk, RN => n313, Q
                           => Flush_BTB_i, QN => N4);
   PC_reg_0_inst : DFFR_X1 port map( D => n287, CK => Clk, RN => n313, Q => 
                           n314, QN => n191);
   PC_reg_1_inst : DFFR_X1 port map( D => n286, CK => Clk, RN => n312, Q => 
                           Iaddr_1_port, QN => n190);
   PC_reg_2_inst : DFFR_X1 port map( D => n285, CK => Clk, RN => n312, Q => 
                           Iaddr_2_port, QN => n189);
   PC_reg_3_inst : DFFR_X1 port map( D => n284, CK => Clk, RN => n313, Q => 
                           Iaddr_3_port, QN => n188);
   PC_reg_4_inst : DFFR_X1 port map( D => n283, CK => Clk, RN => n313, Q => 
                           Iaddr_4_port, QN => n187);
   PC_reg_5_inst : DFFR_X1 port map( D => n282, CK => Clk, RN => n313, Q => 
                           Iaddr_5_port, QN => n186);
   PC_reg_6_inst : DFFR_X1 port map( D => n281, CK => Clk, RN => n313, Q => 
                           Iaddr_6_port, QN => n185);
   PC_reg_7_inst : DFFR_X1 port map( D => n280, CK => Clk, RN => n313, Q => 
                           Iaddr_7_port, QN => n184);
   PC_reg_8_inst : DFFR_X1 port map( D => n279, CK => Clk, RN => n313, Q => 
                           Iaddr_8_port, QN => n183);
   PC_reg_9_inst : DFFR_X1 port map( D => n278, CK => Clk, RN => n313, Q => 
                           Iaddr_9_port, QN => n182);
   PC_reg_10_inst : DFFR_X1 port map( D => n277, CK => Clk, RN => n312, Q => 
                           Iaddr_10_port, QN => n181);
   PC_reg_11_inst : DFFR_X1 port map( D => n276, CK => Clk, RN => n311, Q => 
                           Iaddr_11_port, QN => n180);
   PC_reg_12_inst : DFFR_X1 port map( D => n275, CK => Clk, RN => n311, Q => 
                           Iaddr_12_port, QN => n179);
   PC_reg_13_inst : DFFR_X1 port map( D => n274, CK => Clk, RN => n311, Q => 
                           Iaddr_13_port, QN => n178);
   PC_reg_14_inst : DFFR_X1 port map( D => n273, CK => Clk, RN => n311, Q => 
                           Iaddr_14_port, QN => n177);
   PC_reg_15_inst : DFFR_X1 port map( D => n272, CK => Clk, RN => n311, Q => 
                           Iaddr_15_port, QN => n176);
   PC_reg_16_inst : DFFR_X1 port map( D => n271, CK => Clk, RN => n311, Q => 
                           Iaddr_16_port, QN => n175);
   PC_reg_17_inst : DFFR_X1 port map( D => n270, CK => Clk, RN => n311, Q => 
                           Iaddr_17_port, QN => n174);
   PC_reg_18_inst : DFFR_X1 port map( D => n269, CK => Clk, RN => n311, Q => 
                           Iaddr_18_port, QN => n173);
   PC_reg_19_inst : DFFR_X1 port map( D => n268, CK => Clk, RN => n311, Q => 
                           Iaddr_19_port, QN => n172);
   PC_reg_20_inst : DFFR_X1 port map( D => n267, CK => Clk, RN => n311, Q => 
                           Iaddr_20_port, QN => n171);
   PC_reg_21_inst : DFFR_X1 port map( D => n266, CK => Clk, RN => n312, Q => 
                           Iaddr_21_port, QN => n170);
   PC_reg_22_inst : DFFR_X1 port map( D => n265, CK => Clk, RN => n311, Q => 
                           Iaddr_22_port, QN => n169);
   PC_reg_23_inst : DFFR_X1 port map( D => n264, CK => Clk, RN => n312, Q => 
                           Iaddr_23_port, QN => n168);
   PC_reg_24_inst : DFFR_X1 port map( D => n263, CK => Clk, RN => n311, Q => 
                           Iaddr_24_port, QN => n167);
   PC_reg_25_inst : DFFR_X1 port map( D => n262, CK => Clk, RN => n312, Q => 
                           Iaddr_25_port, QN => n166);
   PC_reg_26_inst : DFFR_X1 port map( D => n261, CK => Clk, RN => n311, Q => 
                           Iaddr_26_port, QN => n165);
   PC_reg_27_inst : DFFR_X1 port map( D => n260, CK => Clk, RN => n312, Q => 
                           Iaddr_27_port, QN => n164);
   PC_reg_28_inst : DFFR_X1 port map( D => n259, CK => Clk, RN => n313, Q => 
                           Iaddr_28_port, QN => n163);
   PC_reg_29_inst : DFFR_X1 port map( D => n258, CK => Clk, RN => n312, Q => 
                           Iaddr_29_port, QN => n162);
   PC_reg_30_inst : DFFR_X1 port map( D => n257, CK => Clk, RN => n311, Q => 
                           Iaddr_30_port, QN => n161);
   NPC_reg_1_inst : DFFR_X1 port map( D => n256, CK => Clk, RN => n312, Q => 
                           NPC_1_port, QN => n160);
   NPC_reg_2_inst : DFFR_X1 port map( D => n255, CK => Clk, RN => n312, Q => 
                           NPC_2_port, QN => n159);
   NPC_reg_3_inst : DFFR_X1 port map( D => n254, CK => Clk, RN => n312, Q => 
                           NPC_3_port, QN => n158);
   NPC_reg_4_inst : DFFR_X1 port map( D => n253, CK => Clk, RN => n313, Q => 
                           NPC_4_port, QN => n157);
   NPC_reg_5_inst : DFFR_X1 port map( D => n252, CK => Clk, RN => n313, Q => 
                           NPC_5_port, QN => n156);
   NPC_reg_6_inst : DFFR_X1 port map( D => n251, CK => Clk, RN => n313, Q => 
                           NPC_6_port, QN => n155);
   NPC_reg_7_inst : DFFR_X1 port map( D => n250, CK => Clk, RN => n313, Q => 
                           NPC_7_port, QN => n154);
   NPC_reg_8_inst : DFFR_X1 port map( D => n249, CK => Clk, RN => n313, Q => 
                           NPC_8_port, QN => n153);
   NPC_reg_9_inst : DFFR_X1 port map( D => n248, CK => Clk, RN => n313, Q => 
                           NPC_9_port, QN => n152);
   NPC_reg_10_inst : DFFR_X1 port map( D => n247, CK => Clk, RN => n311, Q => 
                           NPC_10_port, QN => n151);
   NPC_reg_11_inst : DFFR_X1 port map( D => n246, CK => Clk, RN => n311, Q => 
                           NPC_11_port, QN => n150);
   NPC_reg_12_inst : DFFR_X1 port map( D => n245, CK => Clk, RN => n311, Q => 
                           NPC_12_port, QN => n149);
   NPC_reg_13_inst : DFFR_X1 port map( D => n244, CK => Clk, RN => n311, Q => 
                           NPC_13_port, QN => n148);
   NPC_reg_14_inst : DFFR_X1 port map( D => n243, CK => Clk, RN => n311, Q => 
                           NPC_14_port, QN => n147);
   NPC_reg_15_inst : DFFR_X1 port map( D => n242, CK => Clk, RN => n311, Q => 
                           NPC_15_port, QN => n146);
   NPC_reg_16_inst : DFFR_X1 port map( D => n241, CK => Clk, RN => n311, Q => 
                           NPC_16_port, QN => n145);
   NPC_reg_17_inst : DFFR_X1 port map( D => n240, CK => Clk, RN => n311, Q => 
                           NPC_17_port, QN => n144);
   NPC_reg_18_inst : DFFR_X1 port map( D => n239, CK => Clk, RN => n311, Q => 
                           NPC_18_port, QN => n143);
   NPC_reg_19_inst : DFFR_X1 port map( D => n238, CK => Clk, RN => n311, Q => 
                           NPC_19_port, QN => n142);
   NPC_reg_20_inst : DFFR_X1 port map( D => n237, CK => Clk, RN => n311, Q => 
                           NPC_20_port, QN => n141);
   NPC_reg_21_inst : DFFR_X1 port map( D => n236, CK => Clk, RN => n312, Q => 
                           NPC_21_port, QN => n140);
   NPC_reg_22_inst : DFFR_X1 port map( D => n235, CK => Clk, RN => n311, Q => 
                           NPC_22_port, QN => n139);
   NPC_reg_23_inst : DFFR_X1 port map( D => n234, CK => Clk, RN => n312, Q => 
                           NPC_23_port, QN => n138);
   NPC_reg_24_inst : DFFR_X1 port map( D => n233, CK => Clk, RN => n311, Q => 
                           NPC_24_port, QN => n137);
   NPC_reg_25_inst : DFFR_X1 port map( D => n232, CK => Clk, RN => n312, Q => 
                           NPC_25_port, QN => n136);
   NPC_reg_26_inst : DFFR_X1 port map( D => n231, CK => Clk, RN => n311, Q => 
                           NPC_26_port, QN => n135);
   NPC_reg_27_inst : DFFR_X1 port map( D => n230, CK => Clk, RN => n312, Q => 
                           NPC_27_port, QN => n134);
   NPC_reg_28_inst : DFFR_X1 port map( D => n229, CK => Clk, RN => n313, Q => 
                           NPC_28_port, QN => n133);
   NPC_reg_29_inst : DFFR_X1 port map( D => n228, CK => Clk, RN => n312, Q => 
                           NPC_29_port, QN => n132);
   NPC_reg_30_inst : DFFR_X1 port map( D => n227, CK => Clk, RN => n311, Q => 
                           NPC_30_port, QN => n131);
   NPC_reg_31_inst : DFFR_X1 port map( D => n226, CK => Clk, RN => n313, Q => 
                           NPC_31_port, QN => n130);
   IR_reg_0_inst : DFFR_X1 port map( D => n225, CK => Clk, RN => n312, Q => 
                           INP2_0_port, QN => n129);
   IR_reg_1_inst : DFFR_X1 port map( D => n224, CK => Clk, RN => n312, Q => 
                           INP2_1_port, QN => n128);
   IR_reg_2_inst : DFFR_X1 port map( D => n223, CK => Clk, RN => n312, Q => 
                           INP2_2_port, QN => n127);
   IR_reg_3_inst : DFFR_X1 port map( D => n222, CK => Clk, RN => n312, Q => 
                           INP2_3_port, QN => n126);
   IR_reg_4_inst : DFFR_X1 port map( D => n221, CK => Clk, RN => n312, Q => 
                           INP2_4_port, QN => n125);
   IR_reg_5_inst : DFFR_X1 port map( D => n220, CK => Clk, RN => n312, Q => 
                           INP2_5_port, QN => n124);
   IR_reg_6_inst : DFFR_X1 port map( D => n219, CK => Clk, RN => n312, Q => 
                           INP2_6_port, QN => n123);
   IR_reg_7_inst : DFFR_X1 port map( D => n218, CK => Clk, RN => n312, Q => 
                           INP2_7_port, QN => n122);
   IR_reg_8_inst : DFFR_X1 port map( D => n217, CK => Clk, RN => n312, Q => 
                           INP2_8_port, QN => n121);
   IR_reg_9_inst : DFFR_X1 port map( D => n216, CK => Clk, RN => n312, Q => 
                           INP2_9_port, QN => n120);
   IR_reg_10_inst : DFFR_X1 port map( D => n215, CK => Clk, RN => n312, Q => 
                           INP2_10_port, QN => n119);
   IR_reg_11_inst : DFFR_X1 port map( D => n214, CK => Clk, RN => n312, Q => 
                           INP2_11_port, QN => n118);
   IR_reg_12_inst : DFFR_X1 port map( D => n213, CK => Clk, RN => n312, Q => 
                           INP2_12_port, QN => n117);
   IR_reg_13_inst : DFFR_X1 port map( D => n212, CK => Clk, RN => n312, Q => 
                           INP2_13_port, QN => n116);
   IR_reg_14_inst : DFFR_X1 port map( D => n211, CK => Clk, RN => n312, Q => 
                           INP2_14_port, QN => n115);
   IR_reg_15_inst : DFFR_X1 port map( D => n210, CK => Clk, RN => n312, Q => 
                           INP2_15_port, QN => n114);
   IR_reg_16_inst : DFFR_X1 port map( D => n209, CK => Clk, RN => n312, Q => 
                           IMM26_16_port, QN => n113);
   IR_reg_17_inst : DFFR_X1 port map( D => n208, CK => Clk, RN => n312, Q => 
                           IMM26_17_port, QN => n112);
   IR_reg_18_inst : DFFR_X1 port map( D => n207, CK => Clk, RN => n312, Q => 
                           IMM26_18_port, QN => n111);
   IR_reg_19_inst : DFFR_X1 port map( D => n206, CK => Clk, RN => n312, Q => 
                           IMM26_19_port, QN => n110);
   IR_reg_20_inst : DFFR_X1 port map( D => n205, CK => Clk, RN => n312, Q => 
                           IMM26_20_port, QN => n109);
   IR_reg_21_inst : DFFR_X1 port map( D => n204, CK => Clk, RN => n312, Q => 
                           IMM26_21_port, QN => n108);
   IR_reg_22_inst : DFFR_X1 port map( D => n203, CK => Clk, RN => n312, Q => 
                           IMM26_22_port, QN => n107);
   IR_reg_23_inst : DFFR_X1 port map( D => n202, CK => Clk, RN => n312, Q => 
                           IMM26_23_port, QN => n106);
   IR_reg_24_inst : DFFR_X1 port map( D => n201, CK => Clk, RN => n312, Q => 
                           IMM26_24_port, QN => n105);
   IR_reg_25_inst : DFFR_X1 port map( D => n200, CK => Clk, RN => n312, Q => 
                           IMM26_25_port, QN => n104);
   IR_reg_26_inst : DFFR_X1 port map( D => n199, CK => Clk, RN => n312, Q => 
                           IR_26_port, QN => n103);
   IR_reg_27_inst : DFFR_X1 port map( D => n198, CK => Clk, RN => n312, Q => 
                           IR_27_port, QN => n102);
   IR_reg_28_inst : DFFR_X1 port map( D => n197, CK => Clk, RN => n312, Q => 
                           IR_28_port, QN => n101);
   IR_reg_29_inst : DFFR_X1 port map( D => n196, CK => Clk, RN => n312, Q => 
                           IR_29_port, QN => n100);
   IR_reg_30_inst : DFFR_X1 port map( D => n195, CK => Clk, RN => n313, Q => 
                           IR_30_port, QN => n99);
   IR_reg_31_inst : DFFR_X1 port map( D => n194, CK => Clk, RN => n313, Q => 
                           IR_31_port, QN => n98);
   U3 : OAI21_X1 port map( B1 => n304, B2 => n98, A => n2_port, ZN => n194);
   U4 : NAND2_X1 port map( A1 => Idata(31), A2 => n301, ZN => n2_port);
   U5 : OAI21_X1 port map( B1 => n304, B2 => n99, A => n3, ZN => n195);
   U6 : NAND2_X1 port map( A1 => Idata(30), A2 => n301, ZN => n3);
   U7 : OAI21_X1 port map( B1 => n303, B2 => n100, A => n4_port, ZN => n196);
   U8 : NAND2_X1 port map( A1 => Idata(29), A2 => n301, ZN => n4_port);
   U9 : OAI21_X1 port map( B1 => n303, B2 => n101, A => n5_port, ZN => n197);
   U10 : NAND2_X1 port map( A1 => Idata(28), A2 => n301, ZN => n5_port);
   U11 : OAI21_X1 port map( B1 => n303, B2 => n102, A => n6, ZN => n198);
   U12 : NAND2_X1 port map( A1 => Idata(27), A2 => n301, ZN => n6);
   U13 : OAI21_X1 port map( B1 => n302, B2 => n103, A => n7, ZN => n199);
   U14 : NAND2_X1 port map( A1 => Idata(26), A2 => n301, ZN => n7);
   U15 : OAI21_X1 port map( B1 => n303, B2 => n104, A => n8, ZN => n200);
   U16 : NAND2_X1 port map( A1 => Idata(25), A2 => n301, ZN => n8);
   U17 : OAI21_X1 port map( B1 => n302, B2 => n105, A => n9, ZN => n201);
   U18 : NAND2_X1 port map( A1 => Idata(24), A2 => n300, ZN => n9);
   U19 : OAI21_X1 port map( B1 => n302, B2 => n106, A => n10, ZN => n202);
   U20 : NAND2_X1 port map( A1 => Idata(23), A2 => n301, ZN => n10);
   U21 : OAI21_X1 port map( B1 => n302, B2 => n107, A => n11, ZN => n203);
   U22 : NAND2_X1 port map( A1 => Idata(22), A2 => n300, ZN => n11);
   U23 : OAI21_X1 port map( B1 => n301, B2 => n108, A => n12, ZN => n204);
   U24 : NAND2_X1 port map( A1 => Idata(21), A2 => n300, ZN => n12);
   U25 : OAI21_X1 port map( B1 => n301, B2 => n109, A => n13, ZN => n205);
   U26 : NAND2_X1 port map( A1 => Idata(20), A2 => n300, ZN => n13);
   U27 : OAI21_X1 port map( B1 => n302, B2 => n110, A => n14, ZN => n206);
   U28 : NAND2_X1 port map( A1 => Idata(19), A2 => n300, ZN => n14);
   U29 : OAI21_X1 port map( B1 => n301, B2 => n111, A => n15, ZN => n207);
   U30 : NAND2_X1 port map( A1 => Idata(18), A2 => n300, ZN => n15);
   U31 : OAI21_X1 port map( B1 => n301, B2 => n112, A => n16, ZN => n208);
   U32 : NAND2_X1 port map( A1 => Idata(17), A2 => n300, ZN => n16);
   U33 : OAI21_X1 port map( B1 => n302, B2 => n113, A => n17, ZN => n209);
   U34 : NAND2_X1 port map( A1 => Idata(16), A2 => n300, ZN => n17);
   U35 : OAI21_X1 port map( B1 => n302, B2 => n114, A => n18, ZN => n210);
   U36 : NAND2_X1 port map( A1 => Idata(15), A2 => n300, ZN => n18);
   U37 : OAI21_X1 port map( B1 => n302, B2 => n115, A => n19, ZN => n211);
   U38 : NAND2_X1 port map( A1 => Idata(14), A2 => n300, ZN => n19);
   U39 : OAI21_X1 port map( B1 => n302, B2 => n116, A => n20, ZN => n212);
   U40 : NAND2_X1 port map( A1 => Idata(13), A2 => n300, ZN => n20);
   U41 : OAI21_X1 port map( B1 => n302, B2 => n117, A => n21, ZN => n213);
   U42 : NAND2_X1 port map( A1 => Idata(12), A2 => n299, ZN => n21);
   U43 : OAI21_X1 port map( B1 => n302, B2 => n118, A => n22, ZN => n214);
   U44 : NAND2_X1 port map( A1 => Idata(11), A2 => n299, ZN => n22);
   U45 : OAI21_X1 port map( B1 => n303, B2 => n119, A => n23, ZN => n215);
   U46 : NAND2_X1 port map( A1 => Idata(10), A2 => n299, ZN => n23);
   U47 : OAI21_X1 port map( B1 => n302, B2 => n120, A => n24, ZN => n216);
   U48 : NAND2_X1 port map( A1 => Idata(9), A2 => n299, ZN => n24);
   U49 : OAI21_X1 port map( B1 => n303, B2 => n121, A => n25, ZN => n217);
   U50 : NAND2_X1 port map( A1 => Idata(8), A2 => n299, ZN => n25);
   U51 : OAI21_X1 port map( B1 => n303, B2 => n122, A => n26, ZN => n218);
   U52 : NAND2_X1 port map( A1 => Idata(7), A2 => n299, ZN => n26);
   U53 : OAI21_X1 port map( B1 => n303, B2 => n123, A => n27, ZN => n219);
   U54 : NAND2_X1 port map( A1 => Idata(6), A2 => n299, ZN => n27);
   U55 : OAI21_X1 port map( B1 => n303, B2 => n124, A => n28, ZN => n220);
   U56 : NAND2_X1 port map( A1 => Idata(5), A2 => n299, ZN => n28);
   U57 : OAI21_X1 port map( B1 => n303, B2 => n125, A => n29, ZN => n221);
   U58 : NAND2_X1 port map( A1 => Idata(4), A2 => n299, ZN => n29);
   U59 : OAI21_X1 port map( B1 => n303, B2 => n126, A => n30, ZN => n222);
   U60 : NAND2_X1 port map( A1 => Idata(3), A2 => n299, ZN => n30);
   U61 : OAI21_X1 port map( B1 => n303, B2 => n127, A => n31, ZN => n223);
   U62 : NAND2_X1 port map( A1 => Idata(2), A2 => n299, ZN => n31);
   U63 : OAI21_X1 port map( B1 => n304, B2 => n128, A => n32, ZN => n224);
   U64 : NAND2_X1 port map( A1 => Idata(1), A2 => n299, ZN => n32);
   U65 : OAI21_X1 port map( B1 => n304, B2 => n129, A => n33, ZN => n225);
   U66 : NAND2_X1 port map( A1 => Idata(0), A2 => n300, ZN => n33);
   U67 : OAI21_X1 port map( B1 => n310, B2 => n130, A => n34, ZN => n226);
   U68 : NAND2_X1 port map( A1 => n296, A2 => n307, ZN => n34);
   U69 : OAI21_X1 port map( B1 => n310, B2 => n131, A => n35, ZN => n227);
   U70 : NAND2_X1 port map( A1 => PC_next_30_port, A2 => n307, ZN => n35);
   U71 : OAI21_X1 port map( B1 => n309, B2 => n132, A => n36, ZN => n228);
   U72 : NAND2_X1 port map( A1 => PC_next_29_port, A2 => n307, ZN => n36);
   U73 : OAI21_X1 port map( B1 => n309, B2 => n133, A => n37, ZN => n229);
   U74 : NAND2_X1 port map( A1 => PC_next_28_port, A2 => n307, ZN => n37);
   U75 : OAI21_X1 port map( B1 => n309, B2 => n134, A => n38, ZN => n230);
   U76 : NAND2_X1 port map( A1 => PC_next_27_port, A2 => n307, ZN => n38);
   U77 : OAI21_X1 port map( B1 => n308, B2 => n135, A => n39, ZN => n231);
   U78 : NAND2_X1 port map( A1 => PC_next_26_port, A2 => n307, ZN => n39);
   U79 : OAI21_X1 port map( B1 => n309, B2 => n136, A => n40, ZN => n232);
   U80 : NAND2_X1 port map( A1 => PC_next_25_port, A2 => n307, ZN => n40);
   U81 : OAI21_X1 port map( B1 => n308, B2 => n137, A => n41, ZN => n233);
   U82 : NAND2_X1 port map( A1 => PC_next_24_port, A2 => n306, ZN => n41);
   U83 : OAI21_X1 port map( B1 => n308, B2 => n138, A => n42, ZN => n234);
   U84 : NAND2_X1 port map( A1 => PC_next_23_port, A2 => n307, ZN => n42);
   U85 : OAI21_X1 port map( B1 => n308, B2 => n139, A => n43, ZN => n235);
   U86 : NAND2_X1 port map( A1 => PC_next_22_port, A2 => n306, ZN => n43);
   U87 : OAI21_X1 port map( B1 => n307, B2 => n140, A => n44, ZN => n236);
   U88 : NAND2_X1 port map( A1 => PC_next_21_port, A2 => n306, ZN => n44);
   U89 : OAI21_X1 port map( B1 => n307, B2 => n141, A => n45, ZN => n237);
   U90 : NAND2_X1 port map( A1 => PC_next_20_port, A2 => n306, ZN => n45);
   U91 : OAI21_X1 port map( B1 => n308, B2 => n142, A => n46, ZN => n238);
   U92 : NAND2_X1 port map( A1 => PC_next_19_port, A2 => n306, ZN => n46);
   U93 : OAI21_X1 port map( B1 => n307, B2 => n143, A => n47, ZN => n239);
   U94 : NAND2_X1 port map( A1 => PC_next_18_port, A2 => n306, ZN => n47);
   U95 : OAI21_X1 port map( B1 => n307, B2 => n144, A => n48, ZN => n240);
   U96 : NAND2_X1 port map( A1 => PC_next_17_port, A2 => n306, ZN => n48);
   U97 : OAI21_X1 port map( B1 => n308, B2 => n145, A => n49, ZN => n241);
   U98 : NAND2_X1 port map( A1 => PC_next_16_port, A2 => n306, ZN => n49);
   U99 : OAI21_X1 port map( B1 => n308, B2 => n146, A => n50, ZN => n242);
   U100 : NAND2_X1 port map( A1 => PC_next_15_port, A2 => n306, ZN => n50);
   U101 : OAI21_X1 port map( B1 => n308, B2 => n147, A => n51, ZN => n243);
   U102 : NAND2_X1 port map( A1 => PC_next_14_port, A2 => n306, ZN => n51);
   U103 : OAI21_X1 port map( B1 => n308, B2 => n148, A => n52, ZN => n244);
   U104 : NAND2_X1 port map( A1 => PC_next_13_port, A2 => n306, ZN => n52);
   U105 : OAI21_X1 port map( B1 => n308, B2 => n149, A => n53, ZN => n245);
   U106 : NAND2_X1 port map( A1 => PC_next_12_port, A2 => n305, ZN => n53);
   U107 : OAI21_X1 port map( B1 => n308, B2 => n150, A => n54, ZN => n246);
   U108 : NAND2_X1 port map( A1 => PC_next_11_port, A2 => n305, ZN => n54);
   U109 : OAI21_X1 port map( B1 => n309, B2 => n151, A => n55, ZN => n247);
   U110 : NAND2_X1 port map( A1 => PC_next_10_port, A2 => n305, ZN => n55);
   U111 : OAI21_X1 port map( B1 => n308, B2 => n152, A => n56, ZN => n248);
   U112 : NAND2_X1 port map( A1 => PC_next_9_port, A2 => n305, ZN => n56);
   U113 : OAI21_X1 port map( B1 => n309, B2 => n153, A => n57, ZN => n249);
   U114 : NAND2_X1 port map( A1 => PC_next_8_port, A2 => n305, ZN => n57);
   U115 : OAI21_X1 port map( B1 => n309, B2 => n154, A => n58, ZN => n250);
   U116 : NAND2_X1 port map( A1 => PC_next_7_port, A2 => n305, ZN => n58);
   U117 : OAI21_X1 port map( B1 => n309, B2 => n155, A => n59, ZN => n251);
   U118 : NAND2_X1 port map( A1 => PC_next_6_port, A2 => n305, ZN => n59);
   U119 : OAI21_X1 port map( B1 => n309, B2 => n156, A => n60, ZN => n252);
   U120 : NAND2_X1 port map( A1 => PC_next_5_port, A2 => n305, ZN => n60);
   U121 : OAI21_X1 port map( B1 => n309, B2 => n157, A => n61, ZN => n253);
   U122 : NAND2_X1 port map( A1 => PC_next_4_port, A2 => n305, ZN => n61);
   U123 : OAI21_X1 port map( B1 => n309, B2 => n158, A => n62, ZN => n254);
   U124 : NAND2_X1 port map( A1 => PC_next_3_port, A2 => n305, ZN => n62);
   U125 : OAI21_X1 port map( B1 => n309, B2 => n159, A => n63, ZN => n255);
   U126 : NAND2_X1 port map( A1 => PC_next_2_port, A2 => n305, ZN => n63);
   U127 : OAI21_X1 port map( B1 => n310, B2 => n160, A => n64, ZN => n256);
   U128 : NAND2_X1 port map( A1 => PC_next_1_port, A2 => n305, ZN => n64);
   U129 : OAI21_X1 port map( B1 => PC_LATCH_EN_i, B2 => n161, A => n65, ZN => 
                           n257);
   U130 : NAND2_X1 port map( A1 => PC_LATCH_EN_i, A2 => PC_BUS_30_port, ZN => 
                           n65);
   U131 : OAI21_X1 port map( B1 => PC_LATCH_EN_i, B2 => n162, A => n66, ZN => 
                           n258);
   U132 : NAND2_X1 port map( A1 => PC_BUS_29_port, A2 => PC_LATCH_EN_i, ZN => 
                           n66);
   U133 : OAI21_X1 port map( B1 => PC_LATCH_EN_i, B2 => n163, A => n67, ZN => 
                           n259);
   U134 : NAND2_X1 port map( A1 => PC_BUS_28_port, A2 => PC_LATCH_EN_i, ZN => 
                           n67);
   U135 : OAI21_X1 port map( B1 => PC_LATCH_EN_i, B2 => n164, A => n68, ZN => 
                           n260);
   U136 : NAND2_X1 port map( A1 => PC_BUS_27_port, A2 => PC_LATCH_EN_i, ZN => 
                           n68);
   U137 : OAI21_X1 port map( B1 => PC_LATCH_EN_i, B2 => n165, A => n69, ZN => 
                           n261);
   U138 : NAND2_X1 port map( A1 => PC_BUS_26_port, A2 => PC_LATCH_EN_i, ZN => 
                           n69);
   U139 : OAI21_X1 port map( B1 => PC_LATCH_EN_i, B2 => n166, A => n70, ZN => 
                           n262);
   U140 : NAND2_X1 port map( A1 => PC_BUS_25_port, A2 => PC_LATCH_EN_i, ZN => 
                           n70);
   U141 : OAI21_X1 port map( B1 => PC_LATCH_EN_i, B2 => n167, A => n71, ZN => 
                           n263);
   U142 : NAND2_X1 port map( A1 => PC_BUS_24_port, A2 => PC_LATCH_EN_i, ZN => 
                           n71);
   U143 : OAI21_X1 port map( B1 => PC_LATCH_EN_i, B2 => n168, A => n72, ZN => 
                           n264);
   U144 : NAND2_X1 port map( A1 => PC_BUS_23_port, A2 => PC_LATCH_EN_i, ZN => 
                           n72);
   U145 : OAI21_X1 port map( B1 => PC_LATCH_EN_i, B2 => n169, A => n73, ZN => 
                           n265);
   U146 : NAND2_X1 port map( A1 => PC_BUS_22_port, A2 => PC_LATCH_EN_i, ZN => 
                           n73);
   U147 : OAI21_X1 port map( B1 => PC_LATCH_EN_i, B2 => n170, A => n74, ZN => 
                           n266);
   U148 : NAND2_X1 port map( A1 => PC_BUS_21_port, A2 => PC_LATCH_EN_i, ZN => 
                           n74);
   U149 : OAI21_X1 port map( B1 => PC_LATCH_EN_i, B2 => n171, A => n75, ZN => 
                           n267);
   U150 : NAND2_X1 port map( A1 => PC_BUS_20_port, A2 => PC_LATCH_EN_i, ZN => 
                           n75);
   U151 : OAI21_X1 port map( B1 => PC_LATCH_EN_i, B2 => n172, A => n76, ZN => 
                           n268);
   U152 : NAND2_X1 port map( A1 => PC_BUS_19_port, A2 => PC_LATCH_EN_i, ZN => 
                           n76);
   U153 : OAI21_X1 port map( B1 => PC_LATCH_EN_i, B2 => n173, A => n77, ZN => 
                           n269);
   U154 : NAND2_X1 port map( A1 => PC_BUS_18_port, A2 => PC_LATCH_EN_i, ZN => 
                           n77);
   U155 : OAI21_X1 port map( B1 => PC_LATCH_EN_i, B2 => n174, A => n78, ZN => 
                           n270);
   U156 : NAND2_X1 port map( A1 => PC_BUS_17_port, A2 => PC_LATCH_EN_i, ZN => 
                           n78);
   U157 : OAI21_X1 port map( B1 => PC_LATCH_EN_i, B2 => n175, A => n79, ZN => 
                           n271);
   U158 : NAND2_X1 port map( A1 => PC_BUS_16_port, A2 => PC_LATCH_EN_i, ZN => 
                           n79);
   U159 : OAI21_X1 port map( B1 => PC_LATCH_EN_i, B2 => n176, A => n80, ZN => 
                           n272);
   U160 : NAND2_X1 port map( A1 => PC_BUS_15_port, A2 => PC_LATCH_EN_i, ZN => 
                           n80);
   U161 : OAI21_X1 port map( B1 => PC_LATCH_EN_i, B2 => n177, A => n81, ZN => 
                           n273);
   U162 : NAND2_X1 port map( A1 => PC_BUS_14_port, A2 => PC_LATCH_EN_i, ZN => 
                           n81);
   U163 : OAI21_X1 port map( B1 => PC_LATCH_EN_i, B2 => n178, A => n82, ZN => 
                           n274);
   U164 : NAND2_X1 port map( A1 => PC_BUS_13_port, A2 => PC_LATCH_EN_i, ZN => 
                           n82);
   U165 : OAI21_X1 port map( B1 => PC_LATCH_EN_i, B2 => n179, A => n83, ZN => 
                           n275);
   U166 : NAND2_X1 port map( A1 => PC_BUS_12_port, A2 => PC_LATCH_EN_i, ZN => 
                           n83);
   U167 : OAI21_X1 port map( B1 => PC_LATCH_EN_i, B2 => n180, A => n84, ZN => 
                           n276);
   U168 : NAND2_X1 port map( A1 => PC_BUS_11_port, A2 => PC_LATCH_EN_i, ZN => 
                           n84);
   U169 : OAI21_X1 port map( B1 => PC_LATCH_EN_i, B2 => n181, A => n85, ZN => 
                           n277);
   U170 : NAND2_X1 port map( A1 => PC_BUS_10_port, A2 => PC_LATCH_EN_i, ZN => 
                           n85);
   U171 : OAI21_X1 port map( B1 => PC_LATCH_EN_i, B2 => n182, A => n86, ZN => 
                           n278);
   U172 : NAND2_X1 port map( A1 => PC_BUS_9_port, A2 => PC_LATCH_EN_i, ZN => 
                           n86);
   U173 : OAI21_X1 port map( B1 => PC_LATCH_EN_i, B2 => n183, A => n87, ZN => 
                           n279);
   U174 : NAND2_X1 port map( A1 => PC_BUS_8_port, A2 => PC_LATCH_EN_i, ZN => 
                           n87);
   U175 : OAI21_X1 port map( B1 => PC_LATCH_EN_i, B2 => n184, A => n88, ZN => 
                           n280);
   U176 : NAND2_X1 port map( A1 => PC_BUS_7_port, A2 => PC_LATCH_EN_i, ZN => 
                           n88);
   U177 : OAI21_X1 port map( B1 => PC_LATCH_EN_i, B2 => n185, A => n89, ZN => 
                           n281);
   U178 : NAND2_X1 port map( A1 => PC_BUS_6_port, A2 => PC_LATCH_EN_i, ZN => 
                           n89);
   U179 : OAI21_X1 port map( B1 => PC_LATCH_EN_i, B2 => n186, A => n90, ZN => 
                           n282);
   U180 : NAND2_X1 port map( A1 => PC_BUS_5_port, A2 => PC_LATCH_EN_i, ZN => 
                           n90);
   U181 : OAI21_X1 port map( B1 => PC_LATCH_EN_i, B2 => n187, A => n91, ZN => 
                           n283);
   U182 : NAND2_X1 port map( A1 => PC_BUS_4_port, A2 => PC_LATCH_EN_i, ZN => 
                           n91);
   U183 : OAI21_X1 port map( B1 => PC_LATCH_EN_i, B2 => n188, A => n92, ZN => 
                           n284);
   U184 : NAND2_X1 port map( A1 => PC_BUS_3_port, A2 => PC_LATCH_EN_i, ZN => 
                           n92);
   U185 : OAI21_X1 port map( B1 => PC_LATCH_EN_i, B2 => n189, A => n93, ZN => 
                           n285);
   U186 : NAND2_X1 port map( A1 => PC_BUS_2_port, A2 => PC_LATCH_EN_i, ZN => 
                           n93);
   U187 : OAI21_X1 port map( B1 => PC_LATCH_EN_i, B2 => n190, A => n94, ZN => 
                           n286);
   U188 : NAND2_X1 port map( A1 => PC_BUS_1_port, A2 => PC_LATCH_EN_i, ZN => 
                           n94);
   U189 : OAI21_X1 port map( B1 => PC_LATCH_EN_i, B2 => n191, A => n95, ZN => 
                           n287);
   U190 : NAND2_X1 port map( A1 => PC_BUS_0_port, A2 => PC_LATCH_EN_i, ZN => 
                           n95);
   U192 : NAND2_X1 port map( A1 => PC_BUS_31_port, A2 => PC_LATCH_EN_i, ZN => 
                           n96);
   U193 : OAI21_X1 port map( B1 => n310, B2 => n193, A => n97, ZN => n289);
   U194 : NAND2_X1 port map( A1 => PC_next_0_port, A2 => n306, ZN => n97);
   U195 : INV_X1 port map( A => n290, ZN => RD_4_port);
   U196 : AOI22_X1 port map( A1 => IMM26_20_port, A2 => n291, B1 => N2, B2 => 
                           INP2_15_port, ZN => n290);
   U197 : INV_X1 port map( A => n292, ZN => RD_3_port);
   U198 : AOI22_X1 port map( A1 => IMM26_19_port, A2 => n291, B1 => 
                           INP2_14_port, B2 => N2, ZN => n292);
   U199 : INV_X1 port map( A => n293, ZN => RD_2_port);
   U200 : AOI22_X1 port map( A1 => IMM26_18_port, A2 => n291, B1 => 
                           INP2_13_port, B2 => N2, ZN => n293);
   U201 : INV_X1 port map( A => n294, ZN => RD_1_port);
   U202 : AOI22_X1 port map( A1 => IMM26_17_port, A2 => n291, B1 => 
                           INP2_12_port, B2 => N2, ZN => n294);
   U203 : INV_X1 port map( A => n295, ZN => RD_0_port);
   U204 : AOI22_X1 port map( A1 => IMM26_16_port, A2 => n291, B1 => 
                           INP2_11_port, B2 => N2, ZN => n295);
   U205 : INV_X1 port map( A => N2, ZN => n291);
   NPC_logic_0 : NPC_logic_PC_SIZE32 port map( Flush_BTB => Flush_BTB, 
                           BRANCH_CTRL_SIG => BRANCH_CTRL_SIG, OUTT_NT_i => 
                           OUTT_NT_i, PC_next(31) => PC_next_31_port, 
                           PC_next(30) => PC_next_30_port, PC_next(29) => 
                           PC_next_29_port, PC_next(28) => PC_next_28_port, 
                           PC_next(27) => PC_next_27_port, PC_next(26) => 
                           PC_next_26_port, PC_next(25) => PC_next_25_port, 
                           PC_next(24) => PC_next_24_port, PC_next(23) => 
                           PC_next_23_port, PC_next(22) => PC_next_22_port, 
                           PC_next(21) => PC_next_21_port, PC_next(20) => 
                           PC_next_20_port, PC_next(19) => PC_next_19_port, 
                           PC_next(18) => PC_next_18_port, PC_next(17) => 
                           PC_next_17_port, PC_next(16) => PC_next_16_port, 
                           PC_next(15) => PC_next_15_port, PC_next(14) => 
                           PC_next_14_port, PC_next(13) => PC_next_13_port, 
                           PC_next(12) => PC_next_12_port, PC_next(11) => 
                           PC_next_11_port, PC_next(10) => PC_next_10_port, 
                           PC_next(9) => PC_next_9_port, PC_next(8) => 
                           PC_next_8_port, PC_next(7) => PC_next_7_port, 
                           PC_next(6) => PC_next_6_port, PC_next(5) => 
                           PC_next_5_port, PC_next(4) => PC_next_4_port, 
                           PC_next(3) => PC_next_3_port, PC_next(2) => 
                           PC_next_2_port, PC_next(1) => PC_next_1_port, 
                           PC_next(0) => PC_next_0_port, BRANCH_ALU_OUT(31) => 
                           BRANCH_ALU_OUT_31_port, BRANCH_ALU_OUT(30) => 
                           BRANCH_ALU_OUT_30_port, BRANCH_ALU_OUT(29) => 
                           BRANCH_ALU_OUT_29_port, BRANCH_ALU_OUT(28) => 
                           BRANCH_ALU_OUT_28_port, BRANCH_ALU_OUT(27) => 
                           BRANCH_ALU_OUT_27_port, BRANCH_ALU_OUT(26) => 
                           BRANCH_ALU_OUT_26_port, BRANCH_ALU_OUT(25) => 
                           BRANCH_ALU_OUT_25_port, BRANCH_ALU_OUT(24) => 
                           BRANCH_ALU_OUT_24_port, BRANCH_ALU_OUT(23) => 
                           BRANCH_ALU_OUT_23_port, BRANCH_ALU_OUT(22) => 
                           BRANCH_ALU_OUT_22_port, BRANCH_ALU_OUT(21) => 
                           BRANCH_ALU_OUT_21_port, BRANCH_ALU_OUT(20) => 
                           BRANCH_ALU_OUT_20_port, BRANCH_ALU_OUT(19) => 
                           BRANCH_ALU_OUT_19_port, BRANCH_ALU_OUT(18) => 
                           BRANCH_ALU_OUT_18_port, BRANCH_ALU_OUT(17) => 
                           BRANCH_ALU_OUT_17_port, BRANCH_ALU_OUT(16) => 
                           BRANCH_ALU_OUT_16_port, BRANCH_ALU_OUT(15) => 
                           BRANCH_ALU_OUT_15_port, BRANCH_ALU_OUT(14) => 
                           BRANCH_ALU_OUT_14_port, BRANCH_ALU_OUT(13) => 
                           BRANCH_ALU_OUT_13_port, BRANCH_ALU_OUT(12) => 
                           BRANCH_ALU_OUT_12_port, BRANCH_ALU_OUT(11) => 
                           BRANCH_ALU_OUT_11_port, BRANCH_ALU_OUT(10) => 
                           BRANCH_ALU_OUT_10_port, BRANCH_ALU_OUT(9) => 
                           BRANCH_ALU_OUT_9_port, BRANCH_ALU_OUT(8) => 
                           BRANCH_ALU_OUT_8_port, BRANCH_ALU_OUT(7) => 
                           BRANCH_ALU_OUT_7_port, BRANCH_ALU_OUT(6) => 
                           BRANCH_ALU_OUT_6_port, BRANCH_ALU_OUT(5) => 
                           BRANCH_ALU_OUT_5_port, BRANCH_ALU_OUT(4) => 
                           BRANCH_ALU_OUT_4_port, BRANCH_ALU_OUT(3) => 
                           BRANCH_ALU_OUT_3_port, BRANCH_ALU_OUT(2) => 
                           BRANCH_ALU_OUT_2_port, BRANCH_ALU_OUT(1) => 
                           BRANCH_ALU_OUT_1_port, BRANCH_ALU_OUT(0) => 
                           BRANCH_ALU_OUT_0_port, OUT_PC_target_i(31) => 
                           OUT_PC_target_i_31_port, OUT_PC_target_i(30) => 
                           OUT_PC_target_i_30_port, OUT_PC_target_i(29) => 
                           OUT_PC_target_i_29_port, OUT_PC_target_i(28) => 
                           OUT_PC_target_i_28_port, OUT_PC_target_i(27) => 
                           OUT_PC_target_i_27_port, OUT_PC_target_i(26) => 
                           OUT_PC_target_i_26_port, OUT_PC_target_i(25) => 
                           OUT_PC_target_i_25_port, OUT_PC_target_i(24) => 
                           OUT_PC_target_i_24_port, OUT_PC_target_i(23) => 
                           OUT_PC_target_i_23_port, OUT_PC_target_i(22) => 
                           OUT_PC_target_i_22_port, OUT_PC_target_i(21) => 
                           OUT_PC_target_i_21_port, OUT_PC_target_i(20) => 
                           OUT_PC_target_i_20_port, OUT_PC_target_i(19) => 
                           OUT_PC_target_i_19_port, OUT_PC_target_i(18) => 
                           OUT_PC_target_i_18_port, OUT_PC_target_i(17) => 
                           OUT_PC_target_i_17_port, OUT_PC_target_i(16) => 
                           OUT_PC_target_i_16_port, OUT_PC_target_i(15) => 
                           OUT_PC_target_i_15_port, OUT_PC_target_i(14) => 
                           OUT_PC_target_i_14_port, OUT_PC_target_i(13) => 
                           OUT_PC_target_i_13_port, OUT_PC_target_i(12) => 
                           OUT_PC_target_i_12_port, OUT_PC_target_i(11) => 
                           OUT_PC_target_i_11_port, OUT_PC_target_i(10) => 
                           OUT_PC_target_i_10_port, OUT_PC_target_i(9) => 
                           OUT_PC_target_i_9_port, OUT_PC_target_i(8) => 
                           OUT_PC_target_i_8_port, OUT_PC_target_i(7) => 
                           OUT_PC_target_i_7_port, OUT_PC_target_i(6) => 
                           OUT_PC_target_i_6_port, OUT_PC_target_i(5) => 
                           OUT_PC_target_i_5_port, OUT_PC_target_i(4) => 
                           OUT_PC_target_i_4_port, OUT_PC_target_i(3) => 
                           OUT_PC_target_i_3_port, OUT_PC_target_i(2) => 
                           OUT_PC_target_i_2_port, OUT_PC_target_i(1) => 
                           OUT_PC_target_i_1_port, OUT_PC_target_i(0) => 
                           OUT_PC_target_i_0_port, NPC(31) => NPC_31_port, 
                           NPC(30) => NPC_30_port, NPC(29) => NPC_29_port, 
                           NPC(28) => NPC_28_port, NPC(27) => NPC_27_port, 
                           NPC(26) => NPC_26_port, NPC(25) => NPC_25_port, 
                           NPC(24) => NPC_24_port, NPC(23) => NPC_23_port, 
                           NPC(22) => NPC_22_port, NPC(21) => NPC_21_port, 
                           NPC(20) => NPC_20_port, NPC(19) => NPC_19_port, 
                           NPC(18) => NPC_18_port, NPC(17) => NPC_17_port, 
                           NPC(16) => NPC_16_port, NPC(15) => NPC_15_port, 
                           NPC(14) => NPC_14_port, NPC(13) => NPC_13_port, 
                           NPC(12) => NPC_12_port, NPC(11) => NPC_11_port, 
                           NPC(10) => NPC_10_port, NPC(9) => NPC_9_port, NPC(8)
                           => NPC_8_port, NPC(7) => NPC_7_port, NPC(6) => 
                           NPC_6_port, NPC(5) => NPC_5_port, NPC(4) => 
                           NPC_4_port, NPC(3) => NPC_3_port, NPC(2) => 
                           NPC_2_port, NPC(1) => NPC_1_port, NPC(0) => 
                           NPC_0_port, PC_BUS(31) => PC_BUS_31_port, PC_BUS(30)
                           => PC_BUS_30_port, PC_BUS(29) => PC_BUS_29_port, 
                           PC_BUS(28) => PC_BUS_28_port, PC_BUS(27) => 
                           PC_BUS_27_port, PC_BUS(26) => PC_BUS_26_port, 
                           PC_BUS(25) => PC_BUS_25_port, PC_BUS(24) => 
                           PC_BUS_24_port, PC_BUS(23) => PC_BUS_23_port, 
                           PC_BUS(22) => PC_BUS_22_port, PC_BUS(21) => 
                           PC_BUS_21_port, PC_BUS(20) => PC_BUS_20_port, 
                           PC_BUS(19) => PC_BUS_19_port, PC_BUS(18) => 
                           PC_BUS_18_port, PC_BUS(17) => PC_BUS_17_port, 
                           PC_BUS(16) => PC_BUS_16_port, PC_BUS(15) => 
                           PC_BUS_15_port, PC_BUS(14) => PC_BUS_14_port, 
                           PC_BUS(13) => PC_BUS_13_port, PC_BUS(12) => 
                           PC_BUS_12_port, PC_BUS(11) => PC_BUS_11_port, 
                           PC_BUS(10) => PC_BUS_10_port, PC_BUS(9) => 
                           PC_BUS_9_port, PC_BUS(8) => PC_BUS_8_port, PC_BUS(7)
                           => PC_BUS_7_port, PC_BUS(6) => PC_BUS_6_port, 
                           PC_BUS(5) => PC_BUS_5_port, PC_BUS(4) => 
                           PC_BUS_4_port, PC_BUS(3) => PC_BUS_3_port, PC_BUS(2)
                           => PC_BUS_2_port, PC_BUS(1) => PC_BUS_1_port, 
                           PC_BUS(0) => PC_BUS_0_port);
   CU_I : dlx_cu_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE29 port map( Clk =>
                           Clk, Rst => n311, Flush_BTB => Flush_BTB_i, STALL =>
                           STALL_i, IR_IN(31) => IR_31_port, IR_IN(30) => 
                           IR_30_port, IR_IN(29) => IR_29_port, IR_IN(28) => 
                           IR_28_port, IR_IN(27) => IR_27_port, IR_IN(26) => 
                           IR_26_port, IR_IN(25) => IMM26_25_port, IR_IN(24) =>
                           IMM26_24_port, IR_IN(23) => IMM26_23_port, IR_IN(22)
                           => IMM26_22_port, IR_IN(21) => IMM26_21_port, 
                           IR_IN(20) => IMM26_20_port, IR_IN(19) => 
                           IMM26_19_port, IR_IN(18) => IMM26_18_port, IR_IN(17)
                           => IMM26_17_port, IR_IN(16) => IMM26_16_port, 
                           IR_IN(15) => INP2_15_port, IR_IN(14) => INP2_14_port
                           , IR_IN(13) => INP2_13_port, IR_IN(12) => 
                           INP2_12_port, IR_IN(11) => INP2_11_port, IR_IN(10) 
                           => INP2_10_port, IR_IN(9) => INP2_9_port, IR_IN(8) 
                           => INP2_8_port, IR_IN(7) => INP2_7_port, IR_IN(6) =>
                           INP2_6_port, IR_IN(5) => INP2_5_port, IR_IN(4) => 
                           INP2_4_port, IR_IN(3) => INP2_3_port, IR_IN(2) => 
                           INP2_2_port, IR_IN(1) => INP2_1_port, IR_IN(0) => 
                           INP2_0_port, IR_LATCH_EN => IR_LATCH_EN_i, 
                           NPC_LATCH_EN => NPC_LATCH_EN_i, I_R_type => 
                           I_R_TYPE_i, REGF_LATCH_EN => RegRF_LATCH_EN_i, 
                           RegA_LATCH_EN => RegA_LATCH_EN_i, RegB_LATCH_EN => 
                           RegB_LATCH_EN_i, RegIMM_LATCH_EN => 
                           RegIMM_LATCH_EN_i, RegRD1_LATCH_EN => 
                           RegRD1_LATCH_EN_i, SIGN_UNSIGN => SIGN_UNSIGN_i, 
                           RFR1_EN => RFR1_EN_i, RFR2_EN => RFR2_EN_i, 
                           MUX_IMM_SEL => MUX_IMM_SEL_i, JUMP => JUMP_i, 
                           JUMP_EN => JUMP_EN_i, EQ_COND => EQ_COND_i, MUXA_SEL
                           => MUXA_SEL_i, MUXB_SEL => MUXB_SEL_i, ALU_OUTREG_EN
                           => ALU_OUTREG_EN_i, REGME_LATCH_EN => 
                           REGME_LATCH_EN_i, RegRD2_LATCH_EN => 
                           RegRD2_LATCH_EN_i, ALU_OPCODE(0) => 
                           ALU_OPCODE_i_4_port, ALU_OPCODE(1) => 
                           ALU_OPCODE_i_3_port, ALU_OPCODE(2) => 
                           ALU_OPCODE_i_2_port, ALU_OPCODE(3) => 
                           ALU_OPCODE_i_1_port, ALU_OPCODE(4) => 
                           ALU_OPCODE_i_0_port, DRAM_EN => Denable, DRAM_RE => 
                           Drd, DRAM_WE => Dwd, LMD_LATCH_EN => LMD_LATCH_EN_i,
                           RALUOUT2_LATCH_EN => RALUOUT2_LATCH_EN_i, 
                           RegRD3_LATCH_EN => RegRD3_LATCH_EN_i, PC_LATCH_EN =>
                           PC_LATCH_EN_i, RPCplus8_LATCH_EN => 
                           RPCplus8_LATCH_EN_i, WB_MUX_SEL => WB_MUX_SEL_i, 
                           RF_WE => RF_WE_i, ROUT_LATCH_EN => n_1117, JandL => 
                           JandL_i, REGWRITE_DX => REGWRITE_DX_i, REGWRITE_XM 
                           => REGWRITE_XM_i, REGWRITE_MW => REGWRITE_MW_i, 
                           MEMREAD_DX => MEMREAD_DX_i);
   DP_I : datapath_NUMBIT32_ADDRESS_WIDTH_RF5_ADDRESS_WIDTH_DM32 port map( CLK 
                           => Clk, RST => n311, INP1(31) => NPC_31_port, 
                           INP1(30) => NPC_30_port, INP1(29) => NPC_29_port, 
                           INP1(28) => NPC_28_port, INP1(27) => NPC_27_port, 
                           INP1(26) => NPC_26_port, INP1(25) => NPC_25_port, 
                           INP1(24) => NPC_24_port, INP1(23) => NPC_23_port, 
                           INP1(22) => NPC_22_port, INP1(21) => NPC_21_port, 
                           INP1(20) => NPC_20_port, INP1(19) => NPC_19_port, 
                           INP1(18) => NPC_18_port, INP1(17) => NPC_17_port, 
                           INP1(16) => NPC_16_port, INP1(15) => NPC_15_port, 
                           INP1(14) => NPC_14_port, INP1(13) => NPC_13_port, 
                           INP1(12) => NPC_12_port, INP1(11) => NPC_11_port, 
                           INP1(10) => NPC_10_port, INP1(9) => NPC_9_port, 
                           INP1(8) => NPC_8_port, INP1(7) => NPC_7_port, 
                           INP1(6) => NPC_6_port, INP1(5) => NPC_5_port, 
                           INP1(4) => NPC_4_port, INP1(3) => NPC_3_port, 
                           INP1(2) => NPC_2_port, INP1(1) => NPC_1_port, 
                           INP1(0) => NPC_0_port, INP2(15) => INP2_15_port, 
                           INP2(14) => INP2_14_port, INP2(13) => INP2_13_port, 
                           INP2(12) => INP2_12_port, INP2(11) => INP2_11_port, 
                           INP2(10) => INP2_10_port, INP2(9) => INP2_9_port, 
                           INP2(8) => INP2_8_port, INP2(7) => INP2_7_port, 
                           INP2(6) => INP2_6_port, INP2(5) => INP2_5_port, 
                           INP2(4) => INP2_4_port, INP2(3) => INP2_3_port, 
                           INP2(2) => INP2_2_port, INP2(1) => INP2_1_port, 
                           INP2(0) => INP2_0_port, IMM26(25) => IMM26_25_port, 
                           IMM26(24) => IMM26_24_port, IMM26(23) => 
                           IMM26_23_port, IMM26(22) => IMM26_22_port, IMM26(21)
                           => IMM26_21_port, IMM26(20) => IMM26_20_port, 
                           IMM26(19) => IMM26_19_port, IMM26(18) => 
                           IMM26_18_port, IMM26(17) => IMM26_17_port, IMM26(16)
                           => IMM26_16_port, IMM26(15) => INP2_15_port, 
                           IMM26(14) => INP2_14_port, IMM26(13) => INP2_13_port
                           , IMM26(12) => INP2_12_port, IMM26(11) => 
                           INP2_11_port, IMM26(10) => INP2_10_port, IMM26(9) =>
                           INP2_9_port, IMM26(8) => INP2_8_port, IMM26(7) => 
                           INP2_7_port, IMM26(6) => INP2_6_port, IMM26(5) => 
                           INP2_5_port, IMM26(4) => INP2_4_port, IMM26(3) => 
                           INP2_3_port, IMM26(2) => INP2_2_port, IMM26(1) => 
                           INP2_1_port, IMM26(0) => INP2_0_port, RS1(4) => 
                           IMM26_25_port, RS1(3) => IMM26_24_port, RS1(2) => 
                           IMM26_23_port, RS1(1) => IMM26_22_port, RS1(0) => 
                           IMM26_21_port, RS2(4) => IMM26_20_port, RS2(3) => 
                           IMM26_19_port, RS2(2) => IMM26_18_port, RS2(1) => 
                           IMM26_17_port, RS2(0) => IMM26_16_port, RD(4) => 
                           RD_4_port, RD(3) => RD_3_port, RD(2) => RD_2_port, 
                           RD(1) => RD_1_port, RD(0) => RD_0_port, 
                           REGF_LATCH_EN => RegRF_LATCH_EN_i, RegA_LATCH_EN => 
                           RegA_LATCH_EN_i, RegB_LATCH_EN => RegB_LATCH_EN_i, 
                           RegIMM_LATCH_EN => RegIMM_LATCH_EN_i, 
                           RegRD1_LATCH_EN => RegRD1_LATCH_EN_i, SIGN_UNSIGN =>
                           SIGN_UNSIGN_i, RFR1_EN => RFR1_EN_i, RFR2_EN => 
                           RFR2_EN_i, MUX_IMM_SEL => MUX_IMM_SEL_i, JUMP => 
                           JUMP_i, JUMP_EN => JUMP_EN_i, EQ_COND => EQ_COND_i, 
                           MUXA_SEL => MUXA_SEL_i, MUXB_SEL => MUXB_SEL_i, 
                           RALUOUT_LATCH_EN => ALU_OUTREG_EN_i, REGME_LATCH_EN 
                           => REGME_LATCH_EN_i, RegRD2_LATCH_EN => 
                           RegRD2_LATCH_EN_i, ALU_OPCODE(0) => 
                           ALU_OPCODE_i_4_port, ALU_OPCODE(1) => 
                           ALU_OPCODE_i_3_port, ALU_OPCODE(2) => 
                           ALU_OPCODE_i_2_port, ALU_OPCODE(3) => 
                           ALU_OPCODE_i_1_port, ALU_OPCODE(4) => 
                           ALU_OPCODE_i_0_port, ADDR_DRAM(31) => Daddr(31), 
                           ADDR_DRAM(30) => Daddr(30), ADDR_DRAM(29) => 
                           Daddr(29), ADDR_DRAM(28) => Daddr(28), ADDR_DRAM(27)
                           => Daddr(27), ADDR_DRAM(26) => Daddr(26), 
                           ADDR_DRAM(25) => Daddr(25), ADDR_DRAM(24) => 
                           Daddr(24), ADDR_DRAM(23) => Daddr(23), ADDR_DRAM(22)
                           => Daddr(22), ADDR_DRAM(21) => Daddr(21), 
                           ADDR_DRAM(20) => Daddr(20), ADDR_DRAM(19) => 
                           Daddr(19), ADDR_DRAM(18) => Daddr(18), ADDR_DRAM(17)
                           => Daddr(17), ADDR_DRAM(16) => Daddr(16), 
                           ADDR_DRAM(15) => Daddr(15), ADDR_DRAM(14) => 
                           Daddr(14), ADDR_DRAM(13) => Daddr(13), ADDR_DRAM(12)
                           => Daddr(12), ADDR_DRAM(11) => Daddr(11), 
                           ADDR_DRAM(10) => Daddr(10), ADDR_DRAM(9) => Daddr(9)
                           , ADDR_DRAM(8) => Daddr(8), ADDR_DRAM(7) => Daddr(7)
                           , ADDR_DRAM(6) => Daddr(6), ADDR_DRAM(5) => Daddr(5)
                           , ADDR_DRAM(4) => Daddr(4), ADDR_DRAM(3) => Daddr(3)
                           , ADDR_DRAM(2) => Daddr(2), ADDR_DRAM(1) => Daddr(1)
                           , ADDR_DRAM(0) => Daddr(0), DATAIN_DRAM(31) => 
                           Ddatain(31), DATAIN_DRAM(30) => Ddatain(30), 
                           DATAIN_DRAM(29) => Ddatain(29), DATAIN_DRAM(28) => 
                           Ddatain(28), DATAIN_DRAM(27) => Ddatain(27), 
                           DATAIN_DRAM(26) => Ddatain(26), DATAIN_DRAM(25) => 
                           Ddatain(25), DATAIN_DRAM(24) => Ddatain(24), 
                           DATAIN_DRAM(23) => Ddatain(23), DATAIN_DRAM(22) => 
                           Ddatain(22), DATAIN_DRAM(21) => Ddatain(21), 
                           DATAIN_DRAM(20) => Ddatain(20), DATAIN_DRAM(19) => 
                           Ddatain(19), DATAIN_DRAM(18) => Ddatain(18), 
                           DATAIN_DRAM(17) => Ddatain(17), DATAIN_DRAM(16) => 
                           Ddatain(16), DATAIN_DRAM(15) => Ddatain(15), 
                           DATAIN_DRAM(14) => Ddatain(14), DATAIN_DRAM(13) => 
                           Ddatain(13), DATAIN_DRAM(12) => Ddatain(12), 
                           DATAIN_DRAM(11) => Ddatain(11), DATAIN_DRAM(10) => 
                           Ddatain(10), DATAIN_DRAM(9) => Ddatain(9), 
                           DATAIN_DRAM(8) => Ddatain(8), DATAIN_DRAM(7) => 
                           Ddatain(7), DATAIN_DRAM(6) => Ddatain(6), 
                           DATAIN_DRAM(5) => Ddatain(5), DATAIN_DRAM(4) => 
                           Ddatain(4), DATAIN_DRAM(3) => Ddatain(3), 
                           DATAIN_DRAM(2) => Ddatain(2), DATAIN_DRAM(1) => 
                           Ddatain(1), DATAIN_DRAM(0) => Ddatain(0), 
                           DATAOUT_DRAM(31) => Ddataout(31), DATAOUT_DRAM(30) 
                           => Ddataout(30), DATAOUT_DRAM(29) => Ddataout(29), 
                           DATAOUT_DRAM(28) => Ddataout(28), DATAOUT_DRAM(27) 
                           => Ddataout(27), DATAOUT_DRAM(26) => Ddataout(26), 
                           DATAOUT_DRAM(25) => Ddataout(25), DATAOUT_DRAM(24) 
                           => Ddataout(24), DATAOUT_DRAM(23) => Ddataout(23), 
                           DATAOUT_DRAM(22) => Ddataout(22), DATAOUT_DRAM(21) 
                           => Ddataout(21), DATAOUT_DRAM(20) => Ddataout(20), 
                           DATAOUT_DRAM(19) => Ddataout(19), DATAOUT_DRAM(18) 
                           => Ddataout(18), DATAOUT_DRAM(17) => Ddataout(17), 
                           DATAOUT_DRAM(16) => Ddataout(16), DATAOUT_DRAM(15) 
                           => Ddataout(15), DATAOUT_DRAM(14) => Ddataout(14), 
                           DATAOUT_DRAM(13) => Ddataout(13), DATAOUT_DRAM(12) 
                           => Ddataout(12), DATAOUT_DRAM(11) => Ddataout(11), 
                           DATAOUT_DRAM(10) => Ddataout(10), DATAOUT_DRAM(9) =>
                           Ddataout(9), DATAOUT_DRAM(8) => Ddataout(8), 
                           DATAOUT_DRAM(7) => Ddataout(7), DATAOUT_DRAM(6) => 
                           Ddataout(6), DATAOUT_DRAM(5) => Ddataout(5), 
                           DATAOUT_DRAM(4) => Ddataout(4), DATAOUT_DRAM(3) => 
                           Ddataout(3), DATAOUT_DRAM(2) => Ddataout(2), 
                           DATAOUT_DRAM(1) => Ddataout(1), DATAOUT_DRAM(0) => 
                           Ddataout(0), LMD_LATCH_EN => LMD_LATCH_EN_i, 
                           RALUOUT2_LATCH_EN => RALUOUT2_LATCH_EN_i, 
                           RegRD3_LATCH_EN => RegRD3_LATCH_EN_i, 
                           RPCplus8_LATCH_EN => RPCplus8_LATCH_EN_i, WB_MUX_SEL
                           => WB_MUX_SEL_i, RF_WE => RF_WE_i, ROUT_LATCH_EN => 
                           ROUT_LATCH_EN_i, JandL => JandL_i, BRANCH_CTRL_SIG 
                           => BRANCH_CTRL_SIG, BRANCH_ALU_OUT(31) => 
                           BRANCH_ALU_OUT_31_port, BRANCH_ALU_OUT(30) => 
                           BRANCH_ALU_OUT_30_port, BRANCH_ALU_OUT(29) => 
                           BRANCH_ALU_OUT_29_port, BRANCH_ALU_OUT(28) => 
                           BRANCH_ALU_OUT_28_port, BRANCH_ALU_OUT(27) => 
                           BRANCH_ALU_OUT_27_port, BRANCH_ALU_OUT(26) => 
                           BRANCH_ALU_OUT_26_port, BRANCH_ALU_OUT(25) => 
                           BRANCH_ALU_OUT_25_port, BRANCH_ALU_OUT(24) => 
                           BRANCH_ALU_OUT_24_port, BRANCH_ALU_OUT(23) => 
                           BRANCH_ALU_OUT_23_port, BRANCH_ALU_OUT(22) => 
                           BRANCH_ALU_OUT_22_port, BRANCH_ALU_OUT(21) => 
                           BRANCH_ALU_OUT_21_port, BRANCH_ALU_OUT(20) => 
                           BRANCH_ALU_OUT_20_port, BRANCH_ALU_OUT(19) => 
                           BRANCH_ALU_OUT_19_port, BRANCH_ALU_OUT(18) => 
                           BRANCH_ALU_OUT_18_port, BRANCH_ALU_OUT(17) => 
                           BRANCH_ALU_OUT_17_port, BRANCH_ALU_OUT(16) => 
                           BRANCH_ALU_OUT_16_port, BRANCH_ALU_OUT(15) => 
                           BRANCH_ALU_OUT_15_port, BRANCH_ALU_OUT(14) => 
                           BRANCH_ALU_OUT_14_port, BRANCH_ALU_OUT(13) => 
                           BRANCH_ALU_OUT_13_port, BRANCH_ALU_OUT(12) => 
                           BRANCH_ALU_OUT_12_port, BRANCH_ALU_OUT(11) => 
                           BRANCH_ALU_OUT_11_port, BRANCH_ALU_OUT(10) => 
                           BRANCH_ALU_OUT_10_port, BRANCH_ALU_OUT(9) => 
                           BRANCH_ALU_OUT_9_port, BRANCH_ALU_OUT(8) => 
                           BRANCH_ALU_OUT_8_port, BRANCH_ALU_OUT(7) => 
                           BRANCH_ALU_OUT_7_port, BRANCH_ALU_OUT(6) => 
                           BRANCH_ALU_OUT_6_port, BRANCH_ALU_OUT(5) => 
                           BRANCH_ALU_OUT_5_port, BRANCH_ALU_OUT(4) => 
                           BRANCH_ALU_OUT_4_port, BRANCH_ALU_OUT(3) => 
                           BRANCH_ALU_OUT_3_port, BRANCH_ALU_OUT(2) => 
                           BRANCH_ALU_OUT_2_port, BRANCH_ALU_OUT(1) => 
                           BRANCH_ALU_OUT_1_port, BRANCH_ALU_OUT(0) => 
                           BRANCH_ALU_OUT_0_port, Data_out(31) => DataOut(31), 
                           Data_out(30) => DataOut(30), Data_out(29) => 
                           DataOut(29), Data_out(28) => DataOut(28), 
                           Data_out(27) => DataOut(27), Data_out(26) => 
                           DataOut(26), Data_out(25) => DataOut(25), 
                           Data_out(24) => DataOut(24), Data_out(23) => 
                           DataOut(23), Data_out(22) => DataOut(22), 
                           Data_out(21) => DataOut(21), Data_out(20) => 
                           DataOut(20), Data_out(19) => DataOut(19), 
                           Data_out(18) => DataOut(18), Data_out(17) => 
                           DataOut(17), Data_out(16) => DataOut(16), 
                           Data_out(15) => DataOut(15), Data_out(14) => 
                           DataOut(14), Data_out(13) => DataOut(13), 
                           Data_out(12) => DataOut(12), Data_out(11) => 
                           DataOut(11), Data_out(10) => DataOut(10), 
                           Data_out(9) => DataOut(9), Data_out(8) => DataOut(8)
                           , Data_out(7) => DataOut(7), Data_out(6) => 
                           DataOut(6), Data_out(5) => DataOut(5), Data_out(4) 
                           => DataOut(4), Data_out(3) => DataOut(3), 
                           Data_out(2) => DataOut(2), Data_out(1) => DataOut(1)
                           , Data_out(0) => DataOut(0), REGWRITE_XM => 
                           REGWRITE_XM_i, REGWRITE_MW => REGWRITE_MW_i);
   BTB_0 : BTB_PC_SIZE32_BTBSIZE5 port map( Reset => n311, Clk => Clk, Enable 
                           => X_Logic1_port, PC_read(31) => n296, PC_read(30) 
                           => PC_next_30_port, PC_read(29) => PC_next_29_port, 
                           PC_read(28) => PC_next_28_port, PC_read(27) => 
                           PC_next_27_port, PC_read(26) => PC_next_26_port, 
                           PC_read(25) => PC_next_25_port, PC_read(24) => 
                           PC_next_24_port, PC_read(23) => PC_next_23_port, 
                           PC_read(22) => PC_next_22_port, PC_read(21) => 
                           PC_next_21_port, PC_read(20) => PC_next_20_port, 
                           PC_read(19) => PC_next_19_port, PC_read(18) => 
                           PC_next_18_port, PC_read(17) => PC_next_17_port, 
                           PC_read(16) => PC_next_16_port, PC_read(15) => 
                           PC_next_15_port, PC_read(14) => PC_next_14_port, 
                           PC_read(13) => PC_next_13_port, PC_read(12) => 
                           PC_next_12_port, PC_read(11) => PC_next_11_port, 
                           PC_read(10) => PC_next_10_port, PC_read(9) => 
                           PC_next_9_port, PC_read(8) => PC_next_8_port, 
                           PC_read(7) => PC_next_7_port, PC_read(6) => 
                           PC_next_6_port, PC_read(5) => PC_next_5_port, 
                           PC_read(4) => PC_next_4_port, PC_read(3) => 
                           PC_next_3_port, PC_read(2) => PC_next_2_port, 
                           PC_read(1) => PC_next_1_port, PC_read(0) => 
                           PC_next_0_port, WR => JUMP_EN_i, PC_write(31) => 
                           NPC_31_port, PC_write(30) => NPC_30_port, 
                           PC_write(29) => NPC_29_port, PC_write(28) => 
                           NPC_28_port, PC_write(27) => NPC_27_port, 
                           PC_write(26) => NPC_26_port, PC_write(25) => 
                           NPC_25_port, PC_write(24) => NPC_24_port, 
                           PC_write(23) => NPC_23_port, PC_write(22) => 
                           NPC_22_port, PC_write(21) => NPC_21_port, 
                           PC_write(20) => NPC_20_port, PC_write(19) => 
                           NPC_19_port, PC_write(18) => NPC_18_port, 
                           PC_write(17) => NPC_17_port, PC_write(16) => 
                           NPC_16_port, PC_write(15) => NPC_15_port, 
                           PC_write(14) => NPC_14_port, PC_write(13) => 
                           NPC_13_port, PC_write(12) => NPC_12_port, 
                           PC_write(11) => NPC_11_port, PC_write(10) => 
                           NPC_10_port, PC_write(9) => NPC_9_port, PC_write(8) 
                           => NPC_8_port, PC_write(7) => NPC_7_port, 
                           PC_write(6) => NPC_6_port, PC_write(5) => NPC_5_port
                           , PC_write(4) => NPC_4_port, PC_write(3) => 
                           NPC_3_port, PC_write(2) => NPC_2_port, PC_write(1) 
                           => NPC_1_port, PC_write(0) => NPC_0_port, SetT_NT =>
                           BRANCH_CTRL_SIG, Set_target(31) => 
                           BRANCH_ALU_OUT_31_port, Set_target(30) => 
                           BRANCH_ALU_OUT_30_port, Set_target(29) => 
                           BRANCH_ALU_OUT_29_port, Set_target(28) => 
                           BRANCH_ALU_OUT_28_port, Set_target(27) => 
                           BRANCH_ALU_OUT_27_port, Set_target(26) => 
                           BRANCH_ALU_OUT_26_port, Set_target(25) => 
                           BRANCH_ALU_OUT_25_port, Set_target(24) => 
                           BRANCH_ALU_OUT_24_port, Set_target(23) => 
                           BRANCH_ALU_OUT_23_port, Set_target(22) => 
                           BRANCH_ALU_OUT_22_port, Set_target(21) => 
                           BRANCH_ALU_OUT_21_port, Set_target(20) => 
                           BRANCH_ALU_OUT_20_port, Set_target(19) => 
                           BRANCH_ALU_OUT_19_port, Set_target(18) => 
                           BRANCH_ALU_OUT_18_port, Set_target(17) => 
                           BRANCH_ALU_OUT_17_port, Set_target(16) => 
                           BRANCH_ALU_OUT_16_port, Set_target(15) => 
                           BRANCH_ALU_OUT_15_port, Set_target(14) => 
                           BRANCH_ALU_OUT_14_port, Set_target(13) => 
                           BRANCH_ALU_OUT_13_port, Set_target(12) => 
                           BRANCH_ALU_OUT_12_port, Set_target(11) => 
                           BRANCH_ALU_OUT_11_port, Set_target(10) => 
                           BRANCH_ALU_OUT_10_port, Set_target(9) => 
                           BRANCH_ALU_OUT_9_port, Set_target(8) => 
                           BRANCH_ALU_OUT_8_port, Set_target(7) => 
                           BRANCH_ALU_OUT_7_port, Set_target(6) => 
                           BRANCH_ALU_OUT_6_port, Set_target(5) => 
                           BRANCH_ALU_OUT_5_port, Set_target(4) => 
                           BRANCH_ALU_OUT_4_port, Set_target(3) => 
                           BRANCH_ALU_OUT_3_port, Set_target(2) => 
                           BRANCH_ALU_OUT_2_port, Set_target(1) => 
                           BRANCH_ALU_OUT_1_port, Set_target(0) => 
                           BRANCH_ALU_OUT_0_port, OUT_PC_target(31) => 
                           OUT_PC_target_i_31_port, OUT_PC_target(30) => 
                           OUT_PC_target_i_30_port, OUT_PC_target(29) => 
                           OUT_PC_target_i_29_port, OUT_PC_target(28) => 
                           OUT_PC_target_i_28_port, OUT_PC_target(27) => 
                           OUT_PC_target_i_27_port, OUT_PC_target(26) => 
                           OUT_PC_target_i_26_port, OUT_PC_target(25) => 
                           OUT_PC_target_i_25_port, OUT_PC_target(24) => 
                           OUT_PC_target_i_24_port, OUT_PC_target(23) => 
                           OUT_PC_target_i_23_port, OUT_PC_target(22) => 
                           OUT_PC_target_i_22_port, OUT_PC_target(21) => 
                           OUT_PC_target_i_21_port, OUT_PC_target(20) => 
                           OUT_PC_target_i_20_port, OUT_PC_target(19) => 
                           OUT_PC_target_i_19_port, OUT_PC_target(18) => 
                           OUT_PC_target_i_18_port, OUT_PC_target(17) => 
                           OUT_PC_target_i_17_port, OUT_PC_target(16) => 
                           OUT_PC_target_i_16_port, OUT_PC_target(15) => 
                           OUT_PC_target_i_15_port, OUT_PC_target(14) => 
                           OUT_PC_target_i_14_port, OUT_PC_target(13) => 
                           OUT_PC_target_i_13_port, OUT_PC_target(12) => 
                           OUT_PC_target_i_12_port, OUT_PC_target(11) => 
                           OUT_PC_target_i_11_port, OUT_PC_target(10) => 
                           OUT_PC_target_i_10_port, OUT_PC_target(9) => 
                           OUT_PC_target_i_9_port, OUT_PC_target(8) => 
                           OUT_PC_target_i_8_port, OUT_PC_target(7) => 
                           OUT_PC_target_i_7_port, OUT_PC_target(6) => 
                           OUT_PC_target_i_6_port, OUT_PC_target(5) => 
                           OUT_PC_target_i_5_port, OUT_PC_target(4) => 
                           OUT_PC_target_i_4_port, OUT_PC_target(3) => 
                           OUT_PC_target_i_3_port, OUT_PC_target(2) => 
                           OUT_PC_target_i_2_port, OUT_PC_target(1) => 
                           OUT_PC_target_i_1_port, OUT_PC_target(0) => 
                           OUT_PC_target_i_0_port, OUTT_NT => OUTT_NT_i, 
                           prevT_NT => prevT_NT_i);
   HU_0 : HazardUnit_NUMBIT32_ADDRESS_WIDTH_RF5_OP_CODE_SIZE6 port map( CLK => 
                           Clk, RST => n311, RS1(4) => IMM26_25_port, RS1(3) =>
                           IMM26_24_port, RS1(2) => IMM26_23_port, RS1(1) => 
                           IMM26_22_port, RS1(0) => IMM26_21_port, RS2(4) => 
                           IMM26_20_port, RS2(3) => IMM26_19_port, RS2(2) => 
                           IMM26_18_port, RS2(1) => IMM26_17_port, RS2(0) => 
                           IMM26_16_port, REGWRITE_DX => REGWRITE_DX_i, 
                           MEMREAD_DX => MEMREAD_DX_i, RD(4) => IMM26_20_port, 
                           RD(3) => IMM26_19_port, RD(2) => IMM26_18_port, 
                           RD(1) => IMM26_17_port, RD(0) => IMM26_16_port, 
                           OPCODE(5) => IR_31_port, OPCODE(4) => IR_30_port, 
                           OPCODE(3) => IR_29_port, OPCODE(2) => IR_28_port, 
                           OPCODE(1) => IR_27_port, OPCODE(0) => IR_26_port, 
                           STALL => STALL_i);
   add_365 : DLX_IR_SIZE32_PC_SIZE32_DW01_inc_1 port map( A(31) => 
                           Iaddr_31_port, A(30) => Iaddr_30_port, A(29) => 
                           Iaddr_29_port, A(28) => Iaddr_28_port, A(27) => 
                           Iaddr_27_port, A(26) => Iaddr_26_port, A(25) => 
                           Iaddr_25_port, A(24) => Iaddr_24_port, A(23) => 
                           Iaddr_23_port, A(22) => Iaddr_22_port, A(21) => 
                           Iaddr_21_port, A(20) => Iaddr_20_port, A(19) => 
                           Iaddr_19_port, A(18) => Iaddr_18_port, A(17) => 
                           Iaddr_17_port, A(16) => Iaddr_16_port, A(15) => 
                           Iaddr_15_port, A(14) => Iaddr_14_port, A(13) => 
                           Iaddr_13_port, A(12) => Iaddr_12_port, A(11) => 
                           Iaddr_11_port, A(10) => Iaddr_10_port, A(9) => 
                           Iaddr_9_port, A(8) => Iaddr_8_port, A(7) => 
                           Iaddr_7_port, A(6) => Iaddr_6_port, A(5) => 
                           Iaddr_5_port, A(4) => Iaddr_4_port, A(3) => 
                           Iaddr_3_port, A(2) => Iaddr_2_port, A(1) => 
                           Iaddr_1_port, A(0) => n314, SUM(31) => 
                           PC_next_31_port, SUM(30) => PC_next_30_port, SUM(29)
                           => PC_next_29_port, SUM(28) => PC_next_28_port, 
                           SUM(27) => PC_next_27_port, SUM(26) => 
                           PC_next_26_port, SUM(25) => PC_next_25_port, SUM(24)
                           => PC_next_24_port, SUM(23) => PC_next_23_port, 
                           SUM(22) => PC_next_22_port, SUM(21) => 
                           PC_next_21_port, SUM(20) => PC_next_20_port, SUM(19)
                           => PC_next_19_port, SUM(18) => PC_next_18_port, 
                           SUM(17) => PC_next_17_port, SUM(16) => 
                           PC_next_16_port, SUM(15) => PC_next_15_port, SUM(14)
                           => PC_next_14_port, SUM(13) => PC_next_13_port, 
                           SUM(12) => PC_next_12_port, SUM(11) => 
                           PC_next_11_port, SUM(10) => PC_next_10_port, SUM(9) 
                           => PC_next_9_port, SUM(8) => PC_next_8_port, SUM(7) 
                           => PC_next_7_port, SUM(6) => PC_next_6_port, SUM(5) 
                           => PC_next_5_port, SUM(4) => PC_next_4_port, SUM(3) 
                           => PC_next_3_port, SUM(2) => PC_next_2_port, SUM(1) 
                           => PC_next_1_port, SUM(0) => PC_next_0_port);
   PC_reg_31_inst : DFFR_X1 port map( D => n288, CK => Clk, RN => n311, Q => 
                           Iaddr_31_port, QN => n192);
   U206 : BUF_X8 port map( A => Rst, Z => n311);
   U207 : CLKBUF_X1 port map( A => PC_next_31_port, Z => n296);
   U208 : INV_X1 port map( A => n191, ZN => Iaddr_0_port);
   U209 : OR2_X1 port map( A1 => PC_LATCH_EN_i, A2 => n192, ZN => n298);
   U210 : NAND2_X1 port map( A1 => n298, A2 => n96, ZN => n288);
   U211 : CLKBUF_X1 port map( A => IR_LATCH_EN_i, Z => n299);
   U212 : CLKBUF_X1 port map( A => IR_LATCH_EN_i, Z => n300);
   U213 : CLKBUF_X1 port map( A => IR_LATCH_EN_i, Z => n301);
   U214 : CLKBUF_X1 port map( A => IR_LATCH_EN_i, Z => n302);
   U215 : CLKBUF_X1 port map( A => IR_LATCH_EN_i, Z => n303);
   U216 : CLKBUF_X1 port map( A => IR_LATCH_EN_i, Z => n304);
   U217 : CLKBUF_X1 port map( A => NPC_LATCH_EN_i, Z => n305);
   U218 : CLKBUF_X1 port map( A => NPC_LATCH_EN_i, Z => n306);
   U219 : CLKBUF_X1 port map( A => NPC_LATCH_EN_i, Z => n307);
   U220 : CLKBUF_X1 port map( A => NPC_LATCH_EN_i, Z => n308);
   U221 : CLKBUF_X1 port map( A => NPC_LATCH_EN_i, Z => n309);
   U222 : CLKBUF_X1 port map( A => NPC_LATCH_EN_i, Z => n310);
   U223 : CLKBUF_X3 port map( A => Rst, Z => n312);
   U224 : CLKBUF_X3 port map( A => Rst, Z => n313);
   ROUT_LATCH_EN_i <= '0';

end SYN_dlx_rtl;
